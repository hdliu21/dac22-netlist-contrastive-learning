
module PlusArgTimeout ( clock, reset, io_count );
  input [31:0] io_count;
  input clock, reset;


endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_IBuf ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module Rocket ( clock, reset, io_interrupts_debug, io_interrupts_mtip, 
        io_interrupts_msip, io_interrupts_meip, io_interrupts_seip, 
        io_imem_might_request, io_imem_req_valid, io_imem_req_bits_pc, 
        io_imem_req_bits_speculative, io_imem_sfence_valid, 
        io_imem_sfence_bits_rs1, io_imem_sfence_bits_rs2, 
        io_imem_sfence_bits_addr, io_imem_resp_ready, io_imem_resp_valid, 
        io_imem_resp_bits_btb_taken, io_imem_resp_bits_btb_bridx, 
        io_imem_resp_bits_btb_entry, io_imem_resp_bits_btb_bht_history, 
        io_imem_resp_bits_pc, io_imem_resp_bits_data, 
        io_imem_resp_bits_xcpt_pf_inst, io_imem_resp_bits_xcpt_ae_inst, 
        io_imem_resp_bits_replay, io_imem_btb_update_valid, 
        io_imem_btb_update_bits_prediction_entry, io_imem_btb_update_bits_pc, 
        io_imem_btb_update_bits_isValid, io_imem_btb_update_bits_br_pc, 
        io_imem_btb_update_bits_cfiType, io_imem_bht_update_valid, 
        io_imem_bht_update_bits_prediction_history, io_imem_bht_update_bits_pc, 
        io_imem_bht_update_bits_branch, io_imem_bht_update_bits_taken, 
        io_imem_bht_update_bits_mispredict, io_imem_flush_icache, 
        io_dmem_req_ready, io_dmem_req_valid, io_dmem_req_bits_addr, 
        io_dmem_req_bits_tag, io_dmem_req_bits_cmd, io_dmem_req_bits_size, 
        io_dmem_req_bits_signed, io_dmem_req_bits_dprv, io_dmem_s1_kill, 
        io_dmem_s1_data_data, io_dmem_s2_nack, io_dmem_resp_valid, 
        io_dmem_resp_bits_tag, io_dmem_resp_bits_size, io_dmem_resp_bits_data, 
        io_dmem_resp_bits_replay, io_dmem_resp_bits_has_data, 
        io_dmem_resp_bits_data_word_bypass, io_dmem_replay_next, 
        io_dmem_s2_xcpt_ma_ld, io_dmem_s2_xcpt_ma_st, io_dmem_s2_xcpt_pf_ld, 
        io_dmem_s2_xcpt_pf_st, io_dmem_s2_xcpt_ae_ld, io_dmem_s2_xcpt_ae_st, 
        io_dmem_ordered, io_dmem_perf_release, io_dmem_perf_grant, 
        io_ptw_ptbr_mode, io_ptw_ptbr_ppn, io_ptw_sfence_valid, 
        io_ptw_sfence_bits_rs1, io_ptw_sfence_bits_rs2, 
        io_ptw_sfence_bits_addr, io_ptw_status_debug, io_ptw_status_dprv, 
        io_ptw_status_prv, io_ptw_status_mxr, io_ptw_status_sum, 
        io_ptw_pmp_0_cfg_l, io_ptw_pmp_0_cfg_a, io_ptw_pmp_0_cfg_x, 
        io_ptw_pmp_0_cfg_w, io_ptw_pmp_0_cfg_r, io_ptw_pmp_0_addr, 
        io_ptw_pmp_0_mask, io_ptw_pmp_1_cfg_l, io_ptw_pmp_1_cfg_a, 
        io_ptw_pmp_1_cfg_x, io_ptw_pmp_1_cfg_w, io_ptw_pmp_1_cfg_r, 
        io_ptw_pmp_1_addr, io_ptw_pmp_1_mask, io_ptw_pmp_2_cfg_l, 
        io_ptw_pmp_2_cfg_a, io_ptw_pmp_2_cfg_x, io_ptw_pmp_2_cfg_w, 
        io_ptw_pmp_2_cfg_r, io_ptw_pmp_2_addr, io_ptw_pmp_2_mask, 
        io_ptw_pmp_3_cfg_l, io_ptw_pmp_3_cfg_a, io_ptw_pmp_3_cfg_x, 
        io_ptw_pmp_3_cfg_w, io_ptw_pmp_3_cfg_r, io_ptw_pmp_3_addr, 
        io_ptw_pmp_3_mask, io_ptw_pmp_4_cfg_l, io_ptw_pmp_4_cfg_a, 
        io_ptw_pmp_4_cfg_x, io_ptw_pmp_4_cfg_w, io_ptw_pmp_4_cfg_r, 
        io_ptw_pmp_4_addr, io_ptw_pmp_4_mask, io_ptw_pmp_5_cfg_l, 
        io_ptw_pmp_5_cfg_a, io_ptw_pmp_5_cfg_x, io_ptw_pmp_5_cfg_w, 
        io_ptw_pmp_5_cfg_r, io_ptw_pmp_5_addr, io_ptw_pmp_5_mask, 
        io_ptw_pmp_6_cfg_l, io_ptw_pmp_6_cfg_a, io_ptw_pmp_6_cfg_x, 
        io_ptw_pmp_6_cfg_w, io_ptw_pmp_6_cfg_r, io_ptw_pmp_6_addr, 
        io_ptw_pmp_6_mask, io_ptw_pmp_7_cfg_l, io_ptw_pmp_7_cfg_a, 
        io_ptw_pmp_7_cfg_x, io_ptw_pmp_7_cfg_w, io_ptw_pmp_7_cfg_r, 
        io_ptw_pmp_7_addr, io_ptw_pmp_7_mask, io_ptw_customCSRs_csrs_0_value, 
        io_fpu_inst, io_fpu_fromint_data, io_fpu_fcsr_rm, 
        io_fpu_fcsr_flags_valid, io_fpu_fcsr_flags_bits, io_fpu_store_data, 
        io_fpu_toint_data, io_fpu_dmem_resp_val, io_fpu_dmem_resp_type, 
        io_fpu_dmem_resp_tag, io_fpu_dmem_resp_data, io_fpu_valid, 
        io_fpu_fcsr_rdy, io_fpu_nack_mem, io_fpu_illegal_rm, io_fpu_killx, 
        io_fpu_killm, io_fpu_dec_wen, io_fpu_dec_ren1, io_fpu_dec_ren2, 
        io_fpu_dec_ren3, io_fpu_sboard_set, io_fpu_sboard_clr, 
        io_fpu_sboard_clra, io_wfi );
  output [39:0] io_imem_req_bits_pc;
  output [38:0] io_imem_sfence_bits_addr;
  input [4:0] io_imem_resp_bits_btb_entry;
  input [7:0] io_imem_resp_bits_btb_bht_history;
  input [39:0] io_imem_resp_bits_pc;
  input [31:0] io_imem_resp_bits_data;
  output [4:0] io_imem_btb_update_bits_prediction_entry;
  output [38:0] io_imem_btb_update_bits_pc;
  output [38:0] io_imem_btb_update_bits_br_pc;
  output [1:0] io_imem_btb_update_bits_cfiType;
  output [7:0] io_imem_bht_update_bits_prediction_history;
  output [38:0] io_imem_bht_update_bits_pc;
  output [39:0] io_dmem_req_bits_addr;
  output [6:0] io_dmem_req_bits_tag;
  output [4:0] io_dmem_req_bits_cmd;
  output [1:0] io_dmem_req_bits_size;
  output [1:0] io_dmem_req_bits_dprv;
  output [63:0] io_dmem_s1_data_data;
  input [6:0] io_dmem_resp_bits_tag;
  input [1:0] io_dmem_resp_bits_size;
  input [63:0] io_dmem_resp_bits_data;
  input [63:0] io_dmem_resp_bits_data_word_bypass;
  output [3:0] io_ptw_ptbr_mode;
  output [43:0] io_ptw_ptbr_ppn;
  output [38:0] io_ptw_sfence_bits_addr;
  output [1:0] io_ptw_status_dprv;
  output [1:0] io_ptw_status_prv;
  output [1:0] io_ptw_pmp_0_cfg_a;
  output [29:0] io_ptw_pmp_0_addr;
  output [31:0] io_ptw_pmp_0_mask;
  output [1:0] io_ptw_pmp_1_cfg_a;
  output [29:0] io_ptw_pmp_1_addr;
  output [31:0] io_ptw_pmp_1_mask;
  output [1:0] io_ptw_pmp_2_cfg_a;
  output [29:0] io_ptw_pmp_2_addr;
  output [31:0] io_ptw_pmp_2_mask;
  output [1:0] io_ptw_pmp_3_cfg_a;
  output [29:0] io_ptw_pmp_3_addr;
  output [31:0] io_ptw_pmp_3_mask;
  output [1:0] io_ptw_pmp_4_cfg_a;
  output [29:0] io_ptw_pmp_4_addr;
  output [31:0] io_ptw_pmp_4_mask;
  output [1:0] io_ptw_pmp_5_cfg_a;
  output [29:0] io_ptw_pmp_5_addr;
  output [31:0] io_ptw_pmp_5_mask;
  output [1:0] io_ptw_pmp_6_cfg_a;
  output [29:0] io_ptw_pmp_6_addr;
  output [31:0] io_ptw_pmp_6_mask;
  output [1:0] io_ptw_pmp_7_cfg_a;
  output [29:0] io_ptw_pmp_7_addr;
  output [31:0] io_ptw_pmp_7_mask;
  output [63:0] io_ptw_customCSRs_csrs_0_value;
  output [31:0] io_fpu_inst;
  output [63:0] io_fpu_fromint_data;
  output [2:0] io_fpu_fcsr_rm;
  input [4:0] io_fpu_fcsr_flags_bits;
  input [63:0] io_fpu_store_data;
  input [63:0] io_fpu_toint_data;
  output [2:0] io_fpu_dmem_resp_type;
  output [4:0] io_fpu_dmem_resp_tag;
  output [63:0] io_fpu_dmem_resp_data;
  input [4:0] io_fpu_sboard_clra;
  input clock, reset, io_interrupts_debug, io_interrupts_mtip,
         io_interrupts_msip, io_interrupts_meip, io_interrupts_seip,
         io_imem_resp_valid, io_imem_resp_bits_btb_taken,
         io_imem_resp_bits_btb_bridx, io_imem_resp_bits_xcpt_pf_inst,
         io_imem_resp_bits_xcpt_ae_inst, io_imem_resp_bits_replay,
         io_dmem_req_ready, io_dmem_s2_nack, io_dmem_resp_valid,
         io_dmem_resp_bits_replay, io_dmem_resp_bits_has_data,
         io_dmem_replay_next, io_dmem_s2_xcpt_ma_ld, io_dmem_s2_xcpt_ma_st,
         io_dmem_s2_xcpt_pf_ld, io_dmem_s2_xcpt_pf_st, io_dmem_s2_xcpt_ae_ld,
         io_dmem_s2_xcpt_ae_st, io_dmem_ordered, io_dmem_perf_release,
         io_dmem_perf_grant, io_fpu_fcsr_flags_valid, io_fpu_fcsr_rdy,
         io_fpu_nack_mem, io_fpu_illegal_rm, io_fpu_dec_wen, io_fpu_dec_ren1,
         io_fpu_dec_ren2, io_fpu_dec_ren3, io_fpu_sboard_set,
         io_fpu_sboard_clr;
  output io_imem_might_request, io_imem_req_valid,
         io_imem_req_bits_speculative, io_imem_sfence_valid,
         io_imem_sfence_bits_rs1, io_imem_sfence_bits_rs2, io_imem_resp_ready,
         io_imem_btb_update_valid, io_imem_btb_update_bits_isValid,
         io_imem_bht_update_valid, io_imem_bht_update_bits_branch,
         io_imem_bht_update_bits_taken, io_imem_bht_update_bits_mispredict,
         io_imem_flush_icache, io_dmem_req_valid, io_dmem_req_bits_signed,
         io_dmem_s1_kill, io_ptw_sfence_valid, io_ptw_sfence_bits_rs1,
         io_ptw_sfence_bits_rs2, io_ptw_status_debug, io_ptw_status_mxr,
         io_ptw_status_sum, io_ptw_pmp_0_cfg_l, io_ptw_pmp_0_cfg_x,
         io_ptw_pmp_0_cfg_w, io_ptw_pmp_0_cfg_r, io_ptw_pmp_1_cfg_l,
         io_ptw_pmp_1_cfg_x, io_ptw_pmp_1_cfg_w, io_ptw_pmp_1_cfg_r,
         io_ptw_pmp_2_cfg_l, io_ptw_pmp_2_cfg_x, io_ptw_pmp_2_cfg_w,
         io_ptw_pmp_2_cfg_r, io_ptw_pmp_3_cfg_l, io_ptw_pmp_3_cfg_x,
         io_ptw_pmp_3_cfg_w, io_ptw_pmp_3_cfg_r, io_ptw_pmp_4_cfg_l,
         io_ptw_pmp_4_cfg_x, io_ptw_pmp_4_cfg_w, io_ptw_pmp_4_cfg_r,
         io_ptw_pmp_5_cfg_l, io_ptw_pmp_5_cfg_x, io_ptw_pmp_5_cfg_w,
         io_ptw_pmp_5_cfg_r, io_ptw_pmp_6_cfg_l, io_ptw_pmp_6_cfg_x,
         io_ptw_pmp_6_cfg_w, io_ptw_pmp_6_cfg_r, io_ptw_pmp_7_cfg_l,
         io_ptw_pmp_7_cfg_x, io_ptw_pmp_7_cfg_w, io_ptw_pmp_7_cfg_r,
         io_fpu_dmem_resp_val, io_fpu_valid, io_fpu_killx, io_fpu_killm,
         io_wfi;
  wire   io_imem_sfence_valid, io_imem_sfence_bits_rs1,
         io_imem_sfence_bits_rs2, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         ibuf_io_inst_0_valid, ibuf_io_inst_0_bits_replay,
         ibuf_io_inst_0_bits_rvc, csr_io_rw_cmd_2_, csr_io_decode_0_fp_illegal,
         csr_io_decode_0_fp_csr, csr_io_decode_0_read_illegal,
         csr_io_decode_0_write_illegal, csr_io_decode_0_write_flush,
         csr_io_decode_0_system_illegal, csr_io_csr_stall, csr_io_eret,
         csr_io_singleStep, csr_io_exception, csr_io_retire, csr_io_interrupt,
         csr_io_bp_0_control_action, csr_io_bp_0_control_m,
         csr_io_bp_0_control_s, csr_io_bp_0_control_u, csr_io_bp_0_control_x,
         csr_io_bp_0_control_w, csr_io_bp_0_control_r, bpu_io_xcpt_if,
         bpu_io_xcpt_ld, bpu_io_xcpt_st, bpu_io_debug_if, bpu_io_debug_ld,
         bpu_io_debug_st, alu_io_dw, alu_io_adder_out_39_, alu_io_cmp_out,
         div_io_req_ready, div_io_kill, div_io_resp_ready, div_io_resp_valid,
         wb_reg_replay, wb_reg_valid, wb_ctrl_mem, wb_reg_flush_pipe,
         ex_reg_valid, ex_reg_replay, ex_reg_xcpt_interrupt, mem_ctrl_jalr,
         mem_reg_sfence, n_T_844_10_, n_T_911_11, mem_reg_rvc,
         mem_br_target_39_, mem_br_target_38_, mem_br_target_37_,
         mem_br_target_36_, mem_br_target_35_, mem_br_target_34_,
         mem_br_target_33_, mem_br_target_32_, mem_br_target_31_,
         mem_br_target_30_, mem_br_target_29_, mem_br_target_28_,
         mem_br_target_27_, mem_br_target_26_, mem_br_target_25_,
         mem_br_target_24_, mem_br_target_23_, mem_br_target_22_,
         mem_br_target_21_, mem_br_target_20_, mem_br_target_19_,
         mem_br_target_18_, mem_br_target_17_, mem_br_target_16_,
         mem_br_target_15_, mem_br_target_14_, mem_br_target_13_,
         mem_br_target_12_, mem_br_target_11_, mem_br_target_10_,
         mem_br_target_9_, mem_br_target_8_, mem_br_target_7_,
         mem_br_target_6_, mem_br_target_5_, mem_br_target_4_,
         mem_br_target_3_, mem_br_target_2_, mem_br_target_1_, mem_reg_valid,
         id_ctrl_mem_cmd_2_, id_ctrl_wfd, id_ctrl_wxd, id_reg_fence,
         ex_reg_inst_31_, ex_ctrl_wxd, mem_ctrl_wxd, mem_ctrl_mem,
         ex_reg_rs_bypass_1, ex_ctrl_sel_alu1_0_, ex_reg_rvc, ex_ctrl_jalr,
         ex_ctrl_mem, ex_ctrl_div, ex_ctrl_wfd, mem_reg_slow_bypass,
         mem_ctrl_wfd, wb_ctrl_wxd, wb_ctrl_div, wb_ctrl_wfd, blocked,
         id_reg_pause, n_GEN_9, n_T_731, do_bypass_1, n_T_760, ex_reg_load_use,
         mem_reg_replay, mem_reg_xcpt_interrupt, mem_pc_valid, mem_reg_xcpt,
         mem_reg_flush_pipe, ex_ctrl_rxs2, mem_reg_load, mem_reg_store,
         wb_ctrl_fence_i, wb_reg_sfence, n_T_1057, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N271, N274, N275, N279, N282, N283,
         N284, N286, N290, ex_ctrl_jal, N303, N304, N369, N370, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503,
         N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514,
         N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N526,
         N529, N530, N533, N535, N536, N598, N599, N600, N601, N602, N603,
         N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658,
         N659, N660, N661, N672, N673, N678, N679, N682, N683, N684, N685,
         N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696,
         N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707,
         N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729,
         N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740,
         N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751,
         N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, net34469, net34475, net34480, net34485,
         net34490, net34495, net34500, net34505, net34510, net34515, net34520,
         net34525, net34530, net34535, net34540, net34545, net34550, net34555,
         net34560, net34565, net34570, net34575, net34580, net34585, net34590,
         net34595, net34600, net34605, net34610, net34615, net34620, net34625,
         net34630, net34635, net34640, net34645, net34650, net34655, net34660,
         net34665, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n66, n67, n68, n69, n71, n72, n73, n74, n75, n76, n80, n98, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n308, n309, n310, n312, n313, n314,
         n315, n317, n318, n319, n320, n322, n323, n326, n369, n370, n406,
         n407, n546, n555, n559, n560, n561, n569, n570, n572, n576, n586,
         n588, n589, n590, n591, n592, n594, n595, n596, n598, n711, n882,
         n996, n997, n1262, n1279, n1281, n1431, n1531, n1532, n1589, n1612,
         n1628, n1699, n1820, n1821, n1822, n1823, n1828, n1829, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1855, n1856, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2238, n2239, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2492,
         n2493, n2495, n2496, n2497, n2498, n2501, n2507, n2510, n2512, n2514,
         n2515, n2516, n2518, n2521, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2541, n2542, n2543, n2544, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3046, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9417, n9418, n9421, n9422,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         ibuf_SYNOPSYS_UNCONNECTED_7, ibuf_SYNOPSYS_UNCONNECTED_6,
         ibuf_SYNOPSYS_UNCONNECTED_5, ibuf_SYNOPSYS_UNCONNECTED_4,
         ibuf_SYNOPSYS_UNCONNECTED_3, ibuf_SYNOPSYS_UNCONNECTED_2,
         ibuf_SYNOPSYS_UNCONNECTED_1, ibuf_io_inst_0_bits_inst_rs3_4_,
         ibuf_io_inst_0_bits_inst_rs3_2_, ibuf_n121, ibuf_n120, ibuf_n119,
         ibuf_n118, ibuf_n117, ibuf_n116, ibuf_n115, ibuf_n114, ibuf_n113,
         ibuf_n112, ibuf_n111, ibuf_n110, ibuf_n109, ibuf_n108, ibuf_n107,
         ibuf_n106, ibuf_n105, ibuf_n104, ibuf_n103, ibuf_n102, ibuf_n101,
         ibuf_n100, ibuf_n99, ibuf_n98, ibuf_n97, ibuf_n96, ibuf_n95, ibuf_n94,
         ibuf_n93, ibuf_n92, ibuf_n91, ibuf_n90, ibuf_n89, ibuf_n88, ibuf_n87,
         ibuf_n86, ibuf_n85, ibuf_n84, ibuf_n83, ibuf_n82, ibuf_n81, ibuf_n80,
         ibuf_n79, ibuf_n78, ibuf_n77, ibuf_n76, ibuf_n75, ibuf_n74, ibuf_n73,
         ibuf_n72, ibuf_n71, ibuf_n70, ibuf_n69, ibuf_n68, ibuf_n67, ibuf_n66,
         ibuf_n65, ibuf_n64, ibuf_n63, ibuf_n62, ibuf_n61, ibuf_n60, ibuf_n59,
         ibuf_n58, ibuf_n57, ibuf_n56, ibuf_n55, ibuf_n54, ibuf_n53, ibuf_n52,
         ibuf_n51, ibuf_n50, ibuf_n49, ibuf_n48, ibuf_n47, ibuf_n46, ibuf_n45,
         ibuf_n43, ibuf_n42, ibuf_n41, ibuf_n39, ibuf_n38, ibuf_n37, ibuf_n36,
         ibuf_n35, ibuf_n34, ibuf_n33, ibuf_n32, ibuf_n31, ibuf_n30, ibuf_n29,
         ibuf_n28, ibuf_n27, ibuf_n26, ibuf_n25, ibuf_n24, ibuf_n23, ibuf_n20,
         ibuf_n19, ibuf_n18, ibuf_n11, ibuf_n10, ibuf_n9, ibuf_n8, ibuf_n7,
         ibuf_n5, ibuf_n40, ibuf_n12, ibuf_net35341, ibuf_N51,
         ibuf_buf__xcpt_ae_inst, ibuf_buf__xcpt_pf_inst, ibuf_n_T_55_84_,
         ibuf_n_T_55_85_, ibuf_n_T_55_91_, ibuf_n_T_27_0_, ibuf_buf__replay,
         ibuf_n131, ibuf_n130, ibuf_n129, ibuf_n128, ibuf_n127, ibuf_n126,
         ibuf_n125, ibuf_n124, ibuf_n123, ibuf_n122, ibuf_RVCExpander_n353,
         ibuf_RVCExpander_n352, ibuf_RVCExpander_n351, ibuf_RVCExpander_n350,
         ibuf_RVCExpander_n349, ibuf_RVCExpander_n348, ibuf_RVCExpander_n347,
         ibuf_RVCExpander_n346, ibuf_RVCExpander_n345, ibuf_RVCExpander_n344,
         ibuf_RVCExpander_n343, ibuf_RVCExpander_n342, ibuf_RVCExpander_n341,
         ibuf_RVCExpander_n340, ibuf_RVCExpander_n339, ibuf_RVCExpander_n338,
         ibuf_RVCExpander_n337, ibuf_RVCExpander_n336, ibuf_RVCExpander_n335,
         ibuf_RVCExpander_n334, ibuf_RVCExpander_n333, ibuf_RVCExpander_n332,
         ibuf_RVCExpander_n331, ibuf_RVCExpander_n330, ibuf_RVCExpander_n329,
         ibuf_RVCExpander_n328, ibuf_RVCExpander_n327, ibuf_RVCExpander_n326,
         ibuf_RVCExpander_n325, ibuf_RVCExpander_n324, ibuf_RVCExpander_n323,
         ibuf_RVCExpander_n322, ibuf_RVCExpander_n321, ibuf_RVCExpander_n320,
         ibuf_RVCExpander_n319, ibuf_RVCExpander_n318, ibuf_RVCExpander_n317,
         ibuf_RVCExpander_n316, ibuf_RVCExpander_n315, ibuf_RVCExpander_n314,
         ibuf_RVCExpander_n313, ibuf_RVCExpander_n312, ibuf_RVCExpander_n311,
         ibuf_RVCExpander_n310, ibuf_RVCExpander_n309, ibuf_RVCExpander_n308,
         ibuf_RVCExpander_n307, ibuf_RVCExpander_n306, ibuf_RVCExpander_n305,
         ibuf_RVCExpander_n304, ibuf_RVCExpander_n303, ibuf_RVCExpander_n302,
         ibuf_RVCExpander_n301, ibuf_RVCExpander_n300, ibuf_RVCExpander_n299,
         ibuf_RVCExpander_n298, ibuf_RVCExpander_n297, ibuf_RVCExpander_n296,
         ibuf_RVCExpander_n295, ibuf_RVCExpander_n294, ibuf_RVCExpander_n293,
         ibuf_RVCExpander_n292, ibuf_RVCExpander_n291, ibuf_RVCExpander_n290,
         ibuf_RVCExpander_n289, ibuf_RVCExpander_n288, ibuf_RVCExpander_n287,
         ibuf_RVCExpander_n286, ibuf_RVCExpander_n285, ibuf_RVCExpander_n284,
         ibuf_RVCExpander_n283, ibuf_RVCExpander_n282, ibuf_RVCExpander_n281,
         ibuf_RVCExpander_n280, ibuf_RVCExpander_n279, ibuf_RVCExpander_n278,
         ibuf_RVCExpander_n277, ibuf_RVCExpander_n276, ibuf_RVCExpander_n275,
         ibuf_RVCExpander_n274, ibuf_RVCExpander_n273, ibuf_RVCExpander_n272,
         ibuf_RVCExpander_n271, ibuf_RVCExpander_n270, ibuf_RVCExpander_n269,
         ibuf_RVCExpander_n268, ibuf_RVCExpander_n267, ibuf_RVCExpander_n266,
         ibuf_RVCExpander_n265, ibuf_RVCExpander_n264, ibuf_RVCExpander_n263,
         ibuf_RVCExpander_n262, ibuf_RVCExpander_n261, ibuf_RVCExpander_n260,
         ibuf_RVCExpander_n259, ibuf_RVCExpander_n258, ibuf_RVCExpander_n257,
         ibuf_RVCExpander_n256, ibuf_RVCExpander_n255, ibuf_RVCExpander_n254,
         ibuf_RVCExpander_n253, ibuf_RVCExpander_n252, ibuf_RVCExpander_n251,
         ibuf_RVCExpander_n250, ibuf_RVCExpander_n249, ibuf_RVCExpander_n248,
         ibuf_RVCExpander_n247, ibuf_RVCExpander_n246, ibuf_RVCExpander_n245,
         ibuf_RVCExpander_n244, ibuf_RVCExpander_n243, ibuf_RVCExpander_n242,
         ibuf_RVCExpander_n241, ibuf_RVCExpander_n240, ibuf_RVCExpander_n239,
         ibuf_RVCExpander_n238, ibuf_RVCExpander_n237, ibuf_RVCExpander_n236,
         ibuf_RVCExpander_n235, ibuf_RVCExpander_n234, ibuf_RVCExpander_n233,
         ibuf_RVCExpander_n232, ibuf_RVCExpander_n231, ibuf_RVCExpander_n230,
         ibuf_RVCExpander_n229, ibuf_RVCExpander_n228, ibuf_RVCExpander_n227,
         ibuf_RVCExpander_n226, ibuf_RVCExpander_n225, ibuf_RVCExpander_n224,
         ibuf_RVCExpander_n223, ibuf_RVCExpander_n222, ibuf_RVCExpander_n221,
         ibuf_RVCExpander_n220, ibuf_RVCExpander_n219, ibuf_RVCExpander_n218,
         ibuf_RVCExpander_n217, ibuf_RVCExpander_n216, ibuf_RVCExpander_n215,
         ibuf_RVCExpander_n214, ibuf_RVCExpander_n213, ibuf_RVCExpander_n212,
         ibuf_RVCExpander_n211, ibuf_RVCExpander_n210, ibuf_RVCExpander_n209,
         ibuf_RVCExpander_n208, ibuf_RVCExpander_n207, ibuf_RVCExpander_n206,
         ibuf_RVCExpander_n205, ibuf_RVCExpander_n204, ibuf_RVCExpander_n203,
         ibuf_RVCExpander_n202, ibuf_RVCExpander_n201, ibuf_RVCExpander_n200,
         ibuf_RVCExpander_n199, ibuf_RVCExpander_n198, ibuf_RVCExpander_n197,
         ibuf_RVCExpander_n196, ibuf_RVCExpander_n195, ibuf_RVCExpander_n194,
         ibuf_RVCExpander_n193, ibuf_RVCExpander_n192, ibuf_RVCExpander_n191,
         ibuf_RVCExpander_n190, ibuf_RVCExpander_n189, ibuf_RVCExpander_n188,
         ibuf_RVCExpander_n187, ibuf_RVCExpander_n186, ibuf_RVCExpander_n185,
         ibuf_RVCExpander_n184, ibuf_RVCExpander_n183, ibuf_RVCExpander_n182,
         ibuf_RVCExpander_n181, ibuf_RVCExpander_n180, ibuf_RVCExpander_n179,
         ibuf_RVCExpander_n178, ibuf_RVCExpander_n177, ibuf_RVCExpander_n176,
         ibuf_RVCExpander_n175, ibuf_RVCExpander_n174, ibuf_RVCExpander_n173,
         ibuf_RVCExpander_n172, ibuf_RVCExpander_n171, ibuf_RVCExpander_n170,
         ibuf_RVCExpander_n169, ibuf_RVCExpander_n168, ibuf_RVCExpander_n167,
         ibuf_RVCExpander_n166, ibuf_RVCExpander_n165, ibuf_RVCExpander_n164,
         ibuf_RVCExpander_n163, ibuf_RVCExpander_n162, ibuf_RVCExpander_n161,
         ibuf_RVCExpander_n160, ibuf_RVCExpander_n159, ibuf_RVCExpander_n158,
         ibuf_RVCExpander_n157, ibuf_RVCExpander_n156, ibuf_RVCExpander_n155,
         ibuf_RVCExpander_n154, ibuf_RVCExpander_n153, ibuf_RVCExpander_n152,
         ibuf_RVCExpander_n151, ibuf_RVCExpander_n150, ibuf_RVCExpander_n149,
         ibuf_RVCExpander_n148, ibuf_RVCExpander_n147, ibuf_RVCExpander_n146,
         ibuf_RVCExpander_n145, ibuf_RVCExpander_n144, ibuf_RVCExpander_n143,
         ibuf_RVCExpander_n142, ibuf_RVCExpander_n141, ibuf_RVCExpander_n140,
         ibuf_RVCExpander_n139, ibuf_RVCExpander_n138, ibuf_RVCExpander_n137,
         ibuf_RVCExpander_n136, ibuf_RVCExpander_n135, ibuf_RVCExpander_n134,
         ibuf_RVCExpander_n133, ibuf_RVCExpander_n132, ibuf_RVCExpander_n131,
         ibuf_RVCExpander_n130, ibuf_RVCExpander_n129, ibuf_RVCExpander_n128,
         ibuf_RVCExpander_n127, ibuf_RVCExpander_n126, ibuf_RVCExpander_n125,
         ibuf_RVCExpander_n124, ibuf_RVCExpander_n123, ibuf_RVCExpander_n122,
         ibuf_RVCExpander_n121, ibuf_RVCExpander_n120, ibuf_RVCExpander_n119,
         ibuf_RVCExpander_n118, ibuf_RVCExpander_n117, ibuf_RVCExpander_n116,
         ibuf_RVCExpander_n115, ibuf_RVCExpander_n114, ibuf_RVCExpander_n113,
         ibuf_RVCExpander_n112, ibuf_RVCExpander_n111, ibuf_RVCExpander_n110,
         ibuf_RVCExpander_n109, ibuf_RVCExpander_n108, ibuf_RVCExpander_n107,
         ibuf_RVCExpander_n106, ibuf_RVCExpander_n105, ibuf_RVCExpander_n104,
         ibuf_RVCExpander_n103, ibuf_RVCExpander_n102, ibuf_RVCExpander_n101,
         ibuf_RVCExpander_n100, ibuf_RVCExpander_n99, ibuf_RVCExpander_n98,
         ibuf_RVCExpander_n97, ibuf_RVCExpander_n96, ibuf_RVCExpander_n95,
         ibuf_RVCExpander_n94, ibuf_RVCExpander_n93, ibuf_RVCExpander_n92,
         ibuf_RVCExpander_n91, ibuf_RVCExpander_n90, ibuf_RVCExpander_n89,
         ibuf_RVCExpander_n88, ibuf_RVCExpander_n87, ibuf_RVCExpander_n86,
         ibuf_RVCExpander_n85, ibuf_RVCExpander_n84, ibuf_RVCExpander_n83,
         ibuf_RVCExpander_n82, ibuf_RVCExpander_n81, ibuf_RVCExpander_n80,
         ibuf_RVCExpander_n79, ibuf_RVCExpander_n78, ibuf_RVCExpander_n77,
         ibuf_RVCExpander_n76, ibuf_RVCExpander_n75, ibuf_RVCExpander_n74,
         ibuf_RVCExpander_n73, ibuf_RVCExpander_n72, ibuf_RVCExpander_n71,
         ibuf_RVCExpander_n70, ibuf_RVCExpander_n68, ibuf_RVCExpander_n67,
         ibuf_RVCExpander_n66, ibuf_RVCExpander_n65, ibuf_RVCExpander_n64,
         ibuf_RVCExpander_n63, ibuf_RVCExpander_n62, ibuf_RVCExpander_n61,
         ibuf_RVCExpander_n60, ibuf_RVCExpander_n59, ibuf_RVCExpander_n58,
         ibuf_RVCExpander_n57, ibuf_RVCExpander_n56, ibuf_RVCExpander_n55,
         ibuf_RVCExpander_n54, ibuf_RVCExpander_n53, ibuf_RVCExpander_n52,
         ibuf_RVCExpander_n51, ibuf_RVCExpander_n50, ibuf_RVCExpander_n49,
         ibuf_RVCExpander_n48, ibuf_RVCExpander_n47, ibuf_RVCExpander_n46,
         ibuf_RVCExpander_n40, ibuf_RVCExpander_n39, ibuf_RVCExpander_n38,
         ibuf_RVCExpander_n37, ibuf_RVCExpander_n36, ibuf_RVCExpander_n35,
         ibuf_RVCExpander_n34, ibuf_RVCExpander_n32, ibuf_RVCExpander_n30,
         ibuf_RVCExpander_n29, ibuf_RVCExpander_n28, ibuf_RVCExpander_n27,
         ibuf_RVCExpander_n26, ibuf_RVCExpander_n25, ibuf_RVCExpander_n24,
         ibuf_RVCExpander_n23, ibuf_RVCExpander_n22, ibuf_RVCExpander_n21,
         ibuf_RVCExpander_n20, ibuf_RVCExpander_n19, ibuf_RVCExpander_n18,
         ibuf_RVCExpander_n17, ibuf_RVCExpander_n15, ibuf_RVCExpander_n13,
         ibuf_RVCExpander_n12, ibuf_RVCExpander_n11, ibuf_RVCExpander_n10,
         ibuf_RVCExpander_n9, ibuf_RVCExpander_n8, ibuf_RVCExpander_n7,
         ibuf_RVCExpander_n6, ibuf_RVCExpander_n5, ibuf_RVCExpander_n3,
         ibuf_RVCExpander_n2, ibuf_RVCExpander_n1, ibuf_RVCExpander_n354,
         csr_SYNOPSYS_UNCONNECTED_10, csr_SYNOPSYS_UNCONNECTED_9,
         csr_SYNOPSYS_UNCONNECTED_8, csr_SYNOPSYS_UNCONNECTED_7,
         csr_SYNOPSYS_UNCONNECTED_6, csr_SYNOPSYS_UNCONNECTED_5,
         csr_SYNOPSYS_UNCONNECTED_4, csr_SYNOPSYS_UNCONNECTED_3,
         csr_SYNOPSYS_UNCONNECTED_2, csr_SYNOPSYS_UNCONNECTED_1, csr_n1917,
         csr_n1915, csr_n1914, csr_n1913, csr_n1912, csr_n1911, csr_n1910,
         csr_n1909, csr_n1908, csr_n1907, csr_n1906, csr_n1905, csr_n1904,
         csr_n1903, csr_n1902, csr_n1901, csr_n1900, csr_n1899, csr_n1898,
         csr_n1897, csr_n1896, csr_n1895, csr_n1894, csr_n1893, csr_n1892,
         csr_n1891, csr_n1890, csr_n1889, csr_n1888, csr_n1887, csr_n1886,
         csr_n1885, csr_n1884, csr_n1883, csr_n1882, csr_n1881, csr_n1880,
         csr_n1879, csr_n1878, csr_n1877, csr_n1876, csr_n1875, csr_n1874,
         csr_n1873, csr_n1872, csr_n1871, csr_n1870, csr_n1869, csr_n1868,
         csr_n1867, csr_n1866, csr_n1865, csr_n1864, csr_n1863, csr_n1862,
         csr_n1861, csr_n1860, csr_n1859, csr_n1858, csr_n1857, csr_n1856,
         csr_n1855, csr_n1854, csr_n1853, csr_n1852, csr_n1851, csr_n1850,
         csr_n1849, csr_n1848, csr_n1847, csr_n1846, csr_n1845, csr_n1844,
         csr_n1843, csr_n1842, csr_n1841, csr_n1840, csr_n1839, csr_n1838,
         csr_n1837, csr_n1836, csr_n1835, csr_n1834, csr_n1833, csr_n1832,
         csr_n1831, csr_n1830, csr_n1829, csr_n1828, csr_n1827, csr_n1826,
         csr_n1825, csr_n1824, csr_n1823, csr_n1822, csr_n1821, csr_n1820,
         csr_n1819, csr_n1818, csr_n1817, csr_n1816, csr_n1815, csr_n1814,
         csr_n1813, csr_n1812, csr_n1811, csr_n1810, csr_n1809, csr_n1808,
         csr_n1807, csr_n1806, csr_n1805, csr_n1804, csr_n1803, csr_n1802,
         csr_n1801, csr_n1800, csr_n1799, csr_n1798, csr_n1797, csr_n1796,
         csr_n1795, csr_n1794, csr_n1793, csr_n1792, csr_n1791, csr_n1790,
         csr_n1789, csr_n1788, csr_n1787, csr_n1786, csr_n1785, csr_n1784,
         csr_n1783, csr_n1782, csr_n1781, csr_n1780, csr_n1779, csr_n1778,
         csr_n1777, csr_n1776, csr_n1775, csr_n1774, csr_n1773, csr_n1772,
         csr_n1771, csr_n1770, csr_n1769, csr_n1768, csr_n1767, csr_n1766,
         csr_n1765, csr_n1764, csr_n1763, csr_n1762, csr_n1761, csr_n1760,
         csr_n1759, csr_n1758, csr_n1757, csr_n1756, csr_n1755, csr_n1754,
         csr_n1753, csr_n1752, csr_n1751, csr_n1750, csr_n1749, csr_n1748,
         csr_n1747, csr_n1746, csr_n1745, csr_n1744, csr_n1743, csr_n1742,
         csr_n1741, csr_n1740, csr_n1739, csr_n1738, csr_n1737, csr_n1736,
         csr_n1735, csr_n1734, csr_n1733, csr_n1732, csr_n1731, csr_n1730,
         csr_n1729, csr_n1728, csr_n1727, csr_n1726, csr_n1725, csr_n1724,
         csr_n1723, csr_n1722, csr_n1721, csr_n1720, csr_n1719, csr_n1718,
         csr_n1717, csr_n1716, csr_n1715, csr_n1714, csr_n1713, csr_n1712,
         csr_n1711, csr_n1710, csr_n1709, csr_n1708, csr_n1707, csr_n1706,
         csr_n1705, csr_n1704, csr_n1703, csr_n1702, csr_n1701, csr_n1700,
         csr_n1699, csr_n1698, csr_n1697, csr_n1696, csr_n1695, csr_n1694,
         csr_n1693, csr_n1692, csr_n1691, csr_n1690, csr_n1689, csr_n1688,
         csr_n1687, csr_n1686, csr_n1685, csr_n1684, csr_n1683, csr_n1682,
         csr_n1681, csr_n1680, csr_n1679, csr_n1678, csr_n1677, csr_n1676,
         csr_n1675, csr_n1674, csr_n1673, csr_n1672, csr_n1671, csr_n1670,
         csr_n1669, csr_n1668, csr_n1667, csr_n1666, csr_n1665, csr_n1664,
         csr_n1663, csr_n1662, csr_n1661, csr_n1660, csr_n1659, csr_n1658,
         csr_n1657, csr_n1656, csr_n1655, csr_n1654, csr_n1653, csr_n1652,
         csr_n1651, csr_n1650, csr_n1649, csr_n1648, csr_n1647, csr_n1646,
         csr_n1645, csr_n1644, csr_n1643, csr_n1642, csr_n1641, csr_n1640,
         csr_n1639, csr_n1638, csr_n1637, csr_n1636, csr_n1635, csr_n1634,
         csr_n1633, csr_n1632, csr_n1631, csr_n1630, csr_n1629, csr_n1628,
         csr_n1627, csr_n1626, csr_n1625, csr_n1624, csr_n1623, csr_n1622,
         csr_n1621, csr_n1620, csr_n1619, csr_n1618, csr_n1617, csr_n1616,
         csr_n1615, csr_n1614, csr_n1613, csr_n1612, csr_n1611, csr_n1610,
         csr_n1609, csr_n1608, csr_n1607, csr_n1606, csr_n1605, csr_n1604,
         csr_n1603, csr_n1602, csr_n1601, csr_n1600, csr_n1599, csr_n1598,
         csr_n1597, csr_n1596, csr_n1595, csr_n1594, csr_n1593, csr_n1592,
         csr_n1591, csr_n1590, csr_n1589, csr_n1588, csr_n1587, csr_n1586,
         csr_n1585, csr_n1584, csr_n1583, csr_n1582, csr_n1581, csr_n1580,
         csr_n1579, csr_n1578, csr_n1577, csr_n1576, csr_n1575, csr_n1574,
         csr_n1573, csr_n1572, csr_n1571, csr_n1570, csr_n1569, csr_n1568,
         csr_n1567, csr_n1566, csr_n1565, csr_n1564, csr_n1563, csr_n1562,
         csr_n1561, csr_n1560, csr_n1559, csr_n1558, csr_n1557, csr_n1556,
         csr_n1555, csr_n1554, csr_n1553, csr_n1552, csr_n1551, csr_n1550,
         csr_n1549, csr_n1548, csr_n1547, csr_n1546, csr_n1545, csr_n1544,
         csr_n1543, csr_n1542, csr_n1541, csr_n1540, csr_n1539, csr_n1538,
         csr_n1537, csr_n1536, csr_n1535, csr_n1534, csr_n1533, csr_n1532,
         csr_n1531, csr_n1530, csr_n1529, csr_n1528, csr_n1527, csr_n1526,
         csr_n1525, csr_n1524, csr_n1523, csr_n1522, csr_n1521, csr_n1520,
         csr_n1519, csr_n1518, csr_n1517, csr_n1516, csr_n1515, csr_n1514,
         csr_n1513, csr_n1512, csr_n1511, csr_n1510, csr_n1509, csr_n1508,
         csr_n1507, csr_n1506, csr_n1505, csr_n1504, csr_n1503, csr_n1502,
         csr_n1501, csr_n1500, csr_n1499, csr_n1498, csr_n1497, csr_n1496,
         csr_n1495, csr_n1494, csr_n1493, csr_n1492, csr_n1491, csr_n1490,
         csr_n1489, csr_n1488, csr_n1487, csr_n1486, csr_n1485, csr_n1484,
         csr_n1483, csr_n1482, csr_n1481, csr_n1480, csr_n1479, csr_n1478,
         csr_n1477, csr_n1476, csr_n1475, csr_n1474, csr_n1473, csr_n1472,
         csr_n1471, csr_n1470, csr_n1469, csr_n1468, csr_n1467, csr_n1466,
         csr_n1465, csr_n1464, csr_n1463, csr_n1462, csr_n1461, csr_n1460,
         csr_n1459, csr_n1458, csr_n1457, csr_n1456, csr_n1455, csr_n1454,
         csr_n1453, csr_n1452, csr_n1451, csr_n1450, csr_n1449, csr_n1448,
         csr_n1447, csr_n1446, csr_n1445, csr_n1444, csr_n1443, csr_n1442,
         csr_n1441, csr_n1440, csr_n1439, csr_n1438, csr_n1437, csr_n1436,
         csr_n1435, csr_n1434, csr_n1433, csr_n1432, csr_n1431, csr_n1430,
         csr_n1429, csr_n1428, csr_n1427, csr_n1426, csr_n1425, csr_n1424,
         csr_n1423, csr_n1422, csr_n1421, csr_n1420, csr_n1419, csr_n1418,
         csr_n1417, csr_n1416, csr_n1415, csr_n1414, csr_n1413, csr_n1412,
         csr_n1411, csr_n1410, csr_n1409, csr_n1408, csr_n1407, csr_n1406,
         csr_n1405, csr_n1404, csr_n1403, csr_n1402, csr_n1401, csr_n1400,
         csr_n1399, csr_n1398, csr_n1397, csr_n1396, csr_n1395, csr_n1394,
         csr_n1393, csr_n1392, csr_n1391, csr_n1390, csr_n1389, csr_n1388,
         csr_n1387, csr_n1386, csr_n1385, csr_n1384, csr_n1383, csr_n1382,
         csr_n1381, csr_n1380, csr_n1379, csr_n1378, csr_n1377, csr_n1376,
         csr_n1375, csr_n1374, csr_n1373, csr_n1372, csr_n1371, csr_n1370,
         csr_n1369, csr_n1368, csr_n1367, csr_n1366, csr_n1365, csr_n1364,
         csr_n1363, csr_n1362, csr_n1361, csr_n1360, csr_n1359, csr_n1358,
         csr_n1357, csr_n1356, csr_n1355, csr_n1354, csr_n1353, csr_n1352,
         csr_n1351, csr_n1350, csr_n1349, csr_n1348, csr_n1347, csr_n1345,
         csr_n1344, csr_n1343, csr_n1342, csr_n1341, csr_n1340, csr_n1339,
         csr_n1338, csr_n1337, csr_n1336, csr_n1335, csr_n1334, csr_n1333,
         csr_n1332, csr_n1331, csr_n1330, csr_n1329, csr_n1328, csr_n1327,
         csr_n1326, csr_n1325, csr_n1324, csr_n1323, csr_n1322, csr_n1321,
         csr_n1320, csr_n1319, csr_n1318, csr_n1317, csr_n1316, csr_n1315,
         csr_n1314, csr_n1313, csr_n1312, csr_n1311, csr_n1310, csr_n1309,
         csr_n1308, csr_n1307, csr_n1306, csr_n1305, csr_n1304, csr_n1303,
         csr_n1302, csr_n1301, csr_n1300, csr_n1299, csr_n1298, csr_n1297,
         csr_n1296, csr_n1295, csr_n1294, csr_n1293, csr_n1292, csr_n1291,
         csr_n1290, csr_n1289, csr_n1288, csr_n1287, csr_n1286, csr_n1285,
         csr_n1284, csr_n1283, csr_n1282, csr_n1281, csr_n1280, csr_n1279,
         csr_n1278, csr_n1277, csr_n1276, csr_n1275, csr_n1274, csr_n1273,
         csr_n1272, csr_n1271, csr_n1270, csr_n1269, csr_n1268, csr_n1267,
         csr_n1266, csr_n1265, csr_n1264, csr_n1263, csr_n1262, csr_n1261,
         csr_n1260, csr_n1259, csr_n1258, csr_n1257, csr_n1256, csr_n1255,
         csr_n1254, csr_n1253, csr_n1252, csr_n1251, csr_n1250, csr_n1249,
         csr_n1248, csr_n1247, csr_n1246, csr_n1245, csr_n1244, csr_n1243,
         csr_n1242, csr_n1241, csr_n1240, csr_n1239, csr_n1238, csr_n1237,
         csr_n1236, csr_n1235, csr_n1234, csr_n1233, csr_n1232, csr_n1231,
         csr_n1230, csr_n1229, csr_n1228, csr_n1227, csr_n1226, csr_n1225,
         csr_n1224, csr_n1223, csr_n1222, csr_n1221, csr_n1220, csr_n1219,
         csr_n1218, csr_n1217, csr_n1216, csr_n1215, csr_n1214, csr_n1213,
         csr_n1212, csr_n1211, csr_n1210, csr_n1209, csr_n1208, csr_n1207,
         csr_n1206, csr_n1205, csr_n1204, csr_n1203, csr_n1202, csr_n1201,
         csr_n1200, csr_n1199, csr_n1198, csr_n1197, csr_n1196, csr_n1195,
         csr_n1194, csr_n1193, csr_n1192, csr_n1191, csr_n1190, csr_n1189,
         csr_n1188, csr_n1187, csr_n1186, csr_n1185, csr_n1184, csr_n1183,
         csr_n1182, csr_n1181, csr_n1180, csr_n1179, csr_n1178, csr_n1177,
         csr_n1176, csr_n1175, csr_n1174, csr_n1173, csr_n1172, csr_n1171,
         csr_n1170, csr_n1169, csr_n1168, csr_n1167, csr_n1166, csr_n1165,
         csr_n1164, csr_n1163, csr_n1162, csr_n1161, csr_n1160, csr_n1159,
         csr_n1158, csr_n1157, csr_n1156, csr_n1155, csr_n1154, csr_n1153,
         csr_n1152, csr_n1151, csr_n1150, csr_n1149, csr_n1148, csr_n1147,
         csr_n1146, csr_n1145, csr_n1144, csr_n1143, csr_n1142, csr_n1141,
         csr_n1140, csr_n1139, csr_n1138, csr_n1137, csr_n1136, csr_n1135,
         csr_n1134, csr_n1133, csr_n1132, csr_n1131, csr_n1130, csr_n1129,
         csr_n1128, csr_n1127, csr_n1126, csr_n1125, csr_n1124, csr_n1123,
         csr_n1122, csr_n1121, csr_n1120, csr_n1119, csr_n1118, csr_n1117,
         csr_n1116, csr_n1115, csr_n1114, csr_n1113, csr_n1112, csr_n1111,
         csr_n1110, csr_n1109, csr_n1108, csr_n1107, csr_n1106, csr_n1105,
         csr_n1104, csr_n1103, csr_n1102, csr_n1101, csr_n1100, csr_n1099,
         csr_n1098, csr_n1097, csr_n1096, csr_n1095, csr_n1094, csr_n1093,
         csr_n1092, csr_n1091, csr_n1090, csr_n1089, csr_n1088, csr_n1087,
         csr_n1086, csr_n1085, csr_n1084, csr_n1083, csr_n1082, csr_n1081,
         csr_n1080, csr_n1079, csr_n1078, csr_n1077, csr_n1076, csr_n1075,
         csr_n1074, csr_n1073, csr_n1072, csr_n1071, csr_n1070, csr_n1069,
         csr_n1068, csr_n1067, csr_n1066, csr_n1065, csr_n1064, csr_n1063,
         csr_n1061, csr_n1060, csr_n1059, csr_n1058, csr_n1057, csr_n1056,
         csr_n1055, csr_n1054, csr_n1053, csr_n1052, csr_n1051, csr_n1050,
         csr_n1049, csr_n1048, csr_n1047, csr_n1046, csr_n1045, csr_n1044,
         csr_n1043, csr_n1042, csr_n1040, csr_n1039, csr_n1038, csr_n1037,
         csr_n1036, csr_n1035, csr_n1034, csr_n1033, csr_n1032, csr_n1031,
         csr_n1030, csr_n1029, csr_n1028, csr_n1027, csr_n1026, csr_n1025,
         csr_n1024, csr_n1023, csr_n1022, csr_n1021, csr_n1020, csr_n1019,
         csr_n1018, csr_n1017, csr_n1016, csr_n1015, csr_n1014, csr_n1013,
         csr_n1012, csr_n1011, csr_n1010, csr_n1009, csr_n1008, csr_n1007,
         csr_n1006, csr_n1005, csr_n1004, csr_n1003, csr_n1002, csr_n1001,
         csr_n1000, csr_n999, csr_n998, csr_n997, csr_n996, csr_n995, csr_n994,
         csr_n993, csr_n992, csr_n991, csr_n990, csr_n989, csr_n988, csr_n987,
         csr_n986, csr_n985, csr_n984, csr_n983, csr_n982, csr_n981, csr_n980,
         csr_n979, csr_n978, csr_n977, csr_n976, csr_n975, csr_n974, csr_n973,
         csr_n972, csr_n971, csr_n970, csr_n969, csr_n968, csr_n967, csr_n966,
         csr_n965, csr_n964, csr_n963, csr_n962, csr_n961, csr_n960, csr_n959,
         csr_n958, csr_n957, csr_n956, csr_n955, csr_n954, csr_n953, csr_n952,
         csr_n951, csr_n950, csr_n949, csr_n948, csr_n947, csr_n946, csr_n945,
         csr_n944, csr_n943, csr_n942, csr_n941, csr_n940, csr_n939, csr_n938,
         csr_n937, csr_n936, csr_n935, csr_n934, csr_n933, csr_n932, csr_n931,
         csr_n930, csr_n929, csr_n928, csr_n927, csr_n926, csr_n925, csr_n924,
         csr_n923, csr_n922, csr_n921, csr_n920, csr_n919, csr_n918, csr_n917,
         csr_n916, csr_n915, csr_n914, csr_n913, csr_n912, csr_n911, csr_n910,
         csr_n909, csr_n908, csr_n907, csr_n906, csr_n905, csr_n904, csr_n903,
         csr_n902, csr_n901, csr_n900, csr_n899, csr_n898, csr_n897, csr_n896,
         csr_n895, csr_n894, csr_n893, csr_n892, csr_n891, csr_n890, csr_n889,
         csr_n888, csr_n887, csr_n886, csr_n885, csr_n884, csr_n883, csr_n882,
         csr_n881, csr_n880, csr_n879, csr_n878, csr_n877, csr_n876, csr_n875,
         csr_n874, csr_n873, csr_n872, csr_n871, csr_n870, csr_n869, csr_n868,
         csr_n867, csr_n866, csr_n865, csr_n864, csr_n863, csr_n862, csr_n861,
         csr_n859, csr_n858, csr_n857, csr_n856, csr_n855, csr_n854, csr_n853,
         csr_n852, csr_n851, csr_n850, csr_n849, csr_n848, csr_n847, csr_n846,
         csr_n845, csr_n844, csr_n843, csr_n842, csr_n841, csr_n840, csr_n839,
         csr_n838, csr_n837, csr_n836, csr_n835, csr_n834, csr_n833, csr_n832,
         csr_n831, csr_n830, csr_n829, csr_n828, csr_n827, csr_n826, csr_n825,
         csr_n824, csr_n823, csr_n822, csr_n821, csr_n820, csr_n819, csr_n818,
         csr_n817, csr_n816, csr_n815, csr_n814, csr_n813, csr_n812, csr_n811,
         csr_n810, csr_n809, csr_n808, csr_n807, csr_n806, csr_n805, csr_n804,
         csr_n803, csr_n802, csr_n801, csr_n800, csr_n799, csr_n798, csr_n797,
         csr_n796, csr_n795, csr_n794, csr_n793, csr_n792, csr_n791, csr_n790,
         csr_n789, csr_n788, csr_n787, csr_n786, csr_n785, csr_n784, csr_n783,
         csr_n782, csr_n781, csr_n780, csr_n779, csr_n778, csr_n777, csr_n776,
         csr_n775, csr_n774, csr_n773, csr_n772, csr_n771, csr_n770, csr_n769,
         csr_n768, csr_n767, csr_n766, csr_n765, csr_n764, csr_n763, csr_n762,
         csr_n761, csr_n760, csr_n759, csr_n758, csr_n757, csr_n756, csr_n755,
         csr_n754, csr_n753, csr_n752, csr_n751, csr_n750, csr_n749, csr_n748,
         csr_n747, csr_n746, csr_n745, csr_n744, csr_n743, csr_n742, csr_n741,
         csr_n740, csr_n739, csr_n738, csr_n737, csr_n736, csr_n735, csr_n734,
         csr_n733, csr_n732, csr_n731, csr_n730, csr_n729, csr_n728, csr_n727,
         csr_n726, csr_n725, csr_n724, csr_n723, csr_n722, csr_n721, csr_n720,
         csr_n719, csr_n718, csr_n717, csr_n716, csr_n715, csr_n714, csr_n713,
         csr_n712, csr_n711, csr_n710, csr_n709, csr_n708, csr_n707, csr_n706,
         csr_n705, csr_n704, csr_n703, csr_n702, csr_n701, csr_n700, csr_n699,
         csr_n698, csr_n697, csr_n696, csr_n695, csr_n694, csr_n693, csr_n692,
         csr_n691, csr_n690, csr_n689, csr_n688, csr_n687, csr_n686, csr_n685,
         csr_n684, csr_n683, csr_n682, csr_n681, csr_n680, csr_n679, csr_n678,
         csr_n677, csr_n676, csr_n675, csr_n674, csr_n673, csr_n672, csr_n671,
         csr_n670, csr_n669, csr_n668, csr_n667, csr_n666, csr_n665, csr_n664,
         csr_n663, csr_n662, csr_n661, csr_n660, csr_n657, csr_n656, csr_n655,
         csr_n654, csr_n653, csr_n652, csr_n651, csr_n650, csr_n649, csr_n648,
         csr_n647, csr_n646, csr_n645, csr_n644, csr_n643, csr_n642, csr_n641,
         csr_n640, csr_n639, csr_n638, csr_n637, csr_n636, csr_n635, csr_n634,
         csr_n633, csr_n632, csr_n631, csr_n630, csr_n629, csr_n628, csr_n627,
         csr_n626, csr_n625, csr_n624, csr_n623, csr_n622, csr_n621, csr_n620,
         csr_n619, csr_n618, csr_n617, csr_n616, csr_n615, csr_n614, csr_n613,
         csr_n612, csr_n611, csr_n610, csr_n609, csr_n608, csr_n607, csr_n606,
         csr_n605, csr_n604, csr_n603, csr_n602, csr_n601, csr_n600, csr_n599,
         csr_n598, csr_n597, csr_n596, csr_n595, csr_n594, csr_n593, csr_n592,
         csr_n591, csr_n590, csr_n589, csr_n588, csr_n587, csr_n586, csr_n585,
         csr_n584, csr_n583, csr_n582, csr_n581, csr_n580, csr_n579, csr_n578,
         csr_n577, csr_n576, csr_n575, csr_n574, csr_n573, csr_n572, csr_n571,
         csr_n570, csr_n569, csr_n568, csr_n567, csr_n566, csr_n565, csr_n564,
         csr_n563, csr_n562, csr_n561, csr_n560, csr_n559, csr_n558, csr_n557,
         csr_n556, csr_n555, csr_n554, csr_n553, csr_n552, csr_n551, csr_n550,
         csr_n549, csr_n548, csr_n547, csr_n546, csr_n545, csr_n544, csr_n543,
         csr_n542, csr_n541, csr_n540, csr_n539, csr_n538, csr_n537, csr_n536,
         csr_n535, csr_n534, csr_n533, csr_n532, csr_n531, csr_n530, csr_n529,
         csr_n528, csr_n527, csr_n526, csr_n525, csr_n524, csr_n523, csr_n522,
         csr_n521, csr_n520, csr_n519, csr_n518, csr_n517, csr_n516, csr_n515,
         csr_n514, csr_n513, csr_n512, csr_n511, csr_n510, csr_n509, csr_n508,
         csr_n507, csr_n506, csr_n505, csr_n504, csr_n503, csr_n502, csr_n501,
         csr_n500, csr_n499, csr_n498, csr_n497, csr_n496, csr_n495, csr_n494,
         csr_n493, csr_n492, csr_n491, csr_n490, csr_n489, csr_n488, csr_n487,
         csr_n486, csr_n485, csr_n484, csr_n483, csr_n482, csr_n481, csr_n480,
         csr_n479, csr_n478, csr_n477, csr_n476, csr_n475, csr_n474, csr_n473,
         csr_n472, csr_n471, csr_n470, csr_n469, csr_n468, csr_n467, csr_n466,
         csr_n465, csr_n464, csr_n463, csr_n462, csr_n461, csr_n460, csr_n459,
         csr_n458, csr_n457, csr_n456, csr_n455, csr_n454, csr_n453, csr_n452,
         csr_n451, csr_n450, csr_n449, csr_n448, csr_n447, csr_n446, csr_n445,
         csr_n444, csr_n443, csr_n442, csr_n441, csr_n440, csr_n439, csr_n438,
         csr_n437, csr_n436, csr_n435, csr_n434, csr_n433, csr_n432, csr_n431,
         csr_n430, csr_n429, csr_n428, csr_n427, csr_n426, csr_n425, csr_n424,
         csr_n423, csr_n422, csr_n421, csr_n420, csr_n419, csr_n418, csr_n417,
         csr_n416, csr_n415, csr_n414, csr_n413, csr_n412, csr_n411, csr_n410,
         csr_n409, csr_n408, csr_n407, csr_n406, csr_n405, csr_n404, csr_n403,
         csr_n402, csr_n401, csr_n400, csr_n399, csr_n398, csr_n397, csr_n396,
         csr_n395, csr_n394, csr_n393, csr_n392, csr_n391, csr_n389, csr_n388,
         csr_n387, csr_n386, csr_n385, csr_n384, csr_n383, csr_n382, csr_n381,
         csr_n380, csr_n379, csr_n378, csr_n376, csr_n375, csr_n374, csr_n373,
         csr_n372, csr_n371, csr_n370, csr_n369, csr_n368, csr_n367, csr_n366,
         csr_n365, csr_n361, csr_n360, csr_n359, csr_n358, csr_n357, csr_n356,
         csr_n355, csr_n354, csr_n353, csr_n352, csr_n351, csr_n350, csr_n349,
         csr_n348, csr_n347, csr_n346, csr_n345, csr_n344, csr_n343, csr_n342,
         csr_n341, csr_n340, csr_n339, csr_n338, csr_n337, csr_n336, csr_n334,
         csr_n333, csr_n332, csr_n331, csr_n330, csr_n329, csr_n328, csr_n327,
         csr_n326, csr_n325, csr_n324, csr_n323, csr_n322, csr_n321, csr_n320,
         csr_n319, csr_n318, csr_n317, csr_n316, csr_n315, csr_n314, csr_n313,
         csr_n312, csr_n311, csr_n310, csr_n309, csr_n308, csr_n307, csr_n306,
         csr_n305, csr_n304, csr_n303, csr_n302, csr_n301, csr_n300, csr_n299,
         csr_n298, csr_n297, csr_n296, csr_n295, csr_n294, csr_n293, csr_n292,
         csr_n291, csr_n290, csr_n289, csr_n288, csr_n286, csr_n285, csr_n284,
         csr_n283, csr_n282, csr_n281, csr_n280, csr_n278, csr_n277, csr_n276,
         csr_n275, csr_n274, csr_n273, csr_n272, csr_n271, csr_n270, csr_n269,
         csr_n268, csr_n267, csr_n265, csr_n264, csr_n263, csr_n262, csr_n261,
         csr_n260, csr_n259, csr_n258, csr_n256, csr_n255, csr_n254, csr_n253,
         csr_n252, csr_n251, csr_n250, csr_n249, csr_n248, csr_n247, csr_n246,
         csr_n245, csr_n244, csr_n242, csr_n241, csr_n240, csr_n239, csr_n238,
         csr_n237, csr_n236, csr_n235, csr_n234, csr_n233, csr_n232, csr_n231,
         csr_n230, csr_n228, csr_n227, csr_n226, csr_n225, csr_n224, csr_n223,
         csr_n222, csr_n221, csr_n220, csr_n219, csr_n218, csr_n217, csr_n216,
         csr_n215, csr_n214, csr_n213, csr_n212, csr_n211, csr_n210, csr_n209,
         csr_n208, csr_n207, csr_n206, csr_n205, csr_n204, csr_n203, csr_n202,
         csr_n201, csr_n196, csr_n195, csr_n193, csr_n192, csr_n191, csr_n190,
         csr_n189, csr_n188, csr_n187, csr_n186, csr_n185, csr_n184, csr_n183,
         csr_n182, csr_n181, csr_n180, csr_n178, csr_n177, csr_n176, csr_n175,
         csr_n174, csr_n173, csr_n172, csr_n171, csr_n170, csr_n169, csr_n168,
         csr_n167, csr_n166, csr_n164, csr_n163, csr_n162, csr_n161, csr_n160,
         csr_n159, csr_n158, csr_n157, csr_n156, csr_n155, csr_n154, csr_n153,
         csr_n152, csr_n151, csr_n150, csr_n149, csr_n148, csr_n147, csr_n146,
         csr_n145, csr_n143, csr_n142, csr_n141, csr_n140, csr_n139, csr_n138,
         csr_n137, csr_n136, csr_n135, csr_n134, csr_n133, csr_n132, csr_n131,
         csr_n130, csr_n129, csr_n128, csr_n127, csr_n126, csr_n125, csr_n124,
         csr_n123, csr_n122, csr_n121, csr_n120, csr_n119, csr_n118, csr_n117,
         csr_n116, csr_n115, csr_n114, csr_n113, csr_n112, csr_n111, csr_n110,
         csr_n109, csr_n108, csr_n107, csr_n106, csr_n105, csr_n104, csr_n103,
         csr_n102, csr_n101, csr_n100, csr_n99, csr_n98, csr_n97, csr_n96,
         csr_n95, csr_n94, csr_n93, csr_n92, csr_n91, csr_n90, csr_n88,
         csr_n87, csr_n86, csr_n85, csr_n84, csr_n83, csr_n82, csr_n81,
         csr_n80, csr_n79, csr_n78, csr_n77, csr_n76, csr_n75, csr_n74,
         csr_n72, csr_n71, csr_n70, csr_n69, csr_n68, csr_n67, csr_n66,
         csr_n65, csr_n64, csr_n63, csr_n62, csr_n61, csr_n60, csr_n59,
         csr_n58, csr_n57, csr_n56, csr_n55, csr_n54, csr_n53, csr_n52,
         csr_n50, csr_n49, csr_n48, csr_n47, csr_n46, csr_n45, csr_n44,
         csr_n43, csr_n42, csr_n41, csr_n40, csr_n39, csr_n38, csr_n37,
         csr_n36, csr_n35, csr_n33, csr_n32, csr_n31, csr_n30, csr_n29,
         csr_n28, csr_n27, csr_n25, csr_n24, csr_n23, csr_n22, csr_n21,
         csr_n20, csr_n19, csr_n18, csr_n17, csr_n15, csr_n14, csr_n13,
         csr_n12, csr_n11, csr_n10, csr_n9, csr_n8, csr_n7, csr_n6, csr_n5,
         csr_n3, csr_n2, csr_n1, csr_n2169, csr_n2168, csr_n2167, csr_n2166,
         csr_n2165, csr_n2163, csr_n2162, csr_n2161, csr_n2160, csr_n2157,
         csr_n2156, csr_n2155, csr_n1346, csr_n1062, csr_n1041, csr_n860,
         csr_n659, csr_n658, csr_n200, csr_n199, csr_n194, csr_n51,
         csr_net35324, csr_net35319, csr_net35314, csr_net35309, csr_net35304,
         csr_net35301, csr_net35298, csr_net35295, csr_net35292, csr_net35289,
         csr_net35286, csr_net35283, csr_net35280, csr_net35277, csr_net35274,
         csr_net35271, csr_net35268, csr_net35265, csr_net35262, csr_net35259,
         csr_net35256, csr_net35253, csr_net35250, csr_net35247, csr_net35244,
         csr_net35241, csr_net35238, csr_net35235, csr_net35232, csr_net35229,
         csr_net35226, csr_net35223, csr_net35220, csr_net35217, csr_net35214,
         csr_net35211, csr_net35208, csr_net35205, csr_net35202, csr_net35199,
         csr_net35196, csr_net35193, csr_net35190, csr_net35187, csr_net35183,
         csr_net35177, csr_net35172, csr_net35167, csr_net35162, csr_net35157,
         csr_net35152, csr_net35147, csr_net35137, csr_net35132, csr_net35127,
         csr_net35122, csr_net35117, csr_net35112, csr_net35107, csr_net35102,
         csr_net35097, csr_net35092, csr_net35087, csr_net35082, csr_net35079,
         csr_net35076, csr_net35073, csr_net35070, csr_net35067, csr_net35064,
         csr_net35061, csr_net35058, csr_net35055, csr_net35052, csr_net35049,
         csr_net35046, csr_net35043, csr_net35040, csr_net35037, csr_net35034,
         csr_net35031, csr_net35028, csr_net35025, csr_net35022, csr_net35019,
         csr_net35016, csr_net35013, csr_net35010, csr_net35007, csr_net35004,
         csr_net35001, csr_net34998, csr_net34995, csr_net34992, csr_net34989,
         csr_net34986, csr_net34983, csr_net34980, csr_net34977, csr_net34974,
         csr_net34971, csr_net34968, csr_net34965, csr_net34961, csr_net34955,
         csr_net34950, csr_net34945, csr_net34940, csr_net34935, csr_net34930,
         csr_net34925, csr_net34920, csr_net34915, csr_net34910, csr_net34905,
         csr_net34900, csr_net34895, csr_net34890, csr_net34885, csr_net34880,
         csr_net34877, csr_net34874, csr_net34871, csr_net34868, csr_net34865,
         csr_net34862, csr_net34859, csr_net34856, csr_net34853, csr_net34850,
         csr_net34847, csr_net34844, csr_net34841, csr_net34838, csr_net34835,
         csr_net34832, csr_net34829, csr_net34826, csr_net34823, csr_net34820,
         csr_net34817, csr_net34814, csr_net34811, csr_net34808, csr_net34805,
         csr_net34802, csr_net34799, csr_net34796, csr_net34793, csr_net34790,
         csr_net34787, csr_net34784, csr_net34781, csr_net34778, csr_net34775,
         csr_net34772, csr_net34769, csr_net34766, csr_net34763, csr_net34759,
         csr_net34753, csr_net34748, csr_net34743, csr_net34738, csr_net34733,
         csr_net34728, csr_net34722, csr_N1948, csr_N1947, csr_N1946,
         csr_N1945, csr_N1944, csr_N1943, csr_N1942, csr_N1941, csr_N1940,
         csr_N1939, csr_N1938, csr_N1937, csr_N1936, csr_N1935, csr_N1934,
         csr_N1933, csr_N1932, csr_N1931, csr_N1930, csr_N1929, csr_N1928,
         csr_N1927, csr_N1926, csr_N1925, csr_N1924, csr_N1923, csr_N1922,
         csr_N1921, csr_N1920, csr_N1919, csr_N1918, csr_N1917, csr_N1916,
         csr_N1915, csr_N1914, csr_N1913, csr_N1912, csr_N1911, csr_N1910,
         csr_N1909, csr_N1908, csr_N1907, csr_N1906, csr_N1905, csr_N1904,
         csr_N1903, csr_N1902, csr_N1901, csr_N1900, csr_N1899, csr_N1898,
         csr_N1897, csr_N1896, csr_N1895, csr_N1894, csr_N1893, csr_N1892,
         csr_N1891, csr_N1890, csr_N1827, csr_N1826, csr_N1825, csr_N1824,
         csr_N1823, csr_N1822, csr_N1821, csr_N1693, csr_N1692, csr_N1691,
         csr_N1622, csr_N1582, csr_N1579, csr_N1577, csr_N1567, csr_N1558,
         csr_N1554, csr_N1553, csr_N1552, csr_N1551, csr_N1550, csr_N1549,
         csr_N1548, csr_N1547, csr_N1546, csr_N1545, csr_N1544, csr_N1543,
         csr_N1542, csr_N1541, csr_N1540, csr_N1539, csr_N1538, csr_N1537,
         csr_N1536, csr_N1535, csr_N1534, csr_N1533, csr_N1532, csr_N1531,
         csr_N1530, csr_N1529, csr_N1528, csr_N1527, csr_N1526, csr_N1525,
         csr_N1524, csr_N1523, csr_N1522, csr_N1521, csr_N1520, csr_N1519,
         csr_N1518, csr_N1517, csr_N1516, csr_N1515, csr_N1514, csr_N1513,
         csr_N1512, csr_N1511, csr_N1510, csr_N1509, csr_N1508, csr_N1507,
         csr_N1506, csr_N1505, csr_N1504, csr_N1503, csr_N1502, csr_N1501,
         csr_N1500, csr_N1499, csr_N1498, csr_N1497, csr_N1496, csr_N1433,
         csr_N1432, csr_N1431, csr_N1430, csr_N1429, csr_N1428, csr_N1426,
         csr_N1422, csr_N1421, csr_N1420, csr_N1419, csr_N1418, csr_N1417,
         csr_N1416, csr_N1415, csr_N1414, csr_N1413, csr_N1412, csr_N1411,
         csr_N1410, csr_N1409, csr_N1408, csr_N1407, csr_N1406, csr_N1405,
         csr_N1404, csr_N1403, csr_N1402, csr_N1401, csr_N1400, csr_N1399,
         csr_N1398, csr_N1397, csr_N1396, csr_N1395, csr_N1394, csr_N1393,
         csr_N1392, csr_N1391, csr_N1390, csr_N1389, csr_N1388, csr_N1387,
         csr_N1386, csr_N1385, csr_N1384, csr_N1383, csr_N1382, csr_N1381,
         csr_N1333, csr_N1274, csr_N1273, csr_N1272, csr_N1271, csr_N1270,
         csr_N1269, csr_N1033, csr_N1032, csr_N1031, csr_N1030, csr_N1029,
         csr_N1028, csr_N1027, csr_N1026, csr_N1025, csr_N1024, csr_N1023,
         csr_N1022, csr_N1021, csr_N1020, csr_N1019, csr_N1018, csr_N1017,
         csr_N1016, csr_N1015, csr_N1014, csr_N1013, csr_N1012, csr_N1011,
         csr_N1010, csr_N1009, csr_N1008, csr_N1007, csr_N1006, csr_N1005,
         csr_N1004, csr_N1003, csr_N1002, csr_N1001, csr_N1000, csr_N999,
         csr_N998, csr_N997, csr_N996, csr_N995, csr_N994, csr_N993, csr_N992,
         csr_N944, csr_N884, csr_N883, csr_N882, csr_N881, csr_N880, csr_N670,
         csr_N617, csr_N615, csr_N613, csr_N611, csr_N609, csr_N607, csr_N604,
         csr_N595, csr_N592, csr_N587, csr_N580, csr_N575, csr_N568, csr_N559,
         csr_N556, csr_N551, csr_N542, csr_N539, csr_N531, csr_N527, csr_N518,
         csr_N515, csr_N487, csr_N485, csr_N479, csr_N475, csr_N469, csr_N467,
         csr_N460, csr_N459, csr_N438, csr_N435, csr_N360, csr_N335, csr_N334,
         csr_N333, csr_N290, csr_N276, csr_n_T_3694_9_, csr_n_T_3678_63_,
         csr_wdata_0_, csr_wdata_1_, csr_wdata_2_, csr_wdata_3_, csr_wdata_4_,
         csr_wdata_5_, csr_wdata_6_, csr_wdata_7_, csr_wdata_8_, csr_wdata_9_,
         csr_wdata_10_, csr_wdata_11_, csr_wdata_12_, csr_wdata_13_,
         csr_wdata_14_, csr_wdata_15_, csr_wdata_16_, csr_wdata_17_,
         csr_wdata_18_, csr_wdata_19_, csr_wdata_20_, csr_wdata_21_,
         csr_wdata_22_, csr_wdata_23_, csr_wdata_24_, csr_wdata_25_,
         csr_wdata_26_, csr_wdata_27_, csr_wdata_28_, csr_wdata_29_,
         csr_wdata_30_, csr_wdata_31_, csr_wdata_32_, csr_wdata_33_,
         csr_wdata_34_, csr_wdata_35_, csr_wdata_36_, csr_wdata_37_,
         csr_wdata_38_, csr_wdata_39_, csr_wdata_40_, csr_wdata_41_,
         csr_wdata_42_, csr_wdata_43_, csr_wdata_44_, csr_wdata_45_,
         csr_wdata_46_, csr_wdata_47_, csr_wdata_48_, csr_wdata_49_,
         csr_wdata_50_, csr_wdata_51_, csr_wdata_52_, csr_wdata_53_,
         csr_wdata_54_, csr_wdata_55_, csr_wdata_56_, csr_wdata_57_,
         csr_wdata_58_, csr_wdata_59_, csr_wdata_60_, csr_wdata_61_,
         csr_wdata_62_, csr_wdata_63_, csr_reg_sepc_1_, csr_reg_sepc_2_,
         csr_reg_sepc_3_, csr_reg_sepc_4_, csr_reg_sepc_5_, csr_reg_sepc_6_,
         csr_reg_sepc_7_, csr_reg_sepc_8_, csr_reg_sepc_9_, csr_reg_sepc_10_,
         csr_reg_sepc_11_, csr_reg_sepc_12_, csr_reg_sepc_13_,
         csr_reg_sepc_14_, csr_reg_sepc_15_, csr_reg_sepc_16_,
         csr_reg_sepc_17_, csr_reg_sepc_18_, csr_reg_sepc_19_,
         csr_reg_sepc_20_, csr_reg_sepc_21_, csr_reg_sepc_22_,
         csr_reg_sepc_23_, csr_reg_sepc_24_, csr_reg_sepc_25_,
         csr_reg_sepc_26_, csr_reg_sepc_27_, csr_reg_sepc_28_,
         csr_reg_sepc_29_, csr_reg_sepc_30_, csr_reg_sepc_31_,
         csr_reg_sepc_32_, csr_reg_sepc_33_, csr_reg_sepc_34_,
         csr_reg_sepc_35_, csr_reg_sepc_36_, csr_reg_sepc_37_,
         csr_reg_sepc_38_, csr_reg_sepc_39_, csr_read_fcsr_0_,
         csr_read_fcsr_1_, csr_read_fcsr_2_, csr_read_fcsr_3_,
         csr_read_fcsr_4_, csr_reg_dpc_1_, csr_reg_dpc_2_, csr_reg_dpc_3_,
         csr_reg_dpc_4_, csr_reg_dpc_5_, csr_reg_dpc_6_, csr_reg_dpc_7_,
         csr_reg_dpc_8_, csr_reg_dpc_9_, csr_reg_dpc_10_, csr_reg_dpc_11_,
         csr_reg_dpc_12_, csr_reg_dpc_13_, csr_reg_dpc_14_, csr_reg_dpc_15_,
         csr_reg_dpc_16_, csr_reg_dpc_17_, csr_reg_dpc_18_, csr_reg_dpc_19_,
         csr_reg_dpc_20_, csr_reg_dpc_21_, csr_reg_dpc_22_, csr_reg_dpc_23_,
         csr_reg_dpc_24_, csr_reg_dpc_25_, csr_reg_dpc_26_, csr_reg_dpc_27_,
         csr_reg_dpc_28_, csr_reg_dpc_29_, csr_reg_dpc_30_, csr_reg_dpc_31_,
         csr_reg_dpc_32_, csr_reg_dpc_33_, csr_reg_dpc_34_, csr_reg_dpc_35_,
         csr_reg_dpc_36_, csr_reg_dpc_37_, csr_reg_dpc_38_, csr_reg_dpc_39_,
         csr_n_T_389_0, csr_n_T_389_1, csr_n_T_389_2, csr_reg_mepc_1_,
         csr_reg_mepc_2_, csr_reg_mepc_3_, csr_reg_mepc_4_, csr_reg_mepc_5_,
         csr_reg_mepc_6_, csr_reg_mepc_7_, csr_reg_mepc_8_, csr_reg_mepc_9_,
         csr_reg_mepc_10_, csr_reg_mepc_11_, csr_reg_mepc_12_,
         csr_reg_mepc_13_, csr_reg_mepc_14_, csr_reg_mepc_15_,
         csr_reg_mepc_16_, csr_reg_mepc_17_, csr_reg_mepc_18_,
         csr_reg_mepc_19_, csr_reg_mepc_20_, csr_reg_mepc_21_,
         csr_reg_mepc_22_, csr_reg_mepc_23_, csr_reg_mepc_24_,
         csr_reg_mepc_25_, csr_reg_mepc_26_, csr_reg_mepc_27_,
         csr_reg_mepc_28_, csr_reg_mepc_29_, csr_reg_mepc_30_,
         csr_reg_mepc_31_, csr_reg_mepc_32_, csr_reg_mepc_33_,
         csr_reg_mepc_34_, csr_reg_mepc_35_, csr_reg_mepc_36_,
         csr_reg_mepc_37_, csr_reg_mepc_38_, csr_reg_mepc_39_, csr_n_T_366_59_,
         csr_reg_stvec_2_, csr_reg_stvec_3_, csr_reg_stvec_4_,
         csr_reg_stvec_5_, csr_reg_stvec_6_, csr_reg_stvec_7_,
         csr_reg_stvec_8_, csr_reg_stvec_9_, csr_reg_stvec_10_,
         csr_reg_stvec_11_, csr_reg_stvec_12_, csr_reg_stvec_13_,
         csr_reg_stvec_14_, csr_reg_stvec_15_, csr_reg_stvec_16_,
         csr_reg_stvec_17_, csr_reg_stvec_18_, csr_reg_stvec_19_,
         csr_reg_stvec_20_, csr_reg_stvec_21_, csr_reg_stvec_22_,
         csr_reg_stvec_23_, csr_reg_stvec_24_, csr_reg_stvec_25_,
         csr_reg_stvec_26_, csr_reg_stvec_27_, csr_reg_stvec_28_,
         csr_reg_stvec_29_, csr_reg_stvec_30_, csr_reg_stvec_31_,
         csr_reg_stvec_32_, csr_reg_stvec_33_, csr_reg_stvec_34_,
         csr_reg_stvec_35_, csr_reg_stvec_36_, csr_reg_stvec_37_,
         csr_reg_stvec_38_, csr_reg_mtvec_2_, csr_reg_mtvec_3_,
         csr_reg_mtvec_4_, csr_reg_mtvec_5_, csr_reg_mtvec_6_,
         csr_reg_mtvec_7_, csr_reg_mtvec_8_, csr_reg_mtvec_9_,
         csr_reg_mtvec_10_, csr_reg_mtvec_11_, csr_reg_mtvec_12_,
         csr_reg_mtvec_13_, csr_reg_mtvec_14_, csr_reg_mtvec_15_,
         csr_reg_mtvec_16_, csr_reg_mtvec_17_, csr_reg_mtvec_18_,
         csr_reg_mtvec_19_, csr_reg_mtvec_20_, csr_reg_mtvec_21_,
         csr_reg_mtvec_22_, csr_reg_mtvec_23_, csr_reg_mtvec_24_,
         csr_reg_mtvec_25_, csr_reg_mtvec_26_, csr_reg_mtvec_27_,
         csr_reg_mtvec_28_, csr_reg_mtvec_29_, csr_reg_mtvec_30_,
         csr_reg_mtvec_31_, csr_reg_mie_1_, csr_reg_mie_3_, csr_reg_mie_5_,
         csr_reg_mie_7_, csr_reg_mie_9_, csr_reg_mie_11_, csr_n_T_61_1,
         csr_n_T_61_5_, csr_n_T_45_0_, csr_n_T_45_1_, csr_n_T_45_2_,
         csr_n_T_45_3_, csr_n_T_45_4_, csr_n_T_45_5_, csr_n_T_45_6_,
         csr_n_T_45_7_, csr_n_T_45_8_, csr_n_T_45_9_, csr_n_T_45_10_,
         csr_n_T_45_11_, csr_n_T_45_12_, csr_n_T_45_13_, csr_n_T_45_14_,
         csr_n_T_45_15_, csr_n_T_45_16_, csr_n_T_45_17_, csr_n_T_45_18_,
         csr_n_T_45_19_, csr_n_T_45_20_, csr_n_T_45_21_, csr_n_T_45_22_,
         csr_n_T_45_23_, csr_n_T_45_24_, csr_n_T_45_25_, csr_n_T_45_26_,
         csr_n_T_45_27_, csr_n_T_45_28_, csr_n_T_45_29_, csr_n_T_45_30_,
         csr_n_T_45_31_, csr_n_T_45_32_, csr_n_T_45_33_, csr_n_T_45_34_,
         csr_n_T_45_35_, csr_n_T_45_36_, csr_n_T_45_37_, csr_n_T_45_38_,
         csr_n_T_45_39_, csr_n_T_45_40_, csr_n_T_45_41_, csr_n_T_45_42_,
         csr_n_T_45_43_, csr_n_T_45_44_, csr_n_T_45_45_, csr_n_T_45_46_,
         csr_n_T_45_47_, csr_n_T_45_48_, csr_n_T_45_49_, csr_n_T_45_50_,
         csr_n_T_45_51_, csr_n_T_45_52_, csr_n_T_45_53_, csr_n_T_45_54_,
         csr_n_T_45_55_, csr_n_T_45_56_, csr_n_T_45_57_, csr_n_T_45_58_,
         csr_n_T_45_59_, csr_n_T_45_60_, csr_n_T_45_61_, csr_n_T_45_62_,
         csr_n_T_45_63_, csr_read_scounteren_0_, csr_read_scounteren_1_,
         csr_read_scounteren_2_, csr_read_mcounteren_0_,
         csr_read_mcounteren_1_, csr_read_mcounteren_2_, csr_read_medeleg_0,
         csr_read_medeleg_2_, csr_read_medeleg_3_, csr_read_medeleg_4_,
         csr_read_medeleg_6, csr_read_medeleg_8, csr_read_medeleg_12,
         csr_read_medeleg_13, csr_read_medeleg_15, csr_read_mideleg_1,
         csr_read_mideleg_5, csr_read_mideleg_9_, csr_n_T_1155_0_,
         csr_n_T_1155_1_, csr_n_T_1155_3, csr_n1967, csr_n1966, csr_n1965,
         csr_n1964, csr_n1963, csr_n1962, csr_n1961, csr_n1960, csr_n1959,
         csr_n1958, csr_n1957, csr_n1956, csr_n1955, csr_n1954, csr_n1953,
         csr_n1952, csr_n1951, csr_n1950, csr_n1949, csr_n1948, csr_n1947,
         csr_n1946, csr_n1945, csr_n1944, csr_n1943, csr_n1942, csr_n1941,
         csr_n1940, csr_n1939, csr_n1938, csr_n1937, csr_n1936, csr_n1935,
         csr_n1934, csr_n1933, csr_n1932, csr_n1931, csr_n_1930_, csr_n_1929_,
         csr_n1928, csr_n1927, csr_n1926, csr_n1925, csr_n1924,
         csr_io_status_isa_0_, csr_n1923, csr_n1922, csr_io_status_isa_12_,
         csr_n1921, csr_n1920, csr_n1919, csr_n1918, csr_io_status_debug,
         csr_add_x_427_n199, csr_add_x_427_n198, csr_add_x_427_n197,
         csr_add_x_427_n196, csr_add_x_427_n195, csr_add_x_427_n194,
         csr_add_x_427_n193, csr_add_x_427_n192, csr_add_x_427_n191,
         csr_add_x_427_n190, csr_add_x_427_n189, csr_add_x_427_n188,
         csr_add_x_427_n187, csr_add_x_427_n186, csr_add_x_427_n185,
         csr_add_x_427_n184, csr_add_x_427_n183, csr_add_x_427_n182,
         csr_add_x_427_n181, csr_add_x_427_n180, csr_add_x_427_n179,
         csr_add_x_427_n178, csr_add_x_427_n177, csr_add_x_427_n176,
         csr_add_x_427_n175, csr_add_x_427_n174, csr_add_x_427_n173,
         csr_add_x_427_n172, csr_add_x_427_n171, csr_add_x_427_n170,
         csr_add_x_427_n169, csr_add_x_427_n168, csr_add_x_427_n167,
         csr_add_x_427_n166, csr_add_x_427_n165, csr_add_x_427_n164,
         csr_add_x_427_n163, csr_add_x_427_n162, csr_add_x_427_n161,
         csr_add_x_427_n160, csr_add_x_427_n159, csr_add_x_427_n93,
         csr_add_x_426_n199, csr_add_x_426_n198, csr_add_x_426_n197,
         csr_add_x_426_n196, csr_add_x_426_n195, csr_add_x_426_n194,
         csr_add_x_426_n193, csr_add_x_426_n192, csr_add_x_426_n191,
         csr_add_x_426_n190, csr_add_x_426_n189, csr_add_x_426_n188,
         csr_add_x_426_n187, csr_add_x_426_n186, csr_add_x_426_n185,
         csr_add_x_426_n184, csr_add_x_426_n183, csr_add_x_426_n182,
         csr_add_x_426_n181, csr_add_x_426_n180, csr_add_x_426_n179,
         csr_add_x_426_n178, csr_add_x_426_n177, csr_add_x_426_n176,
         csr_add_x_426_n175, csr_add_x_426_n174, csr_add_x_426_n173,
         csr_add_x_426_n172, csr_add_x_426_n171, csr_add_x_426_n170,
         csr_add_x_426_n169, csr_add_x_426_n168, csr_add_x_426_n167,
         csr_add_x_426_n166, csr_add_x_426_n165, csr_add_x_426_n164,
         csr_add_x_426_n163, csr_add_x_426_n162, csr_add_x_426_n161,
         csr_add_x_426_n160, csr_add_x_426_n159, csr_add_x_426_n93,
         csr_add_x_425_n199, csr_add_x_425_n198, csr_add_x_425_n197,
         csr_add_x_425_n196, csr_add_x_425_n195, csr_add_x_425_n194,
         csr_add_x_425_n193, csr_add_x_425_n192, csr_add_x_425_n191,
         csr_add_x_425_n190, csr_add_x_425_n189, csr_add_x_425_n188,
         csr_add_x_425_n187, csr_add_x_425_n186, csr_add_x_425_n185,
         csr_add_x_425_n184, csr_add_x_425_n183, csr_add_x_425_n182,
         csr_add_x_425_n181, csr_add_x_425_n180, csr_add_x_425_n179,
         csr_add_x_425_n178, csr_add_x_425_n177, csr_add_x_425_n176,
         csr_add_x_425_n175, csr_add_x_425_n174, csr_add_x_425_n173,
         csr_add_x_425_n172, csr_add_x_425_n171, csr_add_x_425_n170,
         csr_add_x_425_n169, csr_add_x_425_n168, csr_add_x_425_n167,
         csr_add_x_425_n166, csr_add_x_425_n165, csr_add_x_425_n164,
         csr_add_x_425_n163, csr_add_x_425_n162, csr_add_x_425_n161,
         csr_add_x_425_n160, csr_add_x_425_n159, csr_add_x_425_n93,
         csr_add_x_424_n199, csr_add_x_424_n198, csr_add_x_424_n197,
         csr_add_x_424_n196, csr_add_x_424_n195, csr_add_x_424_n194,
         csr_add_x_424_n193, csr_add_x_424_n192, csr_add_x_424_n191,
         csr_add_x_424_n190, csr_add_x_424_n189, csr_add_x_424_n188,
         csr_add_x_424_n187, csr_add_x_424_n186, csr_add_x_424_n185,
         csr_add_x_424_n184, csr_add_x_424_n183, csr_add_x_424_n182,
         csr_add_x_424_n181, csr_add_x_424_n180, csr_add_x_424_n179,
         csr_add_x_424_n178, csr_add_x_424_n177, csr_add_x_424_n176,
         csr_add_x_424_n175, csr_add_x_424_n174, csr_add_x_424_n173,
         csr_add_x_424_n172, csr_add_x_424_n171, csr_add_x_424_n170,
         csr_add_x_424_n169, csr_add_x_424_n168, csr_add_x_424_n167,
         csr_add_x_424_n166, csr_add_x_424_n165, csr_add_x_424_n164,
         csr_add_x_424_n163, csr_add_x_424_n162, csr_add_x_424_n161,
         csr_add_x_424_n160, csr_add_x_424_n159, csr_add_x_424_n93,
         csr_add_x_423_n199, csr_add_x_423_n198, csr_add_x_423_n197,
         csr_add_x_423_n196, csr_add_x_423_n195, csr_add_x_423_n194,
         csr_add_x_423_n193, csr_add_x_423_n192, csr_add_x_423_n191,
         csr_add_x_423_n190, csr_add_x_423_n189, csr_add_x_423_n188,
         csr_add_x_423_n187, csr_add_x_423_n186, csr_add_x_423_n185,
         csr_add_x_423_n184, csr_add_x_423_n183, csr_add_x_423_n182,
         csr_add_x_423_n181, csr_add_x_423_n180, csr_add_x_423_n179,
         csr_add_x_423_n178, csr_add_x_423_n177, csr_add_x_423_n176,
         csr_add_x_423_n175, csr_add_x_423_n174, csr_add_x_423_n173,
         csr_add_x_423_n172, csr_add_x_423_n171, csr_add_x_423_n170,
         csr_add_x_423_n169, csr_add_x_423_n168, csr_add_x_423_n167,
         csr_add_x_423_n166, csr_add_x_423_n165, csr_add_x_423_n164,
         csr_add_x_423_n163, csr_add_x_423_n162, csr_add_x_423_n161,
         csr_add_x_423_n160, csr_add_x_423_n159, csr_add_x_423_n93,
         csr_add_x_422_n199, csr_add_x_422_n198, csr_add_x_422_n197,
         csr_add_x_422_n196, csr_add_x_422_n195, csr_add_x_422_n194,
         csr_add_x_422_n193, csr_add_x_422_n192, csr_add_x_422_n191,
         csr_add_x_422_n190, csr_add_x_422_n189, csr_add_x_422_n188,
         csr_add_x_422_n187, csr_add_x_422_n186, csr_add_x_422_n185,
         csr_add_x_422_n184, csr_add_x_422_n183, csr_add_x_422_n182,
         csr_add_x_422_n181, csr_add_x_422_n180, csr_add_x_422_n179,
         csr_add_x_422_n178, csr_add_x_422_n177, csr_add_x_422_n176,
         csr_add_x_422_n175, csr_add_x_422_n174, csr_add_x_422_n173,
         csr_add_x_422_n172, csr_add_x_422_n171, csr_add_x_422_n170,
         csr_add_x_422_n169, csr_add_x_422_n168, csr_add_x_422_n167,
         csr_add_x_422_n166, csr_add_x_422_n165, csr_add_x_422_n164,
         csr_add_x_422_n163, csr_add_x_422_n162, csr_add_x_422_n161,
         csr_add_x_422_n160, csr_add_x_422_n159, csr_add_x_422_n93,
         csr_add_x_421_n199, csr_add_x_421_n198, csr_add_x_421_n197,
         csr_add_x_421_n196, csr_add_x_421_n195, csr_add_x_421_n194,
         csr_add_x_421_n193, csr_add_x_421_n192, csr_add_x_421_n191,
         csr_add_x_421_n190, csr_add_x_421_n189, csr_add_x_421_n188,
         csr_add_x_421_n187, csr_add_x_421_n186, csr_add_x_421_n185,
         csr_add_x_421_n184, csr_add_x_421_n183, csr_add_x_421_n182,
         csr_add_x_421_n181, csr_add_x_421_n180, csr_add_x_421_n179,
         csr_add_x_421_n178, csr_add_x_421_n177, csr_add_x_421_n176,
         csr_add_x_421_n175, csr_add_x_421_n174, csr_add_x_421_n173,
         csr_add_x_421_n172, csr_add_x_421_n171, csr_add_x_421_n170,
         csr_add_x_421_n169, csr_add_x_421_n168, csr_add_x_421_n167,
         csr_add_x_421_n166, csr_add_x_421_n165, csr_add_x_421_n164,
         csr_add_x_421_n163, csr_add_x_421_n162, csr_add_x_421_n161,
         csr_add_x_421_n160, csr_add_x_421_n159, csr_add_x_421_n93,
         csr_add_x_420_n199, csr_add_x_420_n198, csr_add_x_420_n197,
         csr_add_x_420_n196, csr_add_x_420_n195, csr_add_x_420_n194,
         csr_add_x_420_n193, csr_add_x_420_n192, csr_add_x_420_n191,
         csr_add_x_420_n190, csr_add_x_420_n189, csr_add_x_420_n188,
         csr_add_x_420_n187, csr_add_x_420_n186, csr_add_x_420_n185,
         csr_add_x_420_n184, csr_add_x_420_n183, csr_add_x_420_n182,
         csr_add_x_420_n181, csr_add_x_420_n180, csr_add_x_420_n179,
         csr_add_x_420_n178, csr_add_x_420_n177, csr_add_x_420_n176,
         csr_add_x_420_n175, csr_add_x_420_n174, csr_add_x_420_n173,
         csr_add_x_420_n172, csr_add_x_420_n171, csr_add_x_420_n170,
         csr_add_x_420_n169, csr_add_x_420_n168, csr_add_x_420_n167,
         csr_add_x_420_n166, csr_add_x_420_n165, csr_add_x_420_n164,
         csr_add_x_420_n163, csr_add_x_420_n162, csr_add_x_420_n161,
         csr_add_x_420_n160, csr_add_x_420_n159, csr_add_x_420_n93,
         csr_add_x_381_n411, csr_add_x_381_n410, csr_add_x_381_n409,
         csr_add_x_381_n408, csr_add_x_381_n407, csr_add_x_381_n406,
         csr_add_x_381_n405, csr_add_x_381_n404, csr_add_x_381_n403,
         csr_add_x_381_n402, csr_add_x_381_n401, csr_add_x_381_n400,
         csr_add_x_381_n399, csr_add_x_381_n398, csr_add_x_381_n397,
         csr_add_x_381_n396, csr_add_x_381_n395, csr_add_x_381_n394,
         csr_add_x_381_n393, csr_add_x_381_n392, csr_add_x_381_n391,
         csr_add_x_381_n390, csr_add_x_381_n389, csr_add_x_381_n388,
         csr_add_x_381_n387, csr_add_x_381_n386, csr_add_x_381_n385,
         csr_add_x_381_n384, csr_add_x_381_n383, csr_add_x_381_n382,
         csr_add_x_381_n381, csr_add_x_381_n380, csr_add_x_381_n379,
         csr_add_x_381_n378, csr_add_x_381_n377, csr_add_x_381_n376,
         csr_add_x_381_n375, csr_add_x_381_n374, csr_add_x_381_n373,
         csr_add_x_381_n372, csr_add_x_381_n371, csr_add_x_381_n370,
         csr_add_x_381_n369, csr_add_x_381_n368, csr_add_x_381_n367,
         csr_add_x_381_n366, csr_add_x_381_n365, csr_add_x_381_n364,
         csr_add_x_381_n363, csr_add_x_381_n362, csr_add_x_381_n361,
         csr_add_x_381_n360, csr_add_x_381_n359, csr_add_x_381_n358,
         csr_add_x_381_n357, csr_add_x_381_n356, csr_add_x_381_n355,
         csr_add_x_381_n354, csr_add_x_381_n353, csr_add_x_381_n352,
         csr_add_x_381_n351, csr_add_x_381_n350, csr_add_x_381_n349,
         csr_add_x_381_n348, csr_add_x_381_n347, csr_add_x_381_n346,
         csr_add_x_381_n345, csr_add_x_381_n344, csr_add_x_381_n343,
         csr_add_x_381_n342, csr_add_x_381_n341, csr_add_x_381_n340,
         csr_add_x_381_n339, csr_add_x_381_n338, csr_add_x_381_n337,
         csr_add_x_381_n336, csr_add_x_381_n335, csr_add_x_381_n334,
         csr_add_x_381_n333, csr_add_x_381_n332, csr_add_x_381_n331,
         csr_add_x_381_n330, csr_add_x_381_n329, csr_add_x_381_n328,
         csr_add_x_381_n327, csr_add_x_381_n326, csr_add_x_381_n325,
         csr_add_x_381_n203, csr_add_x_379_n411, csr_add_x_379_n410,
         csr_add_x_379_n409, csr_add_x_379_n408, csr_add_x_379_n407,
         csr_add_x_379_n406, csr_add_x_379_n405, csr_add_x_379_n404,
         csr_add_x_379_n403, csr_add_x_379_n402, csr_add_x_379_n401,
         csr_add_x_379_n400, csr_add_x_379_n399, csr_add_x_379_n398,
         csr_add_x_379_n397, csr_add_x_379_n396, csr_add_x_379_n395,
         csr_add_x_379_n394, csr_add_x_379_n393, csr_add_x_379_n392,
         csr_add_x_379_n391, csr_add_x_379_n390, csr_add_x_379_n389,
         csr_add_x_379_n388, csr_add_x_379_n387, csr_add_x_379_n386,
         csr_add_x_379_n385, csr_add_x_379_n384, csr_add_x_379_n383,
         csr_add_x_379_n382, csr_add_x_379_n381, csr_add_x_379_n380,
         csr_add_x_379_n379, csr_add_x_379_n378, csr_add_x_379_n377,
         csr_add_x_379_n376, csr_add_x_379_n375, csr_add_x_379_n374,
         csr_add_x_379_n373, csr_add_x_379_n372, csr_add_x_379_n371,
         csr_add_x_379_n370, csr_add_x_379_n369, csr_add_x_379_n368,
         csr_add_x_379_n367, csr_add_x_379_n366, csr_add_x_379_n365,
         csr_add_x_379_n364, csr_add_x_379_n363, csr_add_x_379_n362,
         csr_add_x_379_n361, csr_add_x_379_n360, csr_add_x_379_n359,
         csr_add_x_379_n358, csr_add_x_379_n357, csr_add_x_379_n356,
         csr_add_x_379_n355, csr_add_x_379_n354, csr_add_x_379_n353,
         csr_add_x_379_n352, csr_add_x_379_n351, csr_add_x_379_n350,
         csr_add_x_379_n349, csr_add_x_379_n348, csr_add_x_379_n347,
         csr_add_x_379_n346, csr_add_x_379_n345, csr_add_x_379_n344,
         csr_add_x_379_n343, csr_add_x_379_n342, csr_add_x_379_n341,
         csr_add_x_379_n340, csr_add_x_379_n339, csr_add_x_379_n338,
         csr_add_x_379_n337, csr_add_x_379_n336, csr_add_x_379_n335,
         csr_add_x_379_n334, csr_add_x_379_n333, csr_add_x_379_n332,
         csr_add_x_379_n331, csr_add_x_379_n330, csr_add_x_379_n329,
         csr_add_x_379_n328, csr_add_x_379_n327, csr_add_x_379_n326,
         csr_add_x_379_n325, csr_add_x_379_n203, bpu_n166, bpu_n165, bpu_n164,
         bpu_n163, bpu_n162, bpu_n161, bpu_n160, bpu_n159, bpu_n156, bpu_n155,
         bpu_n154, bpu_n153, bpu_n152, bpu_n151, bpu_n150, bpu_n149, bpu_n148,
         bpu_n147, bpu_n146, bpu_n145, bpu_n144, bpu_n143, bpu_n142, bpu_n141,
         bpu_n140, bpu_n139, bpu_n138, bpu_n137, bpu_n136, bpu_n135, bpu_n134,
         bpu_n133, bpu_n132, bpu_n131, bpu_n130, bpu_n129, bpu_n128, bpu_n127,
         bpu_n126, bpu_n125, bpu_n124, bpu_n123, bpu_n122, bpu_n121, bpu_n120,
         bpu_n119, bpu_n118, bpu_n117, bpu_n116, bpu_n115, bpu_n114, bpu_n113,
         bpu_n112, bpu_n111, bpu_n110, bpu_n109, bpu_n108, bpu_n107, bpu_n106,
         bpu_n105, bpu_n104, bpu_n103, bpu_n102, bpu_n101, bpu_n100, bpu_n99,
         bpu_n98, bpu_n97, bpu_n96, bpu_n95, bpu_n94, bpu_n93, bpu_n92,
         bpu_n91, bpu_n90, bpu_n89, bpu_n88, bpu_n87, bpu_n86, bpu_n85,
         bpu_n84, bpu_n83, bpu_n82, bpu_n81, bpu_n80, bpu_n79, bpu_n78,
         bpu_n77, bpu_n76, bpu_n75, bpu_n74, bpu_n73, bpu_n72, bpu_n71,
         bpu_n70, bpu_n69, bpu_n68, bpu_n67, bpu_n66, bpu_n65, bpu_n64,
         bpu_n63, bpu_n62, bpu_n61, bpu_n60, bpu_n59, bpu_n58, bpu_n57,
         bpu_n56, bpu_n55, bpu_n54, bpu_n53, bpu_n52, bpu_n51, bpu_n50,
         bpu_n49, bpu_n48, bpu_n47, bpu_n46, bpu_n45, bpu_n44, bpu_n43,
         bpu_n42, bpu_n41, bpu_n40, bpu_n39, bpu_n38, bpu_n37, bpu_n36,
         bpu_n35, bpu_n34, bpu_n33, bpu_n32, bpu_n31, bpu_n30, bpu_n29,
         bpu_n28, bpu_n27, bpu_n26, bpu_n25, bpu_n24, bpu_n23, bpu_n22,
         bpu_n21, bpu_n20, bpu_n19, bpu_n18, bpu_n17, bpu_n16, bpu_n15,
         bpu_n14, bpu_n13, bpu_n12, bpu_n11, bpu_n10, bpu_n9, bpu_n8, bpu_n7,
         bpu_n6, bpu_n5, bpu_n4, bpu_n3, bpu_n2, bpu_n1, bpu_n_T_73, bpu_n_T_9,
         bpu_gte_x_5_n422, bpu_gte_x_5_n421, bpu_gte_x_5_n420,
         bpu_gte_x_5_n419, bpu_gte_x_5_n418, bpu_gte_x_5_n417,
         bpu_gte_x_5_n416, bpu_gte_x_5_n415, bpu_gte_x_5_n414,
         bpu_gte_x_5_n413, bpu_gte_x_5_n412, bpu_gte_x_5_n411,
         bpu_gte_x_5_n410, bpu_gte_x_5_n409, bpu_gte_x_5_n408,
         bpu_gte_x_5_n407, bpu_gte_x_5_n406, bpu_gte_x_5_n405,
         bpu_gte_x_5_n404, bpu_gte_x_5_n403, bpu_gte_x_5_n402,
         bpu_gte_x_5_n401, bpu_gte_x_5_n400, bpu_gte_x_5_n399,
         bpu_gte_x_5_n398, bpu_gte_x_5_n397, bpu_gte_x_5_n396,
         bpu_gte_x_5_n395, bpu_gte_x_5_n394, bpu_gte_x_5_n393,
         bpu_gte_x_5_n392, bpu_gte_x_5_n391, bpu_gte_x_5_n390,
         bpu_gte_x_5_n389, bpu_gte_x_5_n388, bpu_gte_x_5_n387,
         bpu_gte_x_5_n386, bpu_gte_x_5_n385, bpu_gte_x_5_n384,
         bpu_gte_x_5_n383, bpu_gte_x_5_n382, bpu_gte_x_5_n381,
         bpu_gte_x_5_n380, bpu_gte_x_5_n379, bpu_gte_x_5_n378,
         bpu_gte_x_5_n377, bpu_gte_x_5_n376, bpu_gte_x_5_n375,
         bpu_gte_x_5_n374, bpu_gte_x_5_n373, bpu_gte_x_5_n372,
         bpu_gte_x_5_n371, bpu_gte_x_5_n370, bpu_gte_x_5_n369,
         bpu_gte_x_5_n368, bpu_gte_x_5_n367, bpu_gte_x_5_n366,
         bpu_gte_x_5_n365, bpu_gte_x_5_n364, bpu_gte_x_5_n363,
         bpu_gte_x_5_n362, bpu_gte_x_5_n361, bpu_gte_x_5_n360,
         bpu_gte_x_5_n359, bpu_gte_x_5_n358, bpu_gte_x_5_n357,
         bpu_gte_x_5_n356, bpu_gte_x_5_n355, bpu_gte_x_5_n354,
         bpu_gte_x_5_n353, bpu_gte_x_5_n352, bpu_gte_x_5_n351,
         bpu_gte_x_5_n350, bpu_gte_x_5_n349, bpu_gte_x_5_n348,
         bpu_gte_x_5_n347, bpu_gte_x_5_n346, bpu_gte_x_5_n345,
         bpu_gte_x_5_n344, bpu_gte_x_5_n343, bpu_gte_x_5_n342,
         bpu_gte_x_5_n341, bpu_gte_x_5_n340, bpu_gte_x_5_n339,
         bpu_gte_x_5_n338, bpu_gte_x_5_n337, bpu_gte_x_5_n336,
         bpu_gte_x_5_n335, bpu_gte_x_5_n334, bpu_gte_x_5_n333,
         bpu_gte_x_5_n331, bpu_gte_x_5_n330, bpu_gte_x_5_n329,
         bpu_gte_x_5_n328, bpu_gte_x_5_n327, bpu_gte_x_5_n326,
         bpu_gte_x_5_n325, bpu_gte_x_5_n324, bpu_gte_x_5_n323,
         bpu_gte_x_5_n322, bpu_gte_x_5_n321, bpu_gte_x_5_n320,
         bpu_gte_x_5_n318, bpu_gte_x_5_n317, bpu_gte_x_5_n316,
         bpu_gte_x_5_n315, bpu_gte_x_5_n314, bpu_gte_x_5_n313,
         bpu_gte_x_5_n312, bpu_gte_x_5_n311, bpu_gte_x_5_n310,
         bpu_gte_x_5_n309, bpu_gte_x_5_n308, bpu_gte_x_5_n307,
         bpu_gte_x_5_n306, bpu_gte_x_5_n305, bpu_gte_x_5_n304,
         bpu_gte_x_5_n303, bpu_gte_x_5_n302, bpu_gte_x_5_n301,
         bpu_gte_x_5_n300, bpu_gte_x_5_n299, bpu_gte_x_5_n298,
         bpu_gte_x_5_n296, bpu_gte_x_5_n295, bpu_gte_x_5_n294,
         bpu_gte_x_5_n293, bpu_gte_x_5_n292, bpu_gte_x_5_n291,
         bpu_gte_x_5_n290, bpu_gte_x_5_n289, bpu_gte_x_5_n288,
         bpu_gte_x_5_n287, bpu_gte_x_5_n286, bpu_gte_x_5_n285,
         bpu_gte_x_5_n284, bpu_gte_x_2_n423, bpu_gte_x_2_n422,
         bpu_gte_x_2_n421, bpu_gte_x_2_n420, bpu_gte_x_2_n419,
         bpu_gte_x_2_n418, bpu_gte_x_2_n417, bpu_gte_x_2_n416,
         bpu_gte_x_2_n415, bpu_gte_x_2_n414, bpu_gte_x_2_n413,
         bpu_gte_x_2_n412, bpu_gte_x_2_n411, bpu_gte_x_2_n410,
         bpu_gte_x_2_n409, bpu_gte_x_2_n408, bpu_gte_x_2_n407,
         bpu_gte_x_2_n406, bpu_gte_x_2_n405, bpu_gte_x_2_n404,
         bpu_gte_x_2_n403, bpu_gte_x_2_n402, bpu_gte_x_2_n401,
         bpu_gte_x_2_n400, bpu_gte_x_2_n399, bpu_gte_x_2_n398,
         bpu_gte_x_2_n397, bpu_gte_x_2_n396, bpu_gte_x_2_n395,
         bpu_gte_x_2_n394, bpu_gte_x_2_n393, bpu_gte_x_2_n392,
         bpu_gte_x_2_n391, bpu_gte_x_2_n390, bpu_gte_x_2_n389,
         bpu_gte_x_2_n388, bpu_gte_x_2_n387, bpu_gte_x_2_n386,
         bpu_gte_x_2_n385, bpu_gte_x_2_n384, bpu_gte_x_2_n383,
         bpu_gte_x_2_n382, bpu_gte_x_2_n381, bpu_gte_x_2_n380,
         bpu_gte_x_2_n379, bpu_gte_x_2_n378, bpu_gte_x_2_n377,
         bpu_gte_x_2_n376, bpu_gte_x_2_n375, bpu_gte_x_2_n374,
         bpu_gte_x_2_n373, bpu_gte_x_2_n372, bpu_gte_x_2_n371,
         bpu_gte_x_2_n370, bpu_gte_x_2_n369, bpu_gte_x_2_n368,
         bpu_gte_x_2_n367, bpu_gte_x_2_n366, bpu_gte_x_2_n365,
         bpu_gte_x_2_n364, bpu_gte_x_2_n363, bpu_gte_x_2_n362,
         bpu_gte_x_2_n361, bpu_gte_x_2_n360, bpu_gte_x_2_n359,
         bpu_gte_x_2_n358, bpu_gte_x_2_n357, bpu_gte_x_2_n356,
         bpu_gte_x_2_n355, bpu_gte_x_2_n354, bpu_gte_x_2_n353,
         bpu_gte_x_2_n352, bpu_gte_x_2_n351, bpu_gte_x_2_n350,
         bpu_gte_x_2_n349, bpu_gte_x_2_n348, bpu_gte_x_2_n347,
         bpu_gte_x_2_n346, bpu_gte_x_2_n345, bpu_gte_x_2_n344,
         bpu_gte_x_2_n343, bpu_gte_x_2_n342, bpu_gte_x_2_n341,
         bpu_gte_x_2_n340, bpu_gte_x_2_n339, bpu_gte_x_2_n338,
         bpu_gte_x_2_n337, bpu_gte_x_2_n336, bpu_gte_x_2_n335,
         bpu_gte_x_2_n334, bpu_gte_x_2_n333, bpu_gte_x_2_n332,
         bpu_gte_x_2_n331, bpu_gte_x_2_n330, bpu_gte_x_2_n329,
         bpu_gte_x_2_n328, bpu_gte_x_2_n327, bpu_gte_x_2_n326,
         bpu_gte_x_2_n325, bpu_gte_x_2_n324, bpu_gte_x_2_n323,
         bpu_gte_x_2_n322, bpu_gte_x_2_n321, bpu_gte_x_2_n320,
         bpu_gte_x_2_n319, bpu_gte_x_2_n318, bpu_gte_x_2_n317,
         bpu_gte_x_2_n316, bpu_gte_x_2_n315, bpu_gte_x_2_n314,
         bpu_gte_x_2_n313, bpu_gte_x_2_n312, bpu_gte_x_2_n311,
         bpu_gte_x_2_n310, bpu_gte_x_2_n309, bpu_gte_x_2_n308,
         bpu_gte_x_2_n307, bpu_gte_x_2_n306, bpu_gte_x_2_n305,
         bpu_gte_x_2_n304, bpu_gte_x_2_n303, bpu_gte_x_2_n302,
         bpu_gte_x_2_n300, bpu_gte_x_2_n299, bpu_gte_x_2_n297,
         bpu_gte_x_2_n296, bpu_gte_x_2_n295, bpu_gte_x_2_n294,
         bpu_gte_x_2_n293, bpu_gte_x_2_n292, bpu_gte_x_2_n291,
         bpu_gte_x_2_n290, bpu_gte_x_2_n289, bpu_gte_x_2_n288,
         bpu_gte_x_2_n287, bpu_gte_x_2_n286, bpu_gte_x_2_n285,
         bpu_gte_x_2_n284, alu_SYNOPSYS_UNCONNECTED_1, alu_n606, alu_n605,
         alu_n604, alu_n603, alu_n602, alu_n601, alu_n600, alu_n599, alu_n598,
         alu_n597, alu_n596, alu_n595, alu_n594, alu_n593, alu_n592, alu_n591,
         alu_n590, alu_n589, alu_n588, alu_n587, alu_n586, alu_n585, alu_n584,
         alu_n583, alu_n582, alu_n581, alu_n580, alu_n579, alu_n578, alu_n577,
         alu_n576, alu_n575, alu_n574, alu_n573, alu_n572, alu_n571, alu_n570,
         alu_n569, alu_n568, alu_n567, alu_n566, alu_n565, alu_n564, alu_n563,
         alu_n562, alu_n561, alu_n560, alu_n559, alu_n558, alu_n557, alu_n556,
         alu_n555, alu_n554, alu_n553, alu_n552, alu_n551, alu_n550, alu_n549,
         alu_n548, alu_n547, alu_n546, alu_n545, alu_n544, alu_n543, alu_n542,
         alu_n541, alu_n540, alu_n539, alu_n538, alu_n537, alu_n536, alu_n535,
         alu_n534, alu_n533, alu_n532, alu_n531, alu_n530, alu_n529, alu_n528,
         alu_n527, alu_n526, alu_n525, alu_n524, alu_n523, alu_n522, alu_n521,
         alu_n520, alu_n519, alu_n518, alu_n517, alu_n516, alu_n515, alu_n514,
         alu_n513, alu_n512, alu_n511, alu_n510, alu_n509, alu_n508, alu_n507,
         alu_n506, alu_n505, alu_n504, alu_n503, alu_n502, alu_n501, alu_n500,
         alu_n499, alu_n498, alu_n497, alu_n496, alu_n495, alu_n494, alu_n493,
         alu_n492, alu_n491, alu_n490, alu_n489, alu_n488, alu_n487, alu_n486,
         alu_n485, alu_n484, alu_n483, alu_n482, alu_n481, alu_n480, alu_n479,
         alu_n478, alu_n477, alu_n476, alu_n475, alu_n474, alu_n473, alu_n472,
         alu_n471, alu_n470, alu_n469, alu_n468, alu_n467, alu_n466, alu_n465,
         alu_n464, alu_n463, alu_n462, alu_n461, alu_n460, alu_n459, alu_n458,
         alu_n457, alu_n456, alu_n455, alu_n454, alu_n453, alu_n452, alu_n451,
         alu_n450, alu_n449, alu_n448, alu_n447, alu_n446, alu_n445, alu_n444,
         alu_n443, alu_n442, alu_n441, alu_n440, alu_n439, alu_n438, alu_n437,
         alu_n436, alu_n435, alu_n434, alu_n433, alu_n432, alu_n431, alu_n430,
         alu_n429, alu_n428, alu_n427, alu_n426, alu_n425, alu_n424, alu_n423,
         alu_n422, alu_n421, alu_n420, alu_n419, alu_n418, alu_n417, alu_n416,
         alu_n415, alu_n414, alu_n413, alu_n412, alu_n411, alu_n410, alu_n409,
         alu_n408, alu_n407, alu_n406, alu_n405, alu_n404, alu_n403, alu_n402,
         alu_n401, alu_n400, alu_n399, alu_n398, alu_n397, alu_n396, alu_n395,
         alu_n394, alu_n393, alu_n392, alu_n391, alu_n390, alu_n389, alu_n388,
         alu_n387, alu_n386, alu_n385, alu_n384, alu_n383, alu_n382, alu_n381,
         alu_n380, alu_n379, alu_n378, alu_n377, alu_n376, alu_n375, alu_n374,
         alu_n373, alu_n372, alu_n371, alu_n370, alu_n369, alu_n368, alu_n367,
         alu_n366, alu_n365, alu_n364, alu_n363, alu_n362, alu_n361, alu_n360,
         alu_n359, alu_n358, alu_n357, alu_n356, alu_n355, alu_n354, alu_n353,
         alu_n352, alu_n351, alu_n350, alu_n349, alu_n348, alu_n347, alu_n346,
         alu_n345, alu_n344, alu_n343, alu_n342, alu_n341, alu_n340, alu_n339,
         alu_n338, alu_n337, alu_n336, alu_n335, alu_n334, alu_n333, alu_n332,
         alu_n331, alu_n330, alu_n329, alu_n328, alu_n327, alu_n326, alu_n325,
         alu_n324, alu_n323, alu_n322, alu_n321, alu_n320, alu_n319, alu_n318,
         alu_n317, alu_n316, alu_n315, alu_n314, alu_n313, alu_n312, alu_n311,
         alu_n310, alu_n309, alu_n308, alu_n307, alu_n306, alu_n305, alu_n304,
         alu_n303, alu_n302, alu_n301, alu_n300, alu_n299, alu_n298, alu_n297,
         alu_n296, alu_n295, alu_n294, alu_n293, alu_n292, alu_n291, alu_n290,
         alu_n289, alu_n288, alu_n287, alu_n286, alu_n285, alu_n284, alu_n283,
         alu_n282, alu_n281, alu_n280, alu_n279, alu_n278, alu_n277, alu_n276,
         alu_n275, alu_n274, alu_n273, alu_n272, alu_n271, alu_n270, alu_n269,
         alu_n268, alu_n267, alu_n266, alu_n265, alu_n264, alu_n263, alu_n262,
         alu_n261, alu_n260, alu_n259, alu_n258, alu_n257, alu_n256, alu_n255,
         alu_n254, alu_n253, alu_n252, alu_n251, alu_n250, alu_n249, alu_n248,
         alu_n247, alu_n246, alu_n245, alu_n244, alu_n243, alu_n242, alu_n241,
         alu_n240, alu_n239, alu_n238, alu_n237, alu_n236, alu_n235, alu_n234,
         alu_n233, alu_n232, alu_n231, alu_n230, alu_n229, alu_n228, alu_n227,
         alu_n226, alu_n225, alu_n224, alu_n223, alu_n222, alu_n221, alu_n220,
         alu_n219, alu_n218, alu_n217, alu_n216, alu_n215, alu_n214, alu_n213,
         alu_n212, alu_n211, alu_n210, alu_n209, alu_n208, alu_n207, alu_n206,
         alu_n205, alu_n204, alu_n203, alu_n202, alu_n201, alu_n200, alu_n199,
         alu_n198, alu_n197, alu_n196, alu_n195, alu_n194, alu_n193, alu_n192,
         alu_n191, alu_n190, alu_n189, alu_n188, alu_n187, alu_n186, alu_n185,
         alu_n184, alu_n183, alu_n182, alu_n181, alu_n180, alu_n179, alu_n178,
         alu_n177, alu_n176, alu_n175, alu_n174, alu_n173, alu_n172, alu_n171,
         alu_n170, alu_n169, alu_n168, alu_n167, alu_n166, alu_n165, alu_n164,
         alu_n163, alu_n162, alu_n161, alu_n160, alu_n159, alu_n158, alu_n157,
         alu_n156, alu_n155, alu_n154, alu_n153, alu_n152, alu_n151, alu_n150,
         alu_n149, alu_n148, alu_n147, alu_n146, alu_n145, alu_n144, alu_n143,
         alu_n142, alu_n141, alu_n140, alu_n139, alu_n138, alu_n137, alu_n136,
         alu_n135, alu_n134, alu_n133, alu_n132, alu_n131, alu_n130, alu_n129,
         alu_n128, alu_n127, alu_n126, alu_n125, alu_n124, alu_n123, alu_n122,
         alu_n121, alu_n120, alu_n119, alu_n118, alu_n117, alu_n116, alu_n115,
         alu_n114, alu_n113, alu_n112, alu_n111, alu_n110, alu_n109, alu_n108,
         alu_n107, alu_n106, alu_n105, alu_n104, alu_n103, alu_n102, alu_n101,
         alu_n100, alu_n99, alu_n98, alu_n97, alu_n96, alu_n95, alu_n94,
         alu_n93, alu_n92, alu_n91, alu_n90, alu_n89, alu_n88, alu_n87,
         alu_n86, alu_n85, alu_n84, alu_n83, alu_n82, alu_n81, alu_n80,
         alu_n79, alu_n78, alu_n77, alu_n76, alu_n75, alu_n74, alu_n73,
         alu_n72, alu_n71, alu_n70, alu_n69, alu_n68, alu_n67, alu_n66,
         alu_n65, alu_n64, alu_n63, alu_n62, alu_n61, alu_n60, alu_n59,
         alu_n58, alu_n57, alu_n56, alu_n55, alu_n54, alu_n53, alu_n52,
         alu_n51, alu_n50, alu_n49, alu_n48, alu_n47, alu_n46, alu_n45,
         alu_n43, alu_n42, alu_n41, alu_n40, alu_n39, alu_n38, alu_n37,
         alu_n36, alu_n35, alu_n34, alu_n33, alu_n32, alu_n31, alu_n30,
         alu_n29, alu_n28, alu_n27, alu_n26, alu_n25, alu_n24, alu_n23,
         alu_n22, alu_n21, alu_n20, alu_n19, alu_n18, alu_n17, alu_n16,
         alu_n15, alu_n14, alu_n13, alu_n12, alu_n11, alu_n10, alu_n9, alu_n8,
         alu_n7, alu_n6, alu_n5, alu_n4, alu_n3, alu_n2, alu_n1,
         alu_n_T_101_0_, alu_n_T_101_1_, alu_n_T_101_2_, alu_n_T_101_3_,
         alu_n_T_101_4_, alu_n_T_101_5_, alu_n_T_101_6_, alu_n_T_101_7_,
         alu_n_T_101_8_, alu_n_T_101_9_, alu_n_T_101_10_, alu_n_T_101_11_,
         alu_n_T_101_12_, alu_n_T_101_13_, alu_n_T_101_14_, alu_n_T_101_15_,
         alu_n_T_101_16_, alu_n_T_101_17_, alu_n_T_101_18_, alu_n_T_101_19_,
         alu_n_T_101_20_, alu_n_T_101_21_, alu_n_T_101_22_, alu_n_T_101_23_,
         alu_n_T_101_24_, alu_n_T_101_25_, alu_n_T_101_26_, alu_n_T_101_27_,
         alu_n_T_101_28_, alu_n_T_101_29_, alu_n_T_101_30_, alu_n_T_101_31_,
         alu_n_T_101_32_, alu_n_T_101_33_, alu_n_T_101_34_, alu_n_T_101_35_,
         alu_n_T_101_36_, alu_n_T_101_37_, alu_n_T_101_38_, alu_n_T_101_39_,
         alu_n_T_101_40_, alu_n_T_101_41_, alu_n_T_101_42_, alu_n_T_101_43_,
         alu_n_T_101_44_, alu_n_T_101_45_, alu_n_T_101_46_, alu_n_T_101_47_,
         alu_n_T_101_48_, alu_n_T_101_49_, alu_n_T_101_50_, alu_n_T_101_51_,
         alu_n_T_101_52_, alu_n_T_101_53_, alu_n_T_101_54_, alu_n_T_101_55_,
         alu_n_T_101_56_, alu_n_T_101_57_, alu_n_T_101_58_, alu_n_T_101_59_,
         alu_n_T_101_60_, alu_n_T_101_61_, alu_n_T_101_62_, alu_n_T_101_63_,
         alu_n_T_100_64_, alu_shin_0_, alu_shin_1_, alu_shin_2_, alu_shin_3_,
         alu_shin_4_, alu_shin_5_, alu_shin_6_, alu_shin_7_, alu_shin_8_,
         alu_shin_9_, alu_shin_10_, alu_shin_11_, alu_shin_12_, alu_shin_13_,
         alu_shin_14_, alu_shin_15_, alu_shin_16_, alu_shin_17_, alu_shin_18_,
         alu_shin_19_, alu_shin_20_, alu_shin_21_, alu_shin_22_, alu_shin_23_,
         alu_shin_24_, alu_shin_25_, alu_shin_26_, alu_shin_27_, alu_shin_28_,
         alu_shin_29_, alu_shin_30_, alu_shin_31_, alu_shin_32_, alu_shin_33_,
         alu_shin_34_, alu_shin_35_, alu_shin_36_, alu_shin_37_, alu_shin_38_,
         alu_shin_39_, alu_shin_40_, alu_shin_41_, alu_shin_42_, alu_shin_43_,
         alu_shin_44_, alu_shin_45_, alu_shin_46_, alu_shin_47_, alu_shin_48_,
         alu_shin_49_, alu_shin_50_, alu_shin_51_, alu_shin_52_, alu_shin_53_,
         alu_shin_54_, alu_shin_55_, alu_shin_56_, alu_shin_57_, alu_shin_58_,
         alu_shin_59_, alu_shin_60_, alu_shin_61_, alu_shin_62_, alu_shin_63_,
         alu_shamt_5_, alu_in2_inv_0_, alu_in2_inv_1_, alu_in2_inv_2_,
         alu_in2_inv_3_, alu_in2_inv_4_, alu_in2_inv_5_, alu_in2_inv_6_,
         alu_in2_inv_7_, alu_in2_inv_8_, alu_in2_inv_9_, alu_in2_inv_10_,
         alu_in2_inv_11_, alu_in2_inv_12_, alu_in2_inv_13_, alu_in2_inv_14_,
         alu_in2_inv_15_, alu_in2_inv_16_, alu_in2_inv_17_, alu_in2_inv_18_,
         alu_in2_inv_19_, alu_in2_inv_20_, alu_in2_inv_21_, alu_in2_inv_22_,
         alu_in2_inv_23_, alu_in2_inv_24_, alu_in2_inv_25_, alu_in2_inv_26_,
         alu_in2_inv_27_, alu_in2_inv_28_, alu_in2_inv_29_, alu_in2_inv_30_,
         alu_in2_inv_31_, alu_in2_inv_32_, alu_in2_inv_33_, alu_in2_inv_34_,
         alu_in2_inv_35_, alu_in2_inv_36_, alu_in2_inv_37_, alu_in2_inv_38_,
         alu_in2_inv_39_, alu_in2_inv_40_, alu_in2_inv_41_, alu_in2_inv_42_,
         alu_in2_inv_43_, alu_in2_inv_44_, alu_in2_inv_45_, alu_in2_inv_46_,
         alu_in2_inv_47_, alu_in2_inv_48_, alu_in2_inv_49_, alu_in2_inv_50_,
         alu_in2_inv_51_, alu_in2_inv_52_, alu_in2_inv_53_, alu_in2_inv_54_,
         alu_in2_inv_55_, alu_in2_inv_56_, alu_in2_inv_57_, alu_in2_inv_58_,
         alu_in2_inv_59_, alu_in2_inv_60_, alu_in2_inv_61_, alu_in2_inv_62_,
         alu_in2_inv_63_, alu_n630, alu_n629, alu_n628, alu_n627, alu_n626,
         alu_n625, alu_n624, alu_n623, alu_n622, alu_n621, alu_n620, alu_n619,
         alu_n618, alu_n617, alu_n616, alu_n615, alu_n614, alu_n613, alu_n612,
         alu_n611, alu_n610, alu_n609, alu_n608, alu_n607,
         alu_DP_OP_31J40_124_1870_n917, alu_DP_OP_31J40_124_1870_n916,
         alu_DP_OP_31J40_124_1870_n915, alu_DP_OP_31J40_124_1870_n914,
         alu_DP_OP_31J40_124_1870_n913, alu_DP_OP_31J40_124_1870_n912,
         alu_DP_OP_31J40_124_1870_n911, alu_DP_OP_31J40_124_1870_n910,
         alu_DP_OP_31J40_124_1870_n909, alu_DP_OP_31J40_124_1870_n908,
         alu_DP_OP_31J40_124_1870_n907, alu_DP_OP_31J40_124_1870_n906,
         alu_DP_OP_31J40_124_1870_n905, alu_DP_OP_31J40_124_1870_n904,
         alu_DP_OP_31J40_124_1870_n903, alu_DP_OP_31J40_124_1870_n902,
         alu_DP_OP_31J40_124_1870_n901, alu_DP_OP_31J40_124_1870_n900,
         alu_DP_OP_31J40_124_1870_n899, alu_DP_OP_31J40_124_1870_n898,
         alu_DP_OP_31J40_124_1870_n897, alu_DP_OP_31J40_124_1870_n896,
         alu_DP_OP_31J40_124_1870_n895, alu_DP_OP_31J40_124_1870_n894,
         alu_DP_OP_31J40_124_1870_n893, alu_DP_OP_31J40_124_1870_n892,
         alu_DP_OP_31J40_124_1870_n891, alu_DP_OP_31J40_124_1870_n890,
         alu_DP_OP_31J40_124_1870_n889, alu_DP_OP_31J40_124_1870_n888,
         alu_DP_OP_31J40_124_1870_n887, alu_DP_OP_31J40_124_1870_n886,
         alu_DP_OP_31J40_124_1870_n885, alu_DP_OP_31J40_124_1870_n884,
         alu_DP_OP_31J40_124_1870_n883, alu_DP_OP_31J40_124_1870_n882,
         alu_DP_OP_31J40_124_1870_n881, alu_DP_OP_31J40_124_1870_n880,
         alu_DP_OP_31J40_124_1870_n879, alu_DP_OP_31J40_124_1870_n878,
         alu_DP_OP_31J40_124_1870_n877, alu_DP_OP_31J40_124_1870_n876,
         alu_DP_OP_31J40_124_1870_n875, alu_DP_OP_31J40_124_1870_n874,
         alu_DP_OP_31J40_124_1870_n873, alu_DP_OP_31J40_124_1870_n872,
         alu_DP_OP_31J40_124_1870_n871, alu_DP_OP_31J40_124_1870_n870,
         alu_DP_OP_31J40_124_1870_n869, alu_DP_OP_31J40_124_1870_n868,
         alu_DP_OP_31J40_124_1870_n867, alu_DP_OP_31J40_124_1870_n866,
         alu_DP_OP_31J40_124_1870_n865, alu_DP_OP_31J40_124_1870_n864,
         alu_DP_OP_31J40_124_1870_n863, alu_DP_OP_31J40_124_1870_n862,
         alu_DP_OP_31J40_124_1870_n861, alu_DP_OP_31J40_124_1870_n860,
         alu_DP_OP_31J40_124_1870_n859, alu_DP_OP_31J40_124_1870_n858,
         alu_DP_OP_31J40_124_1870_n857, alu_DP_OP_31J40_124_1870_n856,
         alu_DP_OP_31J40_124_1870_n855, alu_DP_OP_31J40_124_1870_n854,
         alu_DP_OP_31J40_124_1870_n853, alu_DP_OP_31J40_124_1870_n852,
         alu_DP_OP_31J40_124_1870_n851, alu_DP_OP_31J40_124_1870_n850,
         alu_DP_OP_31J40_124_1870_n849, alu_DP_OP_31J40_124_1870_n848,
         alu_DP_OP_31J40_124_1870_n847, alu_DP_OP_31J40_124_1870_n846,
         alu_DP_OP_31J40_124_1870_n845, alu_DP_OP_31J40_124_1870_n844,
         alu_DP_OP_31J40_124_1870_n843, alu_DP_OP_31J40_124_1870_n842,
         alu_DP_OP_31J40_124_1870_n841, alu_DP_OP_31J40_124_1870_n840,
         alu_DP_OP_31J40_124_1870_n839, alu_DP_OP_31J40_124_1870_n838,
         alu_DP_OP_31J40_124_1870_n837, alu_DP_OP_31J40_124_1870_n836,
         alu_DP_OP_31J40_124_1870_n835, alu_DP_OP_31J40_124_1870_n834,
         alu_DP_OP_31J40_124_1870_n833, alu_DP_OP_31J40_124_1870_n832,
         alu_DP_OP_31J40_124_1870_n831, alu_DP_OP_31J40_124_1870_n830,
         alu_DP_OP_31J40_124_1870_n829, alu_DP_OP_31J40_124_1870_n828,
         alu_DP_OP_31J40_124_1870_n827, alu_DP_OP_31J40_124_1870_n826,
         alu_DP_OP_31J40_124_1870_n825, alu_DP_OP_31J40_124_1870_n824,
         alu_DP_OP_31J40_124_1870_n823, alu_DP_OP_31J40_124_1870_n822,
         alu_DP_OP_31J40_124_1870_n821, alu_DP_OP_31J40_124_1870_n820,
         alu_DP_OP_31J40_124_1870_n819, alu_DP_OP_31J40_124_1870_n818,
         alu_DP_OP_31J40_124_1870_n817, alu_DP_OP_31J40_124_1870_n816,
         alu_DP_OP_31J40_124_1870_n815, alu_DP_OP_31J40_124_1870_n814,
         alu_DP_OP_31J40_124_1870_n813, alu_DP_OP_31J40_124_1870_n812,
         alu_DP_OP_31J40_124_1870_n811, alu_DP_OP_31J40_124_1870_n810,
         alu_DP_OP_31J40_124_1870_n809, alu_DP_OP_31J40_124_1870_n808,
         alu_DP_OP_31J40_124_1870_n807, alu_DP_OP_31J40_124_1870_n806,
         alu_DP_OP_31J40_124_1870_n805, alu_DP_OP_31J40_124_1870_n804,
         alu_DP_OP_31J40_124_1870_n803, alu_DP_OP_31J40_124_1870_n802,
         alu_DP_OP_31J40_124_1870_n801, alu_DP_OP_31J40_124_1870_n800,
         alu_DP_OP_31J40_124_1870_n799, alu_DP_OP_31J40_124_1870_n798,
         alu_DP_OP_31J40_124_1870_n797, alu_DP_OP_31J40_124_1870_n796,
         alu_DP_OP_31J40_124_1870_n795, alu_DP_OP_31J40_124_1870_n794,
         alu_DP_OP_31J40_124_1870_n793, alu_DP_OP_31J40_124_1870_n792,
         alu_DP_OP_31J40_124_1870_n791, alu_DP_OP_31J40_124_1870_n790,
         alu_DP_OP_31J40_124_1870_n789, alu_DP_OP_31J40_124_1870_n788,
         alu_DP_OP_31J40_124_1870_n787, alu_DP_OP_31J40_124_1870_n786,
         alu_DP_OP_31J40_124_1870_n785, alu_DP_OP_31J40_124_1870_n784,
         alu_DP_OP_31J40_124_1870_n783, alu_DP_OP_31J40_124_1870_n782,
         alu_DP_OP_31J40_124_1870_n781, alu_DP_OP_31J40_124_1870_n780,
         alu_DP_OP_31J40_124_1870_n779, alu_DP_OP_31J40_124_1870_n778,
         alu_DP_OP_31J40_124_1870_n777, alu_DP_OP_31J40_124_1870_n776,
         alu_DP_OP_31J40_124_1870_n775, alu_DP_OP_31J40_124_1870_n774,
         alu_DP_OP_31J40_124_1870_n773, alu_DP_OP_31J40_124_1870_n772,
         alu_DP_OP_31J40_124_1870_n771, alu_DP_OP_31J40_124_1870_n770,
         alu_DP_OP_31J40_124_1870_n769, alu_DP_OP_31J40_124_1870_n768,
         alu_DP_OP_31J40_124_1870_n767, alu_DP_OP_31J40_124_1870_n766,
         alu_DP_OP_31J40_124_1870_n765, alu_DP_OP_31J40_124_1870_n764,
         alu_DP_OP_31J40_124_1870_n763, alu_DP_OP_31J40_124_1870_n762,
         alu_DP_OP_31J40_124_1870_n761, alu_DP_OP_31J40_124_1870_n760,
         alu_DP_OP_31J40_124_1870_n759, alu_DP_OP_31J40_124_1870_n758,
         alu_DP_OP_31J40_124_1870_n757, alu_DP_OP_31J40_124_1870_n756,
         alu_DP_OP_31J40_124_1870_n755, alu_DP_OP_31J40_124_1870_n754,
         alu_DP_OP_31J40_124_1870_n753, alu_DP_OP_31J40_124_1870_n752,
         alu_DP_OP_31J40_124_1870_n751, alu_DP_OP_31J40_124_1870_n750,
         alu_DP_OP_31J40_124_1870_n749, alu_DP_OP_31J40_124_1870_n748,
         alu_DP_OP_31J40_124_1870_n747, alu_DP_OP_31J40_124_1870_n746,
         alu_DP_OP_31J40_124_1870_n745, alu_DP_OP_31J40_124_1870_n744,
         alu_DP_OP_31J40_124_1870_n743, alu_DP_OP_31J40_124_1870_n742,
         alu_DP_OP_31J40_124_1870_n741, alu_DP_OP_31J40_124_1870_n740,
         alu_DP_OP_31J40_124_1870_n739, alu_DP_OP_31J40_124_1870_n738,
         alu_DP_OP_31J40_124_1870_n737, alu_DP_OP_31J40_124_1870_n736,
         alu_DP_OP_31J40_124_1870_n735, alu_DP_OP_31J40_124_1870_n734,
         alu_DP_OP_31J40_124_1870_n733, alu_DP_OP_31J40_124_1870_n732,
         alu_DP_OP_31J40_124_1870_n731, alu_DP_OP_31J40_124_1870_n730,
         alu_DP_OP_31J40_124_1870_n729, alu_DP_OP_31J40_124_1870_n728,
         alu_DP_OP_31J40_124_1870_n727, alu_DP_OP_31J40_124_1870_n726,
         alu_DP_OP_31J40_124_1870_n725, alu_DP_OP_31J40_124_1870_n724,
         alu_DP_OP_31J40_124_1870_n723, alu_DP_OP_31J40_124_1870_n722,
         alu_DP_OP_31J40_124_1870_n721, alu_DP_OP_31J40_124_1870_n720,
         alu_DP_OP_31J40_124_1870_n719, alu_DP_OP_31J40_124_1870_n718,
         alu_DP_OP_31J40_124_1870_n717, alu_DP_OP_31J40_124_1870_n716,
         alu_DP_OP_31J40_124_1870_n715, alu_DP_OP_31J40_124_1870_n714,
         alu_DP_OP_31J40_124_1870_n713, alu_DP_OP_31J40_124_1870_n712,
         alu_DP_OP_31J40_124_1870_n711, alu_DP_OP_31J40_124_1870_n710,
         alu_DP_OP_31J40_124_1870_n709, alu_DP_OP_31J40_124_1870_n708,
         alu_DP_OP_31J40_124_1870_n707, alu_DP_OP_31J40_124_1870_n706,
         alu_DP_OP_31J40_124_1870_n705, alu_DP_OP_31J40_124_1870_n704,
         alu_DP_OP_31J40_124_1870_n703, alu_DP_OP_31J40_124_1870_n442,
         alu_ashr_7_n841, alu_ashr_7_n840, alu_ashr_7_n839, alu_ashr_7_n838,
         alu_ashr_7_n837, alu_ashr_7_n836, alu_ashr_7_n835, alu_ashr_7_n834,
         alu_ashr_7_n833, alu_ashr_7_n832, alu_ashr_7_n831, alu_ashr_7_n830,
         alu_ashr_7_n829, alu_ashr_7_n828, alu_ashr_7_n827, alu_ashr_7_n826,
         alu_ashr_7_n825, alu_ashr_7_n824, alu_ashr_7_n823, alu_ashr_7_n822,
         alu_ashr_7_n821, alu_ashr_7_n820, alu_ashr_7_n819, alu_ashr_7_n818,
         alu_ashr_7_n817, alu_ashr_7_n816, alu_ashr_7_n815, alu_ashr_7_n814,
         alu_ashr_7_n813, alu_ashr_7_n812, alu_ashr_7_n811, alu_ashr_7_n810,
         alu_ashr_7_n809, alu_ashr_7_n808, alu_ashr_7_n807, alu_ashr_7_n806,
         alu_ashr_7_n805, alu_ashr_7_n804, alu_ashr_7_n803, alu_ashr_7_n802,
         alu_ashr_7_n801, alu_ashr_7_n800, alu_ashr_7_n799, alu_ashr_7_n798,
         alu_ashr_7_n797, alu_ashr_7_n796, alu_ashr_7_n795, alu_ashr_7_n794,
         alu_ashr_7_n793, alu_ashr_7_n792, alu_ashr_7_n791, alu_ashr_7_n790,
         alu_ashr_7_n789, alu_ashr_7_n788, alu_ashr_7_n787, alu_ashr_7_n786,
         alu_ashr_7_n785, alu_ashr_7_n784, alu_ashr_7_n783, alu_ashr_7_n782,
         alu_ashr_7_n781, alu_ashr_7_n780, alu_ashr_7_n779, alu_ashr_7_n778,
         alu_ashr_7_n777, alu_ashr_7_n776, alu_ashr_7_n775, alu_ashr_7_n774,
         alu_ashr_7_n773, alu_ashr_7_n772, alu_ashr_7_n771, alu_ashr_7_n770,
         alu_ashr_7_n769, alu_ashr_7_n768, alu_ashr_7_n767, alu_ashr_7_n766,
         alu_ashr_7_n765, alu_ashr_7_n764, alu_ashr_7_n763, alu_ashr_7_n762,
         alu_ashr_7_n761, alu_ashr_7_n760, alu_ashr_7_n759, alu_ashr_7_n758,
         alu_ashr_7_n757, alu_ashr_7_n756, alu_ashr_7_n755, alu_ashr_7_n754,
         alu_ashr_7_n753, alu_ashr_7_n752, alu_ashr_7_n751, alu_ashr_7_n750,
         alu_ashr_7_n749, alu_ashr_7_n748, alu_ashr_7_n747, alu_ashr_7_n746,
         alu_ashr_7_n745, alu_ashr_7_n744, alu_ashr_7_n743, alu_ashr_7_n742,
         alu_ashr_7_n741, alu_ashr_7_n740, alu_ashr_7_n739, alu_ashr_7_n738,
         alu_ashr_7_n737, alu_ashr_7_n736, alu_ashr_7_n735, alu_ashr_7_n734,
         alu_ashr_7_n733, alu_ashr_7_n732, alu_ashr_7_n731, alu_ashr_7_n730,
         alu_ashr_7_n729, alu_ashr_7_n728, alu_ashr_7_n727, alu_ashr_7_n726,
         alu_ashr_7_n725, alu_ashr_7_n724, alu_ashr_7_n723, alu_ashr_7_n722,
         alu_ashr_7_n721, alu_ashr_7_n720, alu_ashr_7_n719, alu_ashr_7_n718,
         alu_ashr_7_n717, alu_ashr_7_n716, alu_ashr_7_n715, alu_ashr_7_n714,
         alu_ashr_7_n713, alu_ashr_7_n712, alu_ashr_7_n711, alu_ashr_7_n710,
         alu_ashr_7_n709, alu_ashr_7_n708, alu_ashr_7_n707, alu_ashr_7_n706,
         alu_ashr_7_n705, alu_ashr_7_n704, alu_ashr_7_n703, alu_ashr_7_n702,
         alu_ashr_7_n701, alu_ashr_7_n700, alu_ashr_7_n699, alu_ashr_7_n698,
         alu_ashr_7_n697, alu_ashr_7_n696, alu_ashr_7_n695, alu_ashr_7_n694,
         alu_ashr_7_n693, alu_ashr_7_n692, alu_ashr_7_n691, alu_ashr_7_n690,
         alu_ashr_7_n689, alu_ashr_7_n688, alu_ashr_7_n687, alu_ashr_7_n686,
         alu_ashr_7_n685, alu_ashr_7_n684, alu_ashr_7_n683, alu_ashr_7_n682,
         alu_ashr_7_n681, alu_ashr_7_n680, alu_ashr_7_n679, alu_ashr_7_n678,
         alu_ashr_7_n677, alu_ashr_7_n676, alu_ashr_7_n675, alu_ashr_7_n674,
         alu_ashr_7_n673, alu_ashr_7_n672, alu_ashr_7_n671, alu_ashr_7_n670,
         alu_ashr_7_n669, alu_ashr_7_n668, alu_ashr_7_n667, alu_ashr_7_n666,
         alu_ashr_7_n665, alu_ashr_7_n664, alu_ashr_7_n663, alu_ashr_7_n662,
         alu_ashr_7_n661, alu_ashr_7_n660, alu_ashr_7_n659, alu_ashr_7_n658,
         alu_ashr_7_n657, alu_ashr_7_n656, alu_ashr_7_n655, alu_ashr_7_n654,
         alu_ashr_7_n653, alu_ashr_7_n652, alu_ashr_7_n651, alu_ashr_7_n650,
         alu_ashr_7_n649, alu_ashr_7_n648, alu_ashr_7_n647, alu_ashr_7_n646,
         alu_ashr_7_n645, alu_ashr_7_n644, alu_ashr_7_n643, alu_ashr_7_n642,
         alu_ashr_7_n641, alu_ashr_7_n640, alu_ashr_7_n639, alu_ashr_7_n638,
         alu_ashr_7_n637, alu_ashr_7_n636, alu_ashr_7_n635, alu_ashr_7_n634,
         alu_ashr_7_n633, alu_ashr_7_n632, alu_ashr_7_n631, alu_ashr_7_n630,
         alu_ashr_7_n629, alu_ashr_7_n628, alu_ashr_7_n627, alu_ashr_7_n626,
         alu_ashr_7_n625, alu_ashr_7_n624, alu_ashr_7_n623, alu_ashr_7_n622,
         alu_ashr_7_n621, alu_ashr_7_n620, alu_ashr_7_n619, alu_ashr_7_n618,
         alu_ashr_7_n617, alu_ashr_7_n616, alu_ashr_7_n615, alu_ashr_7_n614,
         alu_ashr_7_n613, alu_ashr_7_n612, alu_ashr_7_n611, alu_ashr_7_n610,
         alu_ashr_7_n609, alu_ashr_7_n608, alu_ashr_7_n607, alu_ashr_7_n606,
         alu_ashr_7_n605, alu_ashr_7_n604, alu_ashr_7_n603, alu_ashr_7_n602,
         alu_ashr_7_n601, alu_ashr_7_n600, alu_ashr_7_n599, alu_ashr_7_n598,
         alu_ashr_7_n597, alu_ashr_7_n596, alu_ashr_7_n595, alu_ashr_7_n594,
         alu_ashr_7_n593, alu_ashr_7_n592, alu_ashr_7_n591, alu_ashr_7_n590,
         alu_ashr_7_n589, alu_ashr_7_n588, alu_ashr_7_n587, alu_ashr_7_n586,
         alu_ashr_7_n585, alu_ashr_7_n584, alu_ashr_7_n583, alu_ashr_7_n582,
         alu_ashr_7_n581, alu_ashr_7_n580, alu_ashr_7_n579, alu_ashr_7_n578,
         alu_ashr_7_n577, alu_ashr_7_n576, alu_ashr_7_n575, alu_ashr_7_n574,
         alu_ashr_7_n573, alu_ashr_7_n572, alu_ashr_7_n571, alu_ashr_7_n570,
         alu_ashr_7_n569, alu_ashr_7_n568, alu_ashr_7_n567, alu_ashr_7_n566,
         alu_ashr_7_n565, alu_ashr_7_n564, alu_ashr_7_n563, alu_ashr_7_n562,
         alu_ashr_7_n561, alu_ashr_7_n560, alu_ashr_7_n559, alu_ashr_7_n558,
         alu_ashr_7_n557, alu_ashr_7_n556, alu_ashr_7_n555, alu_ashr_7_n554,
         alu_ashr_7_n553, alu_ashr_7_n552, alu_ashr_7_n551, alu_ashr_7_n550,
         alu_ashr_7_n549, alu_ashr_7_n548, alu_ashr_7_n547, alu_ashr_7_n546,
         alu_ashr_7_n545, alu_ashr_7_n544, alu_ashr_7_n543, alu_ashr_7_n542,
         alu_ashr_7_n541, alu_ashr_7_n540, alu_ashr_7_n539, alu_ashr_7_n538,
         alu_ashr_7_n537, alu_ashr_7_n536, alu_ashr_7_n535, alu_ashr_7_n534,
         alu_ashr_7_n533, alu_ashr_7_n532, alu_ashr_7_n531, alu_ashr_7_n530,
         alu_ashr_7_n529, alu_ashr_7_n528, alu_ashr_7_n527, alu_ashr_7_n526,
         alu_ashr_7_n525, alu_ashr_7_n524, alu_ashr_7_n523, alu_ashr_7_n522,
         alu_ashr_7_n521, alu_ashr_7_n520, alu_ashr_7_n519, alu_ashr_7_n518,
         alu_ashr_7_n517, alu_ashr_7_n516, alu_ashr_7_n515, alu_ashr_7_n514,
         alu_ashr_7_n513, alu_ashr_7_n512, alu_ashr_7_n511, alu_ashr_7_n510,
         alu_ashr_7_n509, alu_ashr_7_n508, alu_ashr_7_n507, alu_ashr_7_n506,
         alu_ashr_7_n505, alu_ashr_7_n504, alu_ashr_7_n503, alu_ashr_7_n502,
         alu_ashr_7_n501, alu_ashr_7_n500, alu_ashr_7_n499, alu_ashr_7_n498,
         alu_ashr_7_n497, alu_ashr_7_n496, alu_ashr_7_n495, alu_ashr_7_n493,
         alu_ashr_7_n492, div_SYNOPSYS_UNCONNECTED_64,
         div_SYNOPSYS_UNCONNECTED_63, div_SYNOPSYS_UNCONNECTED_62,
         div_SYNOPSYS_UNCONNECTED_61, div_SYNOPSYS_UNCONNECTED_60,
         div_SYNOPSYS_UNCONNECTED_59, div_SYNOPSYS_UNCONNECTED_58,
         div_SYNOPSYS_UNCONNECTED_57, div_SYNOPSYS_UNCONNECTED_56,
         div_SYNOPSYS_UNCONNECTED_55, div_SYNOPSYS_UNCONNECTED_54,
         div_SYNOPSYS_UNCONNECTED_53, div_SYNOPSYS_UNCONNECTED_52,
         div_SYNOPSYS_UNCONNECTED_51, div_SYNOPSYS_UNCONNECTED_50,
         div_SYNOPSYS_UNCONNECTED_49, div_SYNOPSYS_UNCONNECTED_48,
         div_SYNOPSYS_UNCONNECTED_47, div_SYNOPSYS_UNCONNECTED_46,
         div_SYNOPSYS_UNCONNECTED_45, div_SYNOPSYS_UNCONNECTED_44,
         div_SYNOPSYS_UNCONNECTED_43, div_SYNOPSYS_UNCONNECTED_42,
         div_SYNOPSYS_UNCONNECTED_41, div_SYNOPSYS_UNCONNECTED_40,
         div_SYNOPSYS_UNCONNECTED_39, div_SYNOPSYS_UNCONNECTED_38,
         div_SYNOPSYS_UNCONNECTED_37, div_SYNOPSYS_UNCONNECTED_36,
         div_SYNOPSYS_UNCONNECTED_35, div_SYNOPSYS_UNCONNECTED_34,
         div_SYNOPSYS_UNCONNECTED_33, div_SYNOPSYS_UNCONNECTED_32,
         div_SYNOPSYS_UNCONNECTED_31, div_SYNOPSYS_UNCONNECTED_30,
         div_SYNOPSYS_UNCONNECTED_29, div_SYNOPSYS_UNCONNECTED_28,
         div_SYNOPSYS_UNCONNECTED_27, div_SYNOPSYS_UNCONNECTED_26,
         div_SYNOPSYS_UNCONNECTED_25, div_SYNOPSYS_UNCONNECTED_24,
         div_SYNOPSYS_UNCONNECTED_23, div_SYNOPSYS_UNCONNECTED_22,
         div_SYNOPSYS_UNCONNECTED_21, div_SYNOPSYS_UNCONNECTED_20,
         div_SYNOPSYS_UNCONNECTED_19, div_SYNOPSYS_UNCONNECTED_18,
         div_SYNOPSYS_UNCONNECTED_17, div_SYNOPSYS_UNCONNECTED_16,
         div_SYNOPSYS_UNCONNECTED_15, div_SYNOPSYS_UNCONNECTED_14,
         div_SYNOPSYS_UNCONNECTED_13, div_SYNOPSYS_UNCONNECTED_12,
         div_SYNOPSYS_UNCONNECTED_11, div_SYNOPSYS_UNCONNECTED_10,
         div_SYNOPSYS_UNCONNECTED_9, div_SYNOPSYS_UNCONNECTED_8,
         div_SYNOPSYS_UNCONNECTED_7, div_SYNOPSYS_UNCONNECTED_6,
         div_SYNOPSYS_UNCONNECTED_5, div_SYNOPSYS_UNCONNECTED_4,
         div_SYNOPSYS_UNCONNECTED_3, div_SYNOPSYS_UNCONNECTED_2,
         div_SYNOPSYS_UNCONNECTED_1, div_n1003, div_n1002, div_n1001,
         div_n1000, div_n999, div_n998, div_n997, div_n996, div_n995, div_n994,
         div_n993, div_n992, div_n991, div_n990, div_n989, div_n988, div_n987,
         div_n986, div_n985, div_n984, div_n983, div_n982, div_n981, div_n980,
         div_n979, div_n978, div_n977, div_n976, div_n975, div_n974, div_n973,
         div_n972, div_n971, div_n970, div_n969, div_n968, div_n967, div_n966,
         div_n965, div_n964, div_n963, div_n962, div_n961, div_n960, div_n959,
         div_n958, div_n957, div_n956, div_n955, div_n954, div_n953, div_n952,
         div_n951, div_n950, div_n949, div_n948, div_n947, div_n946, div_n945,
         div_n944, div_n943, div_n942, div_n941, div_n940, div_n939, div_n938,
         div_n937, div_n936, div_n935, div_n934, div_n933, div_n932, div_n931,
         div_n930, div_n929, div_n928, div_n927, div_n926, div_n925, div_n924,
         div_n923, div_n922, div_n921, div_n920, div_n919, div_n918, div_n917,
         div_n916, div_n915, div_n914, div_n913, div_n912, div_n911, div_n910,
         div_n909, div_n908, div_n907, div_n906, div_n905, div_n904, div_n903,
         div_n902, div_n901, div_n900, div_n899, div_n898, div_n897, div_n896,
         div_n895, div_n894, div_n893, div_n892, div_n891, div_n890, div_n889,
         div_n888, div_n887, div_n886, div_n885, div_n884, div_n883, div_n882,
         div_n881, div_n880, div_n879, div_n878, div_n877, div_n876, div_n875,
         div_n874, div_n873, div_n872, div_n871, div_n870, div_n869, div_n868,
         div_n867, div_n866, div_n865, div_n864, div_n863, div_n862, div_n861,
         div_n860, div_n859, div_n858, div_n857, div_n856, div_n855, div_n854,
         div_n853, div_n852, div_n851, div_n850, div_n849, div_n848, div_n847,
         div_n846, div_n845, div_n844, div_n843, div_n842, div_n841, div_n840,
         div_n839, div_n838, div_n837, div_n836, div_n835, div_n834, div_n833,
         div_n832, div_n831, div_n830, div_n829, div_n828, div_n827, div_n826,
         div_n825, div_n824, div_n823, div_n822, div_n821, div_n820, div_n819,
         div_n818, div_n817, div_n816, div_n815, div_n814, div_n813, div_n812,
         div_n811, div_n810, div_n809, div_n808, div_n807, div_n806, div_n805,
         div_n804, div_n803, div_n802, div_n801, div_n800, div_n799, div_n798,
         div_n797, div_n795, div_n792, div_n791, div_n790, div_n789, div_n788,
         div_n787, div_n786, div_n785, div_n784, div_n783, div_n782, div_n781,
         div_n780, div_n779, div_n778, div_n777, div_n776, div_n775, div_n774,
         div_n773, div_n772, div_n771, div_n770, div_n769, div_n768, div_n767,
         div_n766, div_n765, div_n764, div_n763, div_n762, div_n761, div_n760,
         div_n759, div_n758, div_n757, div_n756, div_n755, div_n754, div_n753,
         div_n752, div_n751, div_n750, div_n749, div_n748, div_n747, div_n746,
         div_n745, div_n744, div_n743, div_n742, div_n741, div_n740, div_n739,
         div_n738, div_n737, div_n736, div_n735, div_n734, div_n733, div_n732,
         div_n731, div_n730, div_n729, div_n728, div_n727, div_n726, div_n725,
         div_n724, div_n723, div_n722, div_n721, div_n720, div_n719, div_n718,
         div_n717, div_n716, div_n715, div_n714, div_n713, div_n712, div_n711,
         div_n710, div_n709, div_n708, div_n707, div_n706, div_n705, div_n704,
         div_n703, div_n702, div_n701, div_n700, div_n699, div_n698, div_n697,
         div_n696, div_n695, div_n694, div_n693, div_n692, div_n691, div_n690,
         div_n689, div_n688, div_n687, div_n686, div_n685, div_n684, div_n683,
         div_n682, div_n681, div_n680, div_n679, div_n678, div_n677, div_n676,
         div_n675, div_n674, div_n673, div_n672, div_n671, div_n670, div_n669,
         div_n668, div_n667, div_n666, div_n665, div_n664, div_n663, div_n662,
         div_n661, div_n660, div_n659, div_n658, div_n657, div_n656, div_n655,
         div_n654, div_n653, div_n652, div_n651, div_n650, div_n649, div_n648,
         div_n647, div_n646, div_n645, div_n644, div_n643, div_n642, div_n641,
         div_n640, div_n639, div_n638, div_n637, div_n636, div_n635, div_n634,
         div_n633, div_n632, div_n631, div_n630, div_n629, div_n628, div_n627,
         div_n626, div_n625, div_n624, div_n623, div_n622, div_n621, div_n620,
         div_n619, div_n618, div_n617, div_n616, div_n615, div_n614, div_n613,
         div_n612, div_n611, div_n610, div_n609, div_n608, div_n607, div_n606,
         div_n605, div_n604, div_n603, div_n602, div_n601, div_n600, div_n599,
         div_n598, div_n597, div_n596, div_n595, div_n594, div_n593, div_n592,
         div_n591, div_n590, div_n589, div_n588, div_n587, div_n586, div_n585,
         div_n584, div_n583, div_n582, div_n581, div_n580, div_n579, div_n578,
         div_n577, div_n576, div_n575, div_n574, div_n573, div_n572, div_n571,
         div_n570, div_n569, div_n568, div_n567, div_n566, div_n565, div_n564,
         div_n563, div_n562, div_n561, div_n560, div_n559, div_n558, div_n557,
         div_n556, div_n555, div_n554, div_n553, div_n552, div_n551, div_n550,
         div_n549, div_n548, div_n547, div_n546, div_n545, div_n544, div_n543,
         div_n542, div_n541, div_n540, div_n539, div_n538, div_n537, div_n536,
         div_n535, div_n534, div_n533, div_n532, div_n531, div_n530, div_n529,
         div_n528, div_n527, div_n526, div_n525, div_n524, div_n523, div_n522,
         div_n521, div_n520, div_n519, div_n518, div_n517, div_n516, div_n515,
         div_n514, div_n513, div_n512, div_n511, div_n510, div_n509, div_n508,
         div_n507, div_n506, div_n505, div_n504, div_n503, div_n502, div_n501,
         div_n500, div_n499, div_n498, div_n497, div_n496, div_n495, div_n494,
         div_n493, div_n492, div_n491, div_n490, div_n489, div_n488, div_n487,
         div_n486, div_n485, div_n484, div_n483, div_n482, div_n481, div_n480,
         div_n479, div_n478, div_n477, div_n476, div_n475, div_n474, div_n473,
         div_n472, div_n471, div_n470, div_n469, div_n468, div_n467, div_n466,
         div_n465, div_n464, div_n463, div_n462, div_n461, div_n460, div_n459,
         div_n458, div_n457, div_n456, div_n455, div_n454, div_n453, div_n452,
         div_n451, div_n450, div_n449, div_n448, div_n447, div_n446, div_n445,
         div_n444, div_n443, div_n442, div_n441, div_n440, div_n439, div_n438,
         div_n437, div_n436, div_n435, div_n434, div_n433, div_n432, div_n431,
         div_n430, div_n429, div_n428, div_n427, div_n426, div_n425, div_n424,
         div_n423, div_n422, div_n421, div_n420, div_n419, div_n418, div_n417,
         div_n416, div_n415, div_n414, div_n413, div_n412, div_n411, div_n410,
         div_n409, div_n408, div_n407, div_n406, div_n405, div_n404, div_n403,
         div_n402, div_n401, div_n400, div_n399, div_n398, div_n397, div_n396,
         div_n395, div_n394, div_n393, div_n392, div_n391, div_n390, div_n389,
         div_n388, div_n387, div_n386, div_n385, div_n384, div_n383, div_n382,
         div_n381, div_n380, div_n379, div_n378, div_n377, div_n376, div_n375,
         div_n374, div_n373, div_n372, div_n371, div_n370, div_n369, div_n368,
         div_n367, div_n366, div_n365, div_n364, div_n363, div_n362, div_n361,
         div_n360, div_n359, div_n358, div_n357, div_n356, div_n355, div_n354,
         div_n353, div_n352, div_n351, div_n350, div_n349, div_n348, div_n347,
         div_n346, div_n345, div_n344, div_n343, div_n342, div_n341, div_n340,
         div_n339, div_n338, div_n337, div_n336, div_n335, div_n334, div_n333,
         div_n332, div_n331, div_n330, div_n329, div_n328, div_n327, div_n326,
         div_n325, div_n324, div_n323, div_n322, div_n321, div_n320, div_n319,
         div_n318, div_n317, div_n316, div_n315, div_n314, div_n313, div_n312,
         div_n311, div_n310, div_n309, div_n308, div_n307, div_n306, div_n305,
         div_n304, div_n303, div_n302, div_n301, div_n300, div_n299, div_n298,
         div_n297, div_n295, div_n294, div_n289, div_n288, div_n287, div_n285,
         div_n280, div_n279, div_n276, div_n271, div_n265, div_n262, div_n253,
         div_n245, div_n244, div_n242, div_n235, div_n230, div_n227, div_n226,
         div_n225, div_n224, div_n223, div_n222, div_n221, div_n218, div_n216,
         div_n215, div_n214, div_n213, div_n212, div_n211, div_n210, div_n209,
         div_n208, div_n207, div_n206, div_n204, div_n203, div_n201, div_n200,
         div_n199, div_n198, div_n197, div_n195, div_n194, div_n193, div_n192,
         div_n191, div_n190, div_n189, div_n188, div_n187, div_n186, div_n184,
         div_n183, div_n182, div_n181, div_n180, div_n178, div_n177, div_n176,
         div_n175, div_n174, div_n173, div_n172, div_n165, div_n164, div_n163,
         div_n162, div_n161, div_n160, div_n159, div_n158, div_n157, div_n156,
         div_n155, div_n154, div_n153, div_n152, div_n151, div_n150, div_n149,
         div_n148, div_n147, div_n146, div_n145, div_n141, div_n140, div_n139,
         div_n138, div_n137, div_n136, div_n135, div_n133, div_n132, div_n131,
         div_n130, div_n129, div_n128, div_n127, div_n126, div_n125, div_n124,
         div_n123, div_n121, div_n120, div_n118, div_n117, div_n116, div_n115,
         div_n114, div_n113, div_n112, div_n111, div_n110, div_n109, div_n108,
         div_n106, div_n105, div_n104, div_n103, div_n102, div_n101, div_n100,
         div_n98, div_n97, div_n96, div_n95, div_n93, div_n92, div_n91,
         div_n90, div_n88, div_n87, div_n86, div_n85, div_n83, div_n82,
         div_n81, div_n80, div_n78, div_n77, div_n76, div_n75, div_n73,
         div_n72, div_n71, div_n70, div_n69, div_n68, div_n66, div_n65,
         div_n64, div_n63, div_n62, div_n61, div_n60, div_n59, div_n58,
         div_n56, div_n55, div_n54, div_n53, div_n52, div_n51, div_n50,
         div_n49, div_n48, div_n47, div_n45, div_n44, div_n43, div_n41,
         div_n40, div_n39, div_n38, div_n37, div_n36, div_n35, div_n34,
         div_n33, div_n32, div_n31, div_n30, div_n29, div_n28, div_n27,
         div_n26, div_n25, div_n24, div_n22, div_n21, div_n20, div_n19,
         div_n18, div_n17, div_n16, div_n15, div_n14, div_n13, div_n12,
         div_n11, div_n10, div_n9, div_n8, div_n7, div_n6, div_n5, div_n4,
         div_n3, div_n2, div_n794, div_n793, div_n296, div_n293, div_n292,
         div_n291, div_n290, div_n286, div_n284, div_n283, div_n282, div_n281,
         div_n278, div_n277, div_n275, div_n274, div_n273, div_n272, div_n270,
         div_n269, div_n268, div_n267, div_n266, div_n264, div_n263, div_n261,
         div_n260, div_n259, div_n258, div_n257, div_n256, div_n255, div_n254,
         div_n252, div_n251, div_n250, div_n249, div_n248, div_n247, div_n246,
         div_n243, div_n241, div_n240, div_n239, div_n238, div_n237, div_n236,
         div_n234, div_n233, div_n232, div_n231, div_n229, div_n228, div_n220,
         div_n219, div_n217, div_n205, div_n202, div_n196, div_n185, div_n179,
         div_n171, div_n170, div_n169, div_n168, div_n167, div_n166,
         div_net34705, div_net34700, div_net34695, div_net34690, div_net34684,
         div_N523, div_N522, div_N521, div_N520, div_N519, div_N518, div_N517,
         div_N516, div_N515, div_N514, div_N513, div_N512, div_N511, div_N510,
         div_N509, div_N508, div_N507, div_N506, div_N505, div_N504, div_N503,
         div_N502, div_N501, div_N500, div_N499, div_N498, div_N497, div_N496,
         div_N495, div_N494, div_N493, div_N492, div_N491, div_N490, div_N489,
         div_N488, div_N487, div_N486, div_N485, div_N484, div_N483, div_N482,
         div_N481, div_N480, div_N479, div_N478, div_N477, div_N476, div_N475,
         div_N474, div_N473, div_N472, div_N471, div_N470, div_N469, div_N468,
         div_N467, div_N466, div_N465, div_N464, div_N463, div_N462, div_N461,
         div_N460, div_N459, div_N458, div_N457, div_N456, div_N455, div_N454,
         div_N453, div_N452, div_N451, div_N450, div_N449, div_N448, div_N447,
         div_N446, div_N445, div_N444, div_N443, div_N442, div_N441, div_N440,
         div_N439, div_N438, div_N437, div_N436, div_N435, div_N434, div_N433,
         div_N432, div_N431, div_N430, div_N429, div_N428, div_N427, div_N426,
         div_N425, div_N424, div_N423, div_N422, div_N421, div_N420, div_N419,
         div_N418, div_N417, div_N416, div_N415, div_N414, div_N413, div_N412,
         div_N411, div_N410, div_N409, div_N408, div_N407, div_N406, div_N405,
         div_N404, div_N403, div_N402, div_N401, div_N400, div_N399, div_N398,
         div_N397, div_N396, div_N395, div_N394, div_N387, div_N386, div_N385,
         div_N384, div_N383, div_N382, div_N381, div_N380, div_N379, div_N378,
         div_N377, div_N376, div_N375, div_N374, div_N373, div_N372, div_N371,
         div_N370, div_N369, div_N368, div_N367, div_N366, div_N365, div_N364,
         div_N363, div_N362, div_N361, div_N360, div_N359, div_N358, div_N357,
         div_N356, div_N355, div_N354, div_N353, div_N352, div_N351, div_N350,
         div_N349, div_N348, div_N347, div_N346, div_N345, div_N344, div_N343,
         div_N342, div_N341, div_N340, div_N339, div_N338, div_N337, div_N336,
         div_N335, div_N334, div_N333, div_N332, div_N331, div_N330, div_N329,
         div_N328, div_N327, div_N326, div_N325, div_N324, div_N323, div_N322,
         div_N299, div_N298, div_N297, div_N296, div_N295, div_N294, div_N293,
         div_N285, div_N284, div_N283, div_N282, div_n_T_434_0_,
         div_n_T_434_1_, div_n_T_434_2_, div_n_T_434_3_, div_n_T_434_4_,
         div_n_T_434_5_, div_n_T_430_5_, div_n_T_273_5_, div_n_T_97_6_,
         div_n_T_85_4_, div_n_T_85_5_, div_isHi, div_n_T_71_39_, div_n_T_69_4_,
         div_n_T_69_6_, div_n_T_69_7_, div_n_T_69_8_, div_n_T_69_9_,
         div_neg_out, div_n_T_59_8_, div_n_T_51_0_, div_n_T_51_1_,
         div_n_T_51_3_, div_n_T_51_4_, div_n_T_51_5_, div_n_T_51_6_,
         div_n_T_51_7_, div_n_T_51_8_, div_n_T_51_9_, div_n_T_51_10_,
         div_n_T_51_11_, div_n_T_51_12_, div_n_T_51_13_, div_n_T_51_14_,
         div_n_T_51_15_, div_n_T_51_16_, div_n_T_51_17_, div_n_T_51_18_,
         div_n_T_51_19_, div_n_T_51_20_, div_n_T_51_21_, div_n_T_51_22_,
         div_n_T_51_23_, div_n_T_51_24_, div_n_T_51_25_, div_n_T_51_26_,
         div_n_T_51_27_, div_n_T_51_28_, div_n_T_51_29_, div_n_T_51_30_,
         div_n_T_51_31_, div_n_T_51_32_, div_n_T_51_33_, div_n_T_51_34_,
         div_n_T_51_35_, div_n_T_51_36_, div_n_T_51_37_, div_n_T_51_38_,
         div_n_T_51_39_, div_n_T_51_40_, div_n_T_51_41_, div_n_T_51_42_,
         div_n_T_51_43_, div_n_T_51_44_, div_n_T_51_45_, div_n_T_51_46_,
         div_n_T_51_47_, div_n_T_51_48_, div_n_T_51_49_, div_n_T_51_50_,
         div_n_T_51_51_, div_n_T_51_52_, div_n_T_51_53_, div_n_T_51_54_,
         div_n_T_51_55_, div_n_T_51_56_, div_n_T_51_57_, div_n_T_51_58_,
         div_n_T_51_59_, div_n_T_51_60_, div_n_T_51_61_, div_n_T_51_62_,
         div_n_T_51_63_, div_n_T_51_64_, div_n_T_51_65_, div_n_T_51_66_,
         div_n_T_51_67_, div_n_T_51_68_, div_n_T_51_69_, div_n_T_51_70_,
         div_n_T_51_71_, div_n_T_51_72_, div_n_T_51_73_, div_n_T_51_74_,
         div_n_T_51_75_, div_n_T_51_76_, div_n_T_51_77_, div_n_T_51_78_,
         div_n_T_51_79_, div_n_T_51_80_, div_n_T_51_81_, div_n_T_51_82_,
         div_n_T_51_83_, div_n_T_51_84_, div_n_T_51_85_, div_n_T_51_86_,
         div_n_T_51_87_, div_n_T_51_88_, div_n_T_51_89_, div_n_T_51_90_,
         div_n_T_51_91_, div_n_T_51_92_, div_n_T_51_93_, div_n_T_51_94_,
         div_n_T_51_95_, div_n_T_51_96_, div_n_T_51_97_, div_n_T_51_98_,
         div_n_T_51_99_, div_n_T_51_100_, div_n_T_51_101_, div_n_T_51_102_,
         div_n_T_51_103_, div_n_T_51_104_, div_n_T_51_105_, div_n_T_51_106_,
         div_n_T_51_107_, div_n_T_51_108_, div_n_T_51_109_, div_n_T_51_110_,
         div_n_T_51_111_, div_n_T_51_112_, div_n_T_51_113_, div_n_T_51_114_,
         div_n_T_51_115_, div_n_T_51_116_, div_n_T_51_117_, div_n_T_51_118_,
         div_n_T_51_119_, div_n_T_51_120_, div_n_T_51_121_, div_n_T_51_122_,
         div_n_T_51_123_, div_n_T_51_124_, div_n_T_51_125_, div_n_T_51_126_,
         div_n_T_51_127_, div_n_T_51_128_, div_result_0_, div_result_1_,
         div_result_2_, div_result_3_, div_result_4_, div_result_5_,
         div_result_6_, div_result_7_, div_result_8_, div_result_9_,
         div_result_10_, div_result_11_, div_result_12_, div_result_13_,
         div_result_14_, div_result_15_, div_result_16_, div_result_17_,
         div_result_18_, div_result_19_, div_result_20_, div_result_21_,
         div_result_22_, div_result_23_, div_result_24_, div_result_25_,
         div_result_26_, div_result_27_, div_result_28_, div_result_29_,
         div_result_30_, div_result_31_, div_result_32_, div_result_33_,
         div_result_34_, div_result_35_, div_result_36_, div_result_37_,
         div_result_38_, div_result_39_, div_result_40_, div_result_41_,
         div_result_42_, div_result_43_, div_result_44_, div_result_45_,
         div_result_46_, div_result_47_, div_result_48_, div_result_49_,
         div_result_50_, div_result_51_, div_result_52_, div_result_53_,
         div_result_54_, div_result_55_, div_result_56_, div_result_57_,
         div_result_58_, div_result_59_, div_result_60_, div_result_61_,
         div_result_62_, div_result_63_, div_resHi, div_subtractor_0_,
         div_subtractor_1_, div_subtractor_2_, div_subtractor_3_,
         div_subtractor_4_, div_subtractor_5_, div_subtractor_6_,
         div_subtractor_7_, div_subtractor_8_, div_subtractor_9_,
         div_subtractor_10_, div_subtractor_11_, div_subtractor_12_,
         div_subtractor_13_, div_subtractor_14_, div_subtractor_15_,
         div_subtractor_16_, div_subtractor_17_, div_subtractor_18_,
         div_subtractor_19_, div_subtractor_20_, div_subtractor_21_,
         div_subtractor_22_, div_subtractor_23_, div_subtractor_24_,
         div_subtractor_25_, div_subtractor_26_, div_subtractor_27_,
         div_subtractor_28_, div_subtractor_29_, div_subtractor_30_,
         div_subtractor_31_, div_subtractor_32_, div_subtractor_33_,
         div_subtractor_34_, div_subtractor_35_, div_subtractor_36_,
         div_subtractor_37_, div_subtractor_38_, div_subtractor_39_,
         div_subtractor_40_, div_subtractor_41_, div_subtractor_42_,
         div_subtractor_43_, div_subtractor_44_, div_subtractor_45_,
         div_subtractor_46_, div_subtractor_47_, div_subtractor_48_,
         div_subtractor_49_, div_subtractor_50_, div_subtractor_51_,
         div_subtractor_52_, div_subtractor_53_, div_subtractor_54_,
         div_subtractor_55_, div_subtractor_56_, div_subtractor_57_,
         div_subtractor_58_, div_subtractor_59_, div_subtractor_60_,
         div_subtractor_61_, div_subtractor_62_, div_subtractor_63_,
         div_subtractor_64_, div_divisor_0_, div_divisor_1_, div_divisor_2_,
         div_divisor_3_, div_divisor_4_, div_divisor_5_, div_divisor_6_,
         div_divisor_7_, div_divisor_8_, div_divisor_9_, div_divisor_10_,
         div_divisor_11_, div_divisor_12_, div_divisor_13_, div_divisor_14_,
         div_divisor_15_, div_divisor_16_, div_divisor_17_, div_divisor_18_,
         div_divisor_19_, div_divisor_20_, div_divisor_21_, div_divisor_22_,
         div_divisor_23_, div_divisor_24_, div_divisor_25_, div_divisor_26_,
         div_divisor_27_, div_divisor_28_, div_divisor_29_, div_divisor_30_,
         div_divisor_31_, div_divisor_32_, div_divisor_33_, div_divisor_34_,
         div_divisor_35_, div_divisor_36_, div_divisor_37_, div_divisor_38_,
         div_divisor_39_, div_divisor_40_, div_divisor_41_, div_divisor_42_,
         div_divisor_43_, div_divisor_44_, div_divisor_45_, div_divisor_46_,
         div_divisor_47_, div_divisor_48_, div_divisor_49_, div_divisor_50_,
         div_divisor_51_, div_divisor_52_, div_divisor_53_, div_divisor_54_,
         div_divisor_55_, div_divisor_56_, div_divisor_57_, div_divisor_58_,
         div_divisor_59_, div_divisor_60_, div_divisor_61_, div_divisor_62_,
         div_divisor_63_, div_divisor_64_, div_DP_OP_279J39_124_314_n2787,
         div_DP_OP_279J39_124_314_n2786, div_DP_OP_279J39_124_314_n2785,
         div_DP_OP_279J39_124_314_n2784, div_DP_OP_279J39_124_314_n2783,
         div_DP_OP_279J39_124_314_n2782, div_DP_OP_279J39_124_314_n2781,
         div_DP_OP_279J39_124_314_n2780, div_DP_OP_279J39_124_314_n2779,
         div_DP_OP_279J39_124_314_n2778, div_DP_OP_279J39_124_314_n2777,
         div_DP_OP_279J39_124_314_n2776, div_DP_OP_279J39_124_314_n2775,
         div_DP_OP_279J39_124_314_n2774, div_DP_OP_279J39_124_314_n2773,
         div_DP_OP_279J39_124_314_n2772, div_DP_OP_279J39_124_314_n2771,
         div_DP_OP_279J39_124_314_n2770, div_DP_OP_279J39_124_314_n2769,
         div_DP_OP_279J39_124_314_n2768, div_DP_OP_279J39_124_314_n2767,
         div_DP_OP_279J39_124_314_n2766, div_DP_OP_279J39_124_314_n2765,
         div_DP_OP_279J39_124_314_n2764, div_DP_OP_279J39_124_314_n2763,
         div_DP_OP_279J39_124_314_n2762, div_DP_OP_279J39_124_314_n2761,
         div_DP_OP_279J39_124_314_n2760, div_DP_OP_279J39_124_314_n2759,
         div_DP_OP_279J39_124_314_n2758, div_DP_OP_279J39_124_314_n2757,
         div_DP_OP_279J39_124_314_n2756, div_DP_OP_279J39_124_314_n2755,
         div_DP_OP_279J39_124_314_n2754, div_DP_OP_279J39_124_314_n2753,
         div_DP_OP_279J39_124_314_n2752, div_DP_OP_279J39_124_314_n2751,
         div_DP_OP_279J39_124_314_n2750, div_DP_OP_279J39_124_314_n2749,
         div_DP_OP_279J39_124_314_n2748, div_DP_OP_279J39_124_314_n2747,
         div_DP_OP_279J39_124_314_n2746, div_DP_OP_279J39_124_314_n2745,
         div_DP_OP_279J39_124_314_n2744, div_DP_OP_279J39_124_314_n2743,
         div_DP_OP_279J39_124_314_n2742, div_DP_OP_279J39_124_314_n2741,
         div_DP_OP_279J39_124_314_n2740, div_DP_OP_279J39_124_314_n2739,
         div_DP_OP_279J39_124_314_n2738, div_DP_OP_279J39_124_314_n2737,
         div_DP_OP_279J39_124_314_n2736, div_DP_OP_279J39_124_314_n2735,
         div_DP_OP_279J39_124_314_n2734, div_DP_OP_279J39_124_314_n2733,
         div_DP_OP_279J39_124_314_n2732, div_DP_OP_279J39_124_314_n2731,
         div_DP_OP_279J39_124_314_n2730, div_DP_OP_279J39_124_314_n2729,
         div_DP_OP_279J39_124_314_n2728, div_DP_OP_279J39_124_314_n2727,
         div_DP_OP_279J39_124_314_n2726, div_DP_OP_279J39_124_314_n2725,
         div_DP_OP_279J39_124_314_n2724, div_DP_OP_279J39_124_314_n2723,
         div_DP_OP_279J39_124_314_n2722, div_DP_OP_279J39_124_314_n2721,
         div_DP_OP_279J39_124_314_n2720, div_DP_OP_279J39_124_314_n2719,
         div_DP_OP_279J39_124_314_n2718, div_DP_OP_279J39_124_314_n2717,
         div_DP_OP_279J39_124_314_n2716, div_DP_OP_279J39_124_314_n2715,
         div_DP_OP_279J39_124_314_n2714, div_DP_OP_279J39_124_314_n2713,
         div_DP_OP_279J39_124_314_n2712, div_DP_OP_279J39_124_314_n2711,
         div_DP_OP_279J39_124_314_n2710, div_DP_OP_279J39_124_314_n2709,
         div_DP_OP_279J39_124_314_n2708, div_DP_OP_279J39_124_314_n2707,
         div_DP_OP_279J39_124_314_n2706, div_DP_OP_279J39_124_314_n2705,
         div_DP_OP_279J39_124_314_n2704, div_DP_OP_279J39_124_314_n2703,
         div_DP_OP_279J39_124_314_n2702, div_DP_OP_279J39_124_314_n2701,
         div_DP_OP_279J39_124_314_n2700, div_DP_OP_279J39_124_314_n2699,
         div_DP_OP_279J39_124_314_n2698, div_DP_OP_279J39_124_314_n2697,
         div_DP_OP_279J39_124_314_n2696, div_DP_OP_279J39_124_314_n2695,
         div_DP_OP_279J39_124_314_n2694, div_DP_OP_279J39_124_314_n2693,
         div_DP_OP_279J39_124_314_n2692, div_DP_OP_279J39_124_314_n2691,
         div_DP_OP_279J39_124_314_n2690, div_DP_OP_279J39_124_314_n2689,
         div_DP_OP_279J39_124_314_n2688, div_DP_OP_279J39_124_314_n2687,
         div_DP_OP_279J39_124_314_n2686, div_DP_OP_279J39_124_314_n2685,
         div_DP_OP_279J39_124_314_n2684, div_DP_OP_279J39_124_314_n2683,
         div_DP_OP_279J39_124_314_n2682, div_DP_OP_279J39_124_314_n2681,
         div_DP_OP_279J39_124_314_n2680, div_DP_OP_279J39_124_314_n2679,
         div_DP_OP_279J39_124_314_n2678, div_DP_OP_279J39_124_314_n2677,
         div_DP_OP_279J39_124_314_n2676, div_DP_OP_279J39_124_314_n2675,
         div_DP_OP_279J39_124_314_n2674, div_DP_OP_279J39_124_314_n2673,
         div_DP_OP_279J39_124_314_n2672, div_DP_OP_279J39_124_314_n2671,
         div_DP_OP_279J39_124_314_n2670, div_DP_OP_279J39_124_314_n2669,
         div_DP_OP_279J39_124_314_n2668, div_DP_OP_279J39_124_314_n2667,
         div_DP_OP_279J39_124_314_n2666, div_DP_OP_279J39_124_314_n2665,
         div_DP_OP_279J39_124_314_n2664, div_DP_OP_279J39_124_314_n2663,
         div_DP_OP_279J39_124_314_n2662, div_DP_OP_279J39_124_314_n2661,
         div_DP_OP_279J39_124_314_n2660, div_DP_OP_279J39_124_314_n2659,
         div_DP_OP_279J39_124_314_n2658, div_DP_OP_279J39_124_314_n2657,
         div_DP_OP_279J39_124_314_n2656, div_DP_OP_279J39_124_314_n2655,
         div_DP_OP_279J39_124_314_n2654, div_DP_OP_279J39_124_314_n2653,
         div_DP_OP_279J39_124_314_n2652, div_DP_OP_279J39_124_314_n2651,
         div_DP_OP_279J39_124_314_n2650, div_DP_OP_279J39_124_314_n2649,
         div_DP_OP_279J39_124_314_n2648, div_DP_OP_279J39_124_314_n2647,
         div_DP_OP_279J39_124_314_n2646, div_DP_OP_279J39_124_314_n2645,
         div_DP_OP_279J39_124_314_n2644, div_DP_OP_279J39_124_314_n2643,
         div_DP_OP_279J39_124_314_n2642, div_DP_OP_279J39_124_314_n2641,
         div_DP_OP_279J39_124_314_n2640, div_DP_OP_279J39_124_314_n2639,
         div_DP_OP_279J39_124_314_n2638, div_DP_OP_279J39_124_314_n2637,
         div_DP_OP_279J39_124_314_n2636, div_DP_OP_279J39_124_314_n2635,
         div_DP_OP_279J39_124_314_n2634, div_DP_OP_279J39_124_314_n2633,
         div_DP_OP_279J39_124_314_n2632, div_DP_OP_279J39_124_314_n2631,
         div_DP_OP_279J39_124_314_n2630, div_DP_OP_279J39_124_314_n2629,
         div_DP_OP_279J39_124_314_n2628, div_DP_OP_279J39_124_314_n2627,
         div_DP_OP_279J39_124_314_n2626, div_DP_OP_279J39_124_314_n2625,
         div_DP_OP_279J39_124_314_n2624, div_DP_OP_279J39_124_314_n2623,
         div_DP_OP_279J39_124_314_n2622, div_DP_OP_279J39_124_314_n2621,
         div_DP_OP_279J39_124_314_n2620, div_DP_OP_279J39_124_314_n2619,
         div_DP_OP_279J39_124_314_n2618, div_DP_OP_279J39_124_314_n2617,
         div_DP_OP_279J39_124_314_n2616, div_DP_OP_279J39_124_314_n2615,
         div_DP_OP_279J39_124_314_n2614, div_DP_OP_279J39_124_314_n2613,
         div_DP_OP_279J39_124_314_n2612, div_DP_OP_279J39_124_314_n2611,
         div_DP_OP_279J39_124_314_n2610, div_DP_OP_279J39_124_314_n2609,
         div_DP_OP_279J39_124_314_n2608, div_DP_OP_279J39_124_314_n2607,
         div_DP_OP_279J39_124_314_n2606, div_DP_OP_279J39_124_314_n2605,
         div_DP_OP_279J39_124_314_n2604, div_DP_OP_279J39_124_314_n2603,
         div_DP_OP_279J39_124_314_n2602, div_DP_OP_279J39_124_314_n2601,
         div_DP_OP_279J39_124_314_n2600, div_DP_OP_279J39_124_314_n2599,
         div_DP_OP_279J39_124_314_n2598, div_DP_OP_279J39_124_314_n2597,
         div_DP_OP_279J39_124_314_n2596, div_DP_OP_279J39_124_314_n2595,
         div_DP_OP_279J39_124_314_n2594, div_DP_OP_279J39_124_314_n2593,
         div_DP_OP_279J39_124_314_n2592, div_DP_OP_279J39_124_314_n2591,
         div_DP_OP_279J39_124_314_n2590, div_DP_OP_279J39_124_314_n2589,
         div_DP_OP_279J39_124_314_n2588, div_DP_OP_279J39_124_314_n2587,
         div_DP_OP_279J39_124_314_n2586, div_DP_OP_279J39_124_314_n2585,
         div_DP_OP_279J39_124_314_n2584, div_DP_OP_279J39_124_314_n2583,
         div_DP_OP_279J39_124_314_n2582, div_DP_OP_279J39_124_314_n2581,
         div_DP_OP_279J39_124_314_n2580, div_DP_OP_279J39_124_314_n2579,
         div_DP_OP_279J39_124_314_n2578, div_DP_OP_279J39_124_314_n2577,
         div_DP_OP_279J39_124_314_n2576, div_DP_OP_279J39_124_314_n2575,
         div_DP_OP_279J39_124_314_n2574, div_DP_OP_279J39_124_314_n2573,
         div_DP_OP_279J39_124_314_n2572, div_DP_OP_279J39_124_314_n2571,
         div_DP_OP_279J39_124_314_n2570, div_DP_OP_279J39_124_314_n2569,
         div_DP_OP_279J39_124_314_n2568, div_DP_OP_279J39_124_314_n2567,
         div_DP_OP_279J39_124_314_n2566, div_DP_OP_279J39_124_314_n2565,
         div_DP_OP_279J39_124_314_n2564, div_DP_OP_279J39_124_314_n2563,
         div_DP_OP_279J39_124_314_n2562, div_DP_OP_279J39_124_314_n2561,
         div_DP_OP_279J39_124_314_n2560, div_DP_OP_279J39_124_314_n2559,
         div_DP_OP_279J39_124_314_n2558, div_DP_OP_279J39_124_314_n2557,
         div_DP_OP_279J39_124_314_n2556, div_DP_OP_279J39_124_314_n2555,
         div_DP_OP_279J39_124_314_n2554, div_DP_OP_279J39_124_314_n2553,
         div_DP_OP_279J39_124_314_n2552, div_DP_OP_279J39_124_314_n2551,
         div_DP_OP_279J39_124_314_n2550, div_DP_OP_279J39_124_314_n2549,
         div_DP_OP_279J39_124_314_n2547, div_DP_OP_279J39_124_314_n2546,
         div_DP_OP_279J39_124_314_n2545, div_DP_OP_279J39_124_314_n2544,
         div_DP_OP_279J39_124_314_n2543, div_DP_OP_279J39_124_314_n2542,
         div_DP_OP_279J39_124_314_n2541, div_DP_OP_279J39_124_314_n2539,
         div_DP_OP_279J39_124_314_n2538, div_DP_OP_279J39_124_314_n2537,
         div_DP_OP_279J39_124_314_n2536, div_DP_OP_279J39_124_314_n2535,
         div_DP_OP_279J39_124_314_n2534, div_DP_OP_279J39_124_314_n2533,
         div_DP_OP_279J39_124_314_n2532, div_DP_OP_279J39_124_314_n2530,
         div_DP_OP_279J39_124_314_n2529, div_DP_OP_279J39_124_314_n2528,
         div_DP_OP_279J39_124_314_n2527, div_DP_OP_279J39_124_314_n2235,
         div_DP_OP_279J39_124_314_n2234, div_DP_OP_279J39_124_314_n2233,
         div_DP_OP_279J39_124_314_n2232, div_DP_OP_279J39_124_314_n2231,
         div_DP_OP_279J39_124_314_n2230, div_DP_OP_279J39_124_314_n2229,
         div_DP_OP_279J39_124_314_n2228, div_DP_OP_279J39_124_314_n2227,
         div_DP_OP_279J39_124_314_n2226, div_DP_OP_279J39_124_314_n2225,
         div_DP_OP_279J39_124_314_n2224, div_DP_OP_279J39_124_314_n2223,
         div_DP_OP_279J39_124_314_n2222, div_DP_OP_279J39_124_314_n2221,
         div_DP_OP_279J39_124_314_n2220, div_DP_OP_279J39_124_314_n2219,
         div_DP_OP_279J39_124_314_n2218, div_DP_OP_279J39_124_314_n2217,
         div_DP_OP_279J39_124_314_n2216, div_DP_OP_279J39_124_314_n2215,
         div_DP_OP_279J39_124_314_n2214, div_DP_OP_279J39_124_314_n2213,
         div_DP_OP_279J39_124_314_n2212, div_DP_OP_279J39_124_314_n2211,
         div_DP_OP_279J39_124_314_n2210, div_DP_OP_279J39_124_314_n2209,
         div_DP_OP_279J39_124_314_n2208, div_DP_OP_279J39_124_314_n2207,
         div_DP_OP_279J39_124_314_n2206, div_DP_OP_279J39_124_314_n2205,
         div_DP_OP_279J39_124_314_n2204, div_DP_OP_279J39_124_314_n2203,
         div_DP_OP_279J39_124_314_n2202, div_DP_OP_279J39_124_314_n2201,
         div_DP_OP_279J39_124_314_n2200, div_DP_OP_279J39_124_314_n2199,
         div_DP_OP_279J39_124_314_n2198, div_DP_OP_279J39_124_314_n2197,
         div_DP_OP_279J39_124_314_n2196, div_DP_OP_279J39_124_314_n2195,
         div_DP_OP_279J39_124_314_n2194, div_DP_OP_279J39_124_314_n2193,
         div_DP_OP_279J39_124_314_n2192, div_DP_OP_279J39_124_314_n2191,
         div_DP_OP_279J39_124_314_n2190, div_DP_OP_279J39_124_314_n2189,
         div_DP_OP_279J39_124_314_n2188, div_DP_OP_279J39_124_314_n2187,
         div_DP_OP_279J39_124_314_n2186, div_DP_OP_279J39_124_314_n2185,
         div_DP_OP_279J39_124_314_n2184, div_DP_OP_279J39_124_314_n2183,
         div_DP_OP_279J39_124_314_n2182, div_DP_OP_279J39_124_314_n2181,
         div_DP_OP_279J39_124_314_n2180, div_DP_OP_279J39_124_314_n2179,
         div_DP_OP_279J39_124_314_n2178, div_DP_OP_279J39_124_314_n2177,
         div_DP_OP_279J39_124_314_n2176, div_DP_OP_279J39_124_314_n2175,
         div_DP_OP_279J39_124_314_n2174, div_DP_OP_279J39_124_314_n2173,
         div_DP_OP_279J39_124_314_n2172, div_DP_OP_279J39_124_314_n2171,
         div_DP_OP_279J39_124_314_n2170, div_DP_OP_279J39_124_314_n2169,
         div_DP_OP_279J39_124_314_n2168, div_DP_OP_279J39_124_314_n2167,
         div_DP_OP_279J39_124_314_n2166, div_DP_OP_279J39_124_314_n2165,
         div_DP_OP_279J39_124_314_n2164, div_DP_OP_279J39_124_314_n2163,
         div_DP_OP_279J39_124_314_n2162, div_DP_OP_279J39_124_314_n2161,
         div_DP_OP_279J39_124_314_n2160, div_DP_OP_279J39_124_314_n2159,
         div_DP_OP_279J39_124_314_n2158, div_DP_OP_279J39_124_314_n2157,
         div_DP_OP_279J39_124_314_n2156, div_DP_OP_279J39_124_314_n2155,
         div_DP_OP_279J39_124_314_n2154, div_DP_OP_279J39_124_314_n2153,
         div_DP_OP_279J39_124_314_n2152, div_DP_OP_279J39_124_314_n2151,
         div_DP_OP_279J39_124_314_n2150, div_DP_OP_279J39_124_314_n2149,
         div_DP_OP_279J39_124_314_n2148, div_DP_OP_279J39_124_314_n2147,
         div_DP_OP_279J39_124_314_n2146, div_DP_OP_279J39_124_314_n2145,
         div_DP_OP_279J39_124_314_n2144, div_DP_OP_279J39_124_314_n2143,
         div_DP_OP_279J39_124_314_n2142, div_DP_OP_279J39_124_314_n2141,
         div_DP_OP_279J39_124_314_n2140, div_DP_OP_279J39_124_314_n2139,
         div_DP_OP_279J39_124_314_n2138, div_DP_OP_279J39_124_314_n2137,
         div_DP_OP_279J39_124_314_n2136, div_DP_OP_279J39_124_314_n2135,
         div_DP_OP_279J39_124_314_n2134, div_DP_OP_279J39_124_314_n2133,
         div_DP_OP_279J39_124_314_n2132, div_DP_OP_279J39_124_314_n2131,
         div_DP_OP_279J39_124_314_n2130, div_DP_OP_279J39_124_314_n2129,
         div_DP_OP_279J39_124_314_n2128, div_DP_OP_279J39_124_314_n2127,
         div_DP_OP_279J39_124_314_n2126, div_DP_OP_279J39_124_314_n2125,
         div_DP_OP_279J39_124_314_n2124, div_DP_OP_279J39_124_314_n2123,
         div_DP_OP_279J39_124_314_n2122, div_DP_OP_279J39_124_314_n2121,
         div_DP_OP_279J39_124_314_n2120, div_DP_OP_279J39_124_314_n2119,
         div_DP_OP_279J39_124_314_n2118, div_DP_OP_279J39_124_314_n2117,
         div_DP_OP_279J39_124_314_n2116, div_DP_OP_279J39_124_314_n2115,
         div_DP_OP_279J39_124_314_n2114, div_DP_OP_279J39_124_314_n2113,
         div_DP_OP_279J39_124_314_n2112, div_DP_OP_279J39_124_314_n2111,
         div_DP_OP_279J39_124_314_n2110, div_DP_OP_279J39_124_314_n2109,
         div_DP_OP_279J39_124_314_n2108, div_DP_OP_279J39_124_314_n2107,
         div_DP_OP_279J39_124_314_n2106, div_DP_OP_279J39_124_314_n2105,
         div_DP_OP_279J39_124_314_n2104, div_DP_OP_279J39_124_314_n2103,
         div_DP_OP_279J39_124_314_n2102, div_DP_OP_279J39_124_314_n2101,
         div_DP_OP_279J39_124_314_n2100, div_DP_OP_279J39_124_314_n2099,
         div_DP_OP_279J39_124_314_n2098, div_DP_OP_279J39_124_314_n2097,
         div_DP_OP_279J39_124_314_n2096, div_DP_OP_279J39_124_314_n2095,
         div_DP_OP_279J39_124_314_n2094, div_DP_OP_279J39_124_314_n2093,
         div_DP_OP_279J39_124_314_n2092, div_DP_OP_279J39_124_314_n2091,
         div_DP_OP_279J39_124_314_n2090, div_DP_OP_279J39_124_314_n2089,
         div_DP_OP_279J39_124_314_n2088, div_DP_OP_279J39_124_314_n2087,
         div_DP_OP_279J39_124_314_n2086, div_DP_OP_279J39_124_314_n2085,
         div_DP_OP_279J39_124_314_n2084, div_DP_OP_279J39_124_314_n2083,
         div_DP_OP_279J39_124_314_n2082, div_DP_OP_279J39_124_314_n2081,
         div_DP_OP_279J39_124_314_n2080, div_DP_OP_279J39_124_314_n2079,
         div_DP_OP_279J39_124_314_n2078, div_DP_OP_279J39_124_314_n2077,
         div_DP_OP_279J39_124_314_n2076, div_DP_OP_279J39_124_314_n2075,
         div_DP_OP_279J39_124_314_n2074, div_DP_OP_279J39_124_314_n2073,
         div_DP_OP_279J39_124_314_n2072, div_DP_OP_279J39_124_314_n2071,
         div_DP_OP_279J39_124_314_n2070, div_DP_OP_279J39_124_314_n2069,
         div_DP_OP_279J39_124_314_n2068, div_DP_OP_279J39_124_314_n2067,
         div_DP_OP_279J39_124_314_n2066, div_DP_OP_279J39_124_314_n2065,
         div_DP_OP_279J39_124_314_n2064, div_DP_OP_279J39_124_314_n2063,
         div_DP_OP_279J39_124_314_n2062, div_DP_OP_279J39_124_314_n2061,
         div_DP_OP_279J39_124_314_n2060, div_DP_OP_279J39_124_314_n2059,
         div_DP_OP_279J39_124_314_n2058, div_DP_OP_279J39_124_314_n2057,
         div_DP_OP_279J39_124_314_n2056, div_DP_OP_279J39_124_314_n2055,
         div_DP_OP_279J39_124_314_n2054, div_DP_OP_279J39_124_314_n2053,
         div_DP_OP_279J39_124_314_n2052, div_DP_OP_279J39_124_314_n2051,
         div_DP_OP_279J39_124_314_n2050, div_DP_OP_279J39_124_314_n2049,
         div_DP_OP_279J39_124_314_n2048, div_DP_OP_279J39_124_314_n2047,
         div_DP_OP_279J39_124_314_n2046, div_DP_OP_279J39_124_314_n2045,
         div_DP_OP_279J39_124_314_n2044, div_DP_OP_279J39_124_314_n2043,
         div_DP_OP_279J39_124_314_n2042, div_DP_OP_279J39_124_314_n2041,
         div_DP_OP_279J39_124_314_n2040, div_DP_OP_279J39_124_314_n2039,
         div_DP_OP_279J39_124_314_n2038, div_DP_OP_279J39_124_314_n2037,
         div_DP_OP_279J39_124_314_n2036, div_DP_OP_279J39_124_314_n2035,
         div_DP_OP_279J39_124_314_n2034, div_DP_OP_279J39_124_314_n2033,
         div_DP_OP_279J39_124_314_n2032, div_DP_OP_279J39_124_314_n2031,
         div_DP_OP_279J39_124_314_n2030, div_DP_OP_279J39_124_314_n2029,
         div_DP_OP_279J39_124_314_n2028, div_DP_OP_279J39_124_314_n2027,
         div_DP_OP_279J39_124_314_n2026, div_DP_OP_279J39_124_314_n2025,
         div_DP_OP_279J39_124_314_n2024, div_DP_OP_279J39_124_314_n2023,
         div_DP_OP_279J39_124_314_n2022, div_DP_OP_279J39_124_314_n2021,
         div_DP_OP_279J39_124_314_n2020, div_DP_OP_279J39_124_314_n2019,
         div_DP_OP_279J39_124_314_n2018, div_DP_OP_279J39_124_314_n2017,
         div_DP_OP_279J39_124_314_n2016, div_DP_OP_279J39_124_314_n2015,
         div_DP_OP_279J39_124_314_n2014, div_DP_OP_279J39_124_314_n2013,
         div_DP_OP_279J39_124_314_n2012, div_DP_OP_279J39_124_314_n2011,
         div_DP_OP_279J39_124_314_n2010, div_DP_OP_279J39_124_314_n2009,
         div_DP_OP_279J39_124_314_n2008, div_DP_OP_279J39_124_314_n2007,
         div_DP_OP_279J39_124_314_n2006, div_DP_OP_279J39_124_314_n2005,
         div_DP_OP_279J39_124_314_n2004, div_DP_OP_279J39_124_314_n2003,
         div_DP_OP_279J39_124_314_n2002, div_DP_OP_279J39_124_314_n2001,
         div_DP_OP_279J39_124_314_n2000, div_DP_OP_279J39_124_314_n1999,
         div_DP_OP_279J39_124_314_n1998, div_DP_OP_279J39_124_314_n1997,
         div_DP_OP_279J39_124_314_n1996, div_DP_OP_279J39_124_314_n1995,
         div_DP_OP_279J39_124_314_n1994, div_DP_OP_279J39_124_314_n1993,
         div_DP_OP_279J39_124_314_n1992, div_DP_OP_279J39_124_314_n1991,
         div_DP_OP_279J39_124_314_n1990, div_DP_OP_279J39_124_314_n1989,
         div_DP_OP_279J39_124_314_n1988, div_DP_OP_279J39_124_314_n1987,
         div_DP_OP_279J39_124_314_n1986, div_DP_OP_279J39_124_314_n1985,
         div_DP_OP_279J39_124_314_n1984, div_DP_OP_279J39_124_314_n1983,
         div_DP_OP_279J39_124_314_n1982, div_DP_OP_279J39_124_314_n1981,
         div_DP_OP_279J39_124_314_n1980, div_DP_OP_279J39_124_314_n1979,
         div_DP_OP_279J39_124_314_n1978, div_DP_OP_279J39_124_314_n1977,
         div_DP_OP_279J39_124_314_n1976, div_DP_OP_279J39_124_314_n1975,
         div_DP_OP_279J39_124_314_n1974, div_DP_OP_279J39_124_314_n1973,
         div_DP_OP_279J39_124_314_n1972, div_DP_OP_279J39_124_314_n1971,
         div_DP_OP_279J39_124_314_n1970, div_DP_OP_279J39_124_314_n1969,
         div_DP_OP_279J39_124_314_n1968, div_DP_OP_279J39_124_314_n1967,
         div_DP_OP_279J39_124_314_n1966, div_DP_OP_279J39_124_314_n1965,
         div_DP_OP_279J39_124_314_n1964, div_DP_OP_279J39_124_314_n1963,
         div_DP_OP_279J39_124_314_n1962, div_DP_OP_279J39_124_314_n1961,
         div_DP_OP_279J39_124_314_n1960, div_DP_OP_279J39_124_314_n1959,
         div_DP_OP_279J39_124_314_n1958, div_DP_OP_279J39_124_314_n1957,
         div_DP_OP_279J39_124_314_n1956, div_DP_OP_279J39_124_314_n1955,
         div_DP_OP_279J39_124_314_n1954, div_DP_OP_279J39_124_314_n1953,
         div_DP_OP_279J39_124_314_n1952, div_DP_OP_279J39_124_314_n1951,
         div_DP_OP_279J39_124_314_n1950, div_DP_OP_279J39_124_314_n1949,
         div_DP_OP_279J39_124_314_n1948, div_DP_OP_279J39_124_314_n1947,
         div_DP_OP_279J39_124_314_n1946, div_DP_OP_279J39_124_314_n1945,
         div_DP_OP_279J39_124_314_n1944, div_DP_OP_279J39_124_314_n1943,
         div_DP_OP_279J39_124_314_n1942, div_DP_OP_279J39_124_314_n1941,
         div_DP_OP_279J39_124_314_n1940, div_DP_OP_279J39_124_314_n1939,
         div_DP_OP_279J39_124_314_n1938, div_DP_OP_279J39_124_314_n1937,
         div_DP_OP_279J39_124_314_n1936, div_DP_OP_279J39_124_314_n1935,
         div_DP_OP_279J39_124_314_n1934, div_DP_OP_279J39_124_314_n1933,
         div_DP_OP_279J39_124_314_n1932, div_DP_OP_279J39_124_314_n1931,
         div_DP_OP_279J39_124_314_n1930, div_DP_OP_279J39_124_314_n1929,
         div_DP_OP_279J39_124_314_n1928, div_DP_OP_279J39_124_314_n1927,
         div_DP_OP_279J39_124_314_n1926, div_DP_OP_279J39_124_314_n1925,
         div_DP_OP_279J39_124_314_n1924, div_DP_OP_279J39_124_314_n1923,
         div_DP_OP_279J39_124_314_n1922, div_DP_OP_279J39_124_314_n1921,
         div_DP_OP_279J39_124_314_n1920, div_DP_OP_279J39_124_314_n1919,
         div_DP_OP_279J39_124_314_n1918, div_DP_OP_279J39_124_314_n1917,
         div_DP_OP_279J39_124_314_n1916, div_DP_OP_279J39_124_314_n1915,
         div_DP_OP_279J39_124_314_n1914, div_DP_OP_279J39_124_314_n1913,
         div_DP_OP_279J39_124_314_n1912, div_DP_OP_279J39_124_314_n1911,
         div_DP_OP_279J39_124_314_n1910, div_DP_OP_279J39_124_314_n1909,
         div_DP_OP_279J39_124_314_n1908, div_DP_OP_279J39_124_314_n1907,
         div_DP_OP_279J39_124_314_n1906, div_DP_OP_279J39_124_314_n1905,
         div_DP_OP_279J39_124_314_n1904, div_DP_OP_279J39_124_314_n1903,
         div_DP_OP_279J39_124_314_n1902, div_DP_OP_279J39_124_314_n1901,
         div_DP_OP_279J39_124_314_n1900, div_DP_OP_279J39_124_314_n1899,
         div_DP_OP_279J39_124_314_n1898, div_DP_OP_279J39_124_314_n1897,
         div_DP_OP_279J39_124_314_n1896, div_DP_OP_279J39_124_314_n1895,
         div_DP_OP_279J39_124_314_n1894, div_DP_OP_279J39_124_314_n1893,
         div_DP_OP_279J39_124_314_n1892, div_DP_OP_279J39_124_314_n1891,
         div_DP_OP_279J39_124_314_n1890, div_DP_OP_279J39_124_314_n1889,
         div_DP_OP_279J39_124_314_n1888, div_DP_OP_279J39_124_314_n1887,
         div_DP_OP_279J39_124_314_n1886, div_DP_OP_279J39_124_314_n1885,
         div_DP_OP_279J39_124_314_n1884, div_DP_OP_279J39_124_314_n1883,
         div_DP_OP_279J39_124_314_n1882, div_DP_OP_279J39_124_314_n1881,
         div_DP_OP_279J39_124_314_n1880, div_DP_OP_279J39_124_314_n1879,
         div_DP_OP_279J39_124_314_n1878, div_DP_OP_279J39_124_314_n1877,
         div_DP_OP_279J39_124_314_n1876, div_DP_OP_279J39_124_314_n1875,
         div_DP_OP_279J39_124_314_n1874, div_DP_OP_279J39_124_314_n1873,
         div_DP_OP_279J39_124_314_n1872, div_DP_OP_279J39_124_314_n1871,
         div_DP_OP_279J39_124_314_n1870, div_DP_OP_279J39_124_314_n1869,
         div_DP_OP_279J39_124_314_n1868, div_DP_OP_279J39_124_314_n1867,
         div_DP_OP_279J39_124_314_n1866, div_DP_OP_279J39_124_314_n1865,
         div_DP_OP_279J39_124_314_n1864, div_DP_OP_279J39_124_314_n1863,
         div_DP_OP_279J39_124_314_n1862, div_DP_OP_279J39_124_314_n1861,
         div_DP_OP_279J39_124_314_n1860, div_DP_OP_279J39_124_314_n1859,
         div_DP_OP_279J39_124_314_n1858, div_DP_OP_279J39_124_314_n1857,
         div_DP_OP_279J39_124_314_n1856, div_DP_OP_279J39_124_314_n1855,
         div_DP_OP_279J39_124_314_n1854, div_DP_OP_279J39_124_314_n1853,
         div_DP_OP_279J39_124_314_n1852, div_DP_OP_279J39_124_314_n1851,
         div_DP_OP_279J39_124_314_n1850, div_DP_OP_279J39_124_314_n1849,
         div_DP_OP_279J39_124_314_n1848, div_DP_OP_279J39_124_314_n1847,
         div_DP_OP_279J39_124_314_n1846, div_DP_OP_279J39_124_314_n1845,
         div_DP_OP_279J39_124_314_n1844, div_DP_OP_279J39_124_314_n1843,
         div_DP_OP_279J39_124_314_n1842, div_DP_OP_279J39_124_314_n1841,
         div_DP_OP_279J39_124_314_n1840, div_DP_OP_279J39_124_314_n1839,
         div_DP_OP_279J39_124_314_n1838, div_DP_OP_279J39_124_314_n1837,
         div_DP_OP_279J39_124_314_n1836, div_DP_OP_279J39_124_314_n1835,
         div_DP_OP_279J39_124_314_n1834, div_DP_OP_279J39_124_314_n1833,
         div_DP_OP_279J39_124_314_n1832, div_DP_OP_279J39_124_314_n1831,
         div_DP_OP_279J39_124_314_n1830, div_DP_OP_279J39_124_314_n1829,
         div_DP_OP_279J39_124_314_n1828, div_DP_OP_279J39_124_314_n1827,
         div_DP_OP_279J39_124_314_n1826, div_DP_OP_279J39_124_314_n1825,
         div_DP_OP_279J39_124_314_n1824, div_DP_OP_279J39_124_314_n1823,
         div_DP_OP_279J39_124_314_n1822, div_DP_OP_279J39_124_314_n1821,
         div_DP_OP_279J39_124_314_n1820, div_DP_OP_279J39_124_314_n1819,
         div_DP_OP_279J39_124_314_n1818, div_DP_OP_279J39_124_314_n1817,
         div_DP_OP_279J39_124_314_n1816, div_DP_OP_279J39_124_314_n1815,
         div_DP_OP_279J39_124_314_n1814, div_DP_OP_279J39_124_314_n1813,
         div_DP_OP_279J39_124_314_n1812, div_DP_OP_279J39_124_314_n1811,
         div_DP_OP_279J39_124_314_n1810, div_DP_OP_279J39_124_314_n1809,
         div_DP_OP_279J39_124_314_n1808, div_DP_OP_279J39_124_314_n1807,
         div_DP_OP_279J39_124_314_n1806, div_DP_OP_279J39_124_314_n1805,
         div_DP_OP_279J39_124_314_n1804, div_DP_OP_279J39_124_314_n1803,
         div_DP_OP_279J39_124_314_n1802, div_DP_OP_279J39_124_314_n1801,
         div_DP_OP_279J39_124_314_n1800, div_DP_OP_279J39_124_314_n1799,
         div_DP_OP_279J39_124_314_n1798, div_DP_OP_279J39_124_314_n1797,
         div_DP_OP_279J39_124_314_n1796, div_DP_OP_279J39_124_314_n1795,
         div_DP_OP_279J39_124_314_n1794, div_DP_OP_279J39_124_314_n1793,
         div_DP_OP_279J39_124_314_n1792, div_DP_OP_279J39_124_314_n1791,
         div_DP_OP_279J39_124_314_n1790, div_DP_OP_279J39_124_314_n1789,
         div_DP_OP_279J39_124_314_n1788, div_DP_OP_279J39_124_314_n1787,
         div_DP_OP_279J39_124_314_n1786, div_DP_OP_279J39_124_314_n1785,
         div_DP_OP_279J39_124_314_n1784, div_DP_OP_279J39_124_314_n1783,
         div_DP_OP_279J39_124_314_n1782, div_DP_OP_279J39_124_314_n1781,
         div_DP_OP_279J39_124_314_n1780, div_DP_OP_279J39_124_314_n1779,
         div_DP_OP_279J39_124_314_n1778, div_DP_OP_279J39_124_314_n1777,
         div_DP_OP_279J39_124_314_n1776, div_DP_OP_279J39_124_314_n1775,
         div_DP_OP_279J39_124_314_n1774, div_DP_OP_279J39_124_314_n1773,
         div_DP_OP_279J39_124_314_n1772, div_DP_OP_279J39_124_314_n1771,
         div_DP_OP_279J39_124_314_n1770, div_DP_OP_279J39_124_314_n1769,
         div_DP_OP_279J39_124_314_n1768, div_DP_OP_279J39_124_314_n1767,
         div_DP_OP_279J39_124_314_n1766, div_DP_OP_279J39_124_314_n1765,
         div_DP_OP_279J39_124_314_n1764, div_DP_OP_279J39_124_314_n1763,
         div_DP_OP_279J39_124_314_n1762, div_DP_OP_279J39_124_314_n1761,
         div_DP_OP_279J39_124_314_n1760, div_DP_OP_279J39_124_314_n1759,
         div_DP_OP_279J39_124_314_n1758, div_DP_OP_279J39_124_314_n1757,
         div_DP_OP_279J39_124_314_n1756, div_DP_OP_279J39_124_314_n1755,
         div_DP_OP_279J39_124_314_n1754, div_DP_OP_279J39_124_314_n1753,
         div_DP_OP_279J39_124_314_n1752, div_DP_OP_279J39_124_314_n1751,
         div_DP_OP_279J39_124_314_n1750, div_DP_OP_279J39_124_314_n1749,
         div_DP_OP_279J39_124_314_n1748, div_DP_OP_279J39_124_314_n1747,
         div_DP_OP_279J39_124_314_n1746, div_DP_OP_279J39_124_314_n1745,
         div_DP_OP_279J39_124_314_n1744, div_DP_OP_279J39_124_314_n1743,
         div_DP_OP_279J39_124_314_n1742, div_DP_OP_279J39_124_314_n1741,
         div_DP_OP_279J39_124_314_n1740, div_DP_OP_279J39_124_314_n1739,
         div_DP_OP_279J39_124_314_n1738, div_DP_OP_279J39_124_314_n1737,
         div_DP_OP_279J39_124_314_n1736, div_DP_OP_279J39_124_314_n1735,
         div_DP_OP_279J39_124_314_n1734, div_DP_OP_279J39_124_314_n1733,
         div_DP_OP_279J39_124_314_n1732, div_DP_OP_279J39_124_314_n1731,
         div_DP_OP_279J39_124_314_n1730, div_DP_OP_279J39_124_314_n1729,
         div_DP_OP_279J39_124_314_n1728, div_DP_OP_279J39_124_314_n1727,
         div_DP_OP_279J39_124_314_n1726, div_DP_OP_279J39_124_314_n1725,
         div_DP_OP_279J39_124_314_n1724, div_DP_OP_279J39_124_314_n1723,
         div_DP_OP_279J39_124_314_n1722, div_DP_OP_279J39_124_314_n1721,
         div_DP_OP_279J39_124_314_n1720, div_DP_OP_279J39_124_314_n1719,
         div_DP_OP_279J39_124_314_n1718, div_DP_OP_279J39_124_314_n1717,
         div_DP_OP_279J39_124_314_n1715, div_DP_OP_279J39_124_314_n1714,
         div_DP_OP_279J39_124_314_n1713, div_DP_OP_279J39_124_314_n1712,
         div_DP_OP_279J39_124_314_n1711, div_DP_OP_279J39_124_314_n1710,
         div_DP_OP_279J39_124_314_n1709, div_DP_OP_279J39_124_314_n1708,
         div_DP_OP_279J39_124_314_n1707, div_DP_OP_279J39_124_314_n1706,
         div_DP_OP_279J39_124_314_n1705, div_DP_OP_279J39_124_314_n1704,
         div_DP_OP_279J39_124_314_n1703, div_DP_OP_279J39_124_314_n1702,
         div_DP_OP_279J39_124_314_n1701, div_DP_OP_279J39_124_314_n1700,
         div_DP_OP_279J39_124_314_n1699, div_DP_OP_279J39_124_314_n1698,
         div_DP_OP_279J39_124_314_n1697, div_DP_OP_279J39_124_314_n1696,
         div_DP_OP_279J39_124_314_n1695, div_DP_OP_279J39_124_314_n1694,
         div_DP_OP_279J39_124_314_n1693, div_DP_OP_279J39_124_314_n1692,
         div_DP_OP_279J39_124_314_n1691, div_DP_OP_279J39_124_314_n1690,
         div_DP_OP_279J39_124_314_n1689, div_DP_OP_279J39_124_314_n1688,
         div_DP_OP_279J39_124_314_n1687, div_DP_OP_279J39_124_314_n1686,
         div_DP_OP_279J39_124_314_n1685, div_DP_OP_279J39_124_314_n1684,
         div_DP_OP_279J39_124_314_n1683, div_DP_OP_279J39_124_314_n1682,
         div_DP_OP_279J39_124_314_n1681, div_DP_OP_279J39_124_314_n1680,
         div_DP_OP_279J39_124_314_n1679, div_DP_OP_279J39_124_314_n1678,
         div_DP_OP_279J39_124_314_n1677, div_DP_OP_279J39_124_314_n1676,
         div_DP_OP_279J39_124_314_n1675, div_DP_OP_279J39_124_314_n1674,
         div_DP_OP_279J39_124_314_n1673, div_DP_OP_279J39_124_314_n1672,
         div_DP_OP_279J39_124_314_n1671, div_DP_OP_279J39_124_314_n1670,
         div_DP_OP_279J39_124_314_n1669, div_DP_OP_279J39_124_314_n1668,
         div_DP_OP_279J39_124_314_n1667, div_DP_OP_279J39_124_314_n1666,
         div_DP_OP_279J39_124_314_n1665, div_DP_OP_279J39_124_314_n1664,
         div_DP_OP_279J39_124_314_n1663, div_DP_OP_279J39_124_314_n1662,
         div_DP_OP_279J39_124_314_n1661, div_DP_OP_279J39_124_314_n1660,
         div_DP_OP_279J39_124_314_n1659, div_DP_OP_279J39_124_314_n1658,
         div_DP_OP_279J39_124_314_n1657, div_DP_OP_279J39_124_314_n1656,
         div_DP_OP_279J39_124_314_n1655, div_DP_OP_279J39_124_314_n1654,
         div_DP_OP_279J39_124_314_n1653, div_DP_OP_279J39_124_314_n1650,
         div_DP_OP_279J39_124_314_n1649, div_DP_OP_279J39_124_314_n1648,
         div_DP_OP_279J39_124_314_n1647, div_DP_OP_279J39_124_314_n1646,
         div_DP_OP_279J39_124_314_n1645, div_DP_OP_279J39_124_314_n1644,
         div_DP_OP_279J39_124_314_n1643, div_DP_OP_279J39_124_314_n1642,
         div_DP_OP_279J39_124_314_n1641, div_DP_OP_279J39_124_314_n1640,
         div_DP_OP_279J39_124_314_n1639, div_DP_OP_279J39_124_314_n1638,
         div_DP_OP_279J39_124_314_n1637, div_DP_OP_279J39_124_314_n1636,
         div_DP_OP_279J39_124_314_n1635, div_DP_OP_279J39_124_314_n1634,
         div_DP_OP_279J39_124_314_n1633, div_DP_OP_279J39_124_314_n1632,
         div_DP_OP_279J39_124_314_n1631, div_DP_OP_279J39_124_314_n1630,
         div_DP_OP_279J39_124_314_n1629, div_DP_OP_279J39_124_314_n1628,
         div_DP_OP_279J39_124_314_n1627, div_DP_OP_279J39_124_314_n1626,
         div_DP_OP_279J39_124_314_n1625, div_DP_OP_279J39_124_314_n1624,
         div_DP_OP_279J39_124_314_n1623, div_DP_OP_279J39_124_314_n1622,
         div_DP_OP_279J39_124_314_n1621, div_DP_OP_279J39_124_314_n1620,
         div_DP_OP_279J39_124_314_n1619, div_DP_OP_279J39_124_314_n1618,
         div_DP_OP_279J39_124_314_n1617, div_DP_OP_279J39_124_314_n1616,
         div_DP_OP_279J39_124_314_n1615, div_DP_OP_279J39_124_314_n1614,
         div_DP_OP_279J39_124_314_n1613, div_DP_OP_279J39_124_314_n1612,
         div_DP_OP_279J39_124_314_n1611, div_DP_OP_279J39_124_314_n1610,
         div_DP_OP_279J39_124_314_n1609, div_DP_OP_279J39_124_314_n1608,
         div_DP_OP_279J39_124_314_n1607, div_DP_OP_279J39_124_314_n1606,
         div_DP_OP_279J39_124_314_n1605, div_DP_OP_279J39_124_314_n1604,
         div_DP_OP_279J39_124_314_n1603, div_DP_OP_279J39_124_314_n1602,
         div_DP_OP_279J39_124_314_n1601, div_DP_OP_279J39_124_314_n1600,
         div_DP_OP_279J39_124_314_n1599, div_DP_OP_279J39_124_314_n1598,
         div_DP_OP_279J39_124_314_n1597, div_DP_OP_279J39_124_314_n1596,
         div_DP_OP_279J39_124_314_n1595, div_DP_OP_279J39_124_314_n1594,
         div_DP_OP_279J39_124_314_n1593, div_DP_OP_279J39_124_314_n1592,
         div_DP_OP_279J39_124_314_n1591, div_DP_OP_279J39_124_314_n1590,
         div_DP_OP_279J39_124_314_n1589, div_DP_OP_279J39_124_314_n1588,
         div_DP_OP_279J39_124_314_n1587, div_DP_OP_279J39_124_314_n1586,
         div_DP_OP_279J39_124_314_n1585, div_DP_OP_279J39_124_314_n1584,
         div_DP_OP_279J39_124_314_n1583, div_DP_OP_279J39_124_314_n1582,
         div_DP_OP_279J39_124_314_n1581, div_DP_OP_279J39_124_314_n1580,
         div_DP_OP_279J39_124_314_n1579, div_DP_OP_279J39_124_314_n1578,
         div_DP_OP_279J39_124_314_n1577, div_DP_OP_279J39_124_314_n1576,
         div_DP_OP_279J39_124_314_n1575, div_DP_OP_279J39_124_314_n1574,
         div_DP_OP_279J39_124_314_n1573, div_DP_OP_279J39_124_314_n1572,
         div_DP_OP_279J39_124_314_n1571, div_DP_OP_279J39_124_314_n1570,
         div_DP_OP_279J39_124_314_n1569, div_DP_OP_279J39_124_314_n1568,
         div_DP_OP_279J39_124_314_n1567, div_DP_OP_279J39_124_314_n1566,
         div_DP_OP_279J39_124_314_n1565, div_DP_OP_279J39_124_314_n1564,
         div_DP_OP_279J39_124_314_n1563, div_DP_OP_279J39_124_314_n1562,
         div_DP_OP_279J39_124_314_n1561, div_DP_OP_279J39_124_314_n1560,
         div_DP_OP_279J39_124_314_n1559, div_DP_OP_279J39_124_314_n1558,
         div_DP_OP_279J39_124_314_n1557, div_DP_OP_279J39_124_314_n1556,
         div_DP_OP_279J39_124_314_n1555, div_DP_OP_279J39_124_314_n1554,
         div_DP_OP_279J39_124_314_n1553, div_DP_OP_279J39_124_314_n1552,
         div_DP_OP_279J39_124_314_n1551, div_DP_OP_279J39_124_314_n1550,
         div_DP_OP_279J39_124_314_n1549, div_DP_OP_279J39_124_314_n1548,
         div_DP_OP_279J39_124_314_n1547, div_DP_OP_279J39_124_314_n1546,
         div_DP_OP_279J39_124_314_n1545, div_DP_OP_279J39_124_314_n1544,
         div_DP_OP_279J39_124_314_n1543, div_DP_OP_279J39_124_314_n1542,
         div_DP_OP_279J39_124_314_n1541, div_DP_OP_279J39_124_314_n1540,
         div_DP_OP_279J39_124_314_n1539, div_DP_OP_279J39_124_314_n1538,
         div_DP_OP_279J39_124_314_n1537, div_DP_OP_279J39_124_314_n1536,
         div_DP_OP_279J39_124_314_n1535, div_DP_OP_279J39_124_314_n1534,
         div_DP_OP_279J39_124_314_n1533, div_DP_OP_279J39_124_314_n1532,
         div_DP_OP_279J39_124_314_n1531, div_DP_OP_279J39_124_314_n1530,
         div_DP_OP_279J39_124_314_n1529, div_DP_OP_279J39_124_314_n1528,
         div_DP_OP_279J39_124_314_n1527, div_DP_OP_279J39_124_314_n1526,
         div_DP_OP_279J39_124_314_n1525, div_DP_OP_279J39_124_314_n1524,
         div_DP_OP_279J39_124_314_n1523, div_DP_OP_279J39_124_314_n1522,
         div_DP_OP_279J39_124_314_n1521, div_DP_OP_279J39_124_314_n1520,
         div_DP_OP_279J39_124_314_n1519, div_DP_OP_279J39_124_314_n1518,
         div_DP_OP_279J39_124_314_n1517, div_DP_OP_279J39_124_314_n1516,
         div_DP_OP_279J39_124_314_n1515, div_DP_OP_279J39_124_314_n1514,
         div_DP_OP_279J39_124_314_n1513, div_DP_OP_279J39_124_314_n1512,
         div_DP_OP_279J39_124_314_n1511, div_DP_OP_279J39_124_314_n1510,
         div_DP_OP_279J39_124_314_n1509, div_DP_OP_279J39_124_314_n1508,
         div_DP_OP_279J39_124_314_n1507, div_DP_OP_279J39_124_314_n1506,
         div_DP_OP_279J39_124_314_n1505, div_DP_OP_279J39_124_314_n1504,
         div_DP_OP_279J39_124_314_n1503, div_DP_OP_279J39_124_314_n1502,
         div_DP_OP_279J39_124_314_n1501, div_DP_OP_279J39_124_314_n1500,
         div_DP_OP_279J39_124_314_n1499, div_DP_OP_279J39_124_314_n1498,
         div_DP_OP_279J39_124_314_n1497, div_DP_OP_279J39_124_314_n1496,
         div_DP_OP_279J39_124_314_n1495, div_DP_OP_279J39_124_314_n1494,
         div_DP_OP_279J39_124_314_n1493, div_DP_OP_279J39_124_314_n1492,
         div_DP_OP_279J39_124_314_n1491, div_DP_OP_279J39_124_314_n1490,
         div_DP_OP_279J39_124_314_n1489, div_DP_OP_279J39_124_314_n1488,
         div_DP_OP_279J39_124_314_n1487, div_DP_OP_279J39_124_314_n1486,
         div_DP_OP_279J39_124_314_n1485, div_DP_OP_279J39_124_314_n1484,
         div_DP_OP_279J39_124_314_n1483, div_DP_OP_279J39_124_314_n1482,
         div_DP_OP_279J39_124_314_n1481, div_DP_OP_279J39_124_314_n1480,
         div_DP_OP_279J39_124_314_n1479, div_DP_OP_279J39_124_314_n1478,
         div_DP_OP_279J39_124_314_n1477, div_DP_OP_279J39_124_314_n1476,
         div_DP_OP_279J39_124_314_n1475, div_DP_OP_279J39_124_314_n1474,
         div_DP_OP_279J39_124_314_n1473, div_DP_OP_279J39_124_314_n1472,
         div_DP_OP_279J39_124_314_n1471, div_DP_OP_279J39_124_314_n1470,
         div_DP_OP_279J39_124_314_n1469, div_DP_OP_279J39_124_314_n1468,
         div_DP_OP_279J39_124_314_n1467, div_DP_OP_279J39_124_314_n1466,
         div_DP_OP_279J39_124_314_n1465, div_DP_OP_279J39_124_314_n1464,
         div_DP_OP_279J39_124_314_n1463, div_DP_OP_279J39_124_314_n1462,
         div_DP_OP_279J39_124_314_n1461, div_DP_OP_279J39_124_314_n1460,
         div_DP_OP_279J39_124_314_n1459, div_DP_OP_279J39_124_314_n1458,
         div_DP_OP_279J39_124_314_n1457, div_DP_OP_279J39_124_314_n1456,
         div_DP_OP_279J39_124_314_n1455, div_DP_OP_279J39_124_314_n1454,
         div_DP_OP_279J39_124_314_n1453, div_DP_OP_279J39_124_314_n1452,
         div_DP_OP_279J39_124_314_n1451, div_DP_OP_279J39_124_314_n1450,
         div_DP_OP_279J39_124_314_n1449, div_DP_OP_279J39_124_314_n1448,
         div_DP_OP_279J39_124_314_n1447, div_DP_OP_279J39_124_314_n1446,
         div_DP_OP_279J39_124_314_n1445, div_DP_OP_279J39_124_314_n1444,
         div_DP_OP_279J39_124_314_n1443, div_DP_OP_279J39_124_314_n1442,
         div_DP_OP_279J39_124_314_n1441, div_DP_OP_279J39_124_314_n1440,
         div_DP_OP_279J39_124_314_n1439, div_DP_OP_279J39_124_314_n1438,
         div_DP_OP_279J39_124_314_n1437, div_DP_OP_279J39_124_314_n1436,
         div_DP_OP_279J39_124_314_n1435, div_DP_OP_279J39_124_314_n1434,
         div_DP_OP_279J39_124_314_n1433, div_DP_OP_279J39_124_314_n1432,
         div_DP_OP_279J39_124_314_n1431, div_DP_OP_279J39_124_314_n1430,
         div_DP_OP_279J39_124_314_n1429, div_DP_OP_279J39_124_314_n1428,
         div_DP_OP_279J39_124_314_n1427, div_DP_OP_279J39_124_314_n1426,
         div_DP_OP_279J39_124_314_n1425, div_DP_OP_279J39_124_314_n1424,
         div_DP_OP_279J39_124_314_n1423, div_DP_OP_279J39_124_314_n1422,
         div_DP_OP_279J39_124_314_n1421, div_DP_OP_279J39_124_314_n1420,
         div_DP_OP_279J39_124_314_n1419, div_DP_OP_279J39_124_314_n1418,
         div_DP_OP_279J39_124_314_n1417, div_DP_OP_279J39_124_314_n1416,
         div_DP_OP_279J39_124_314_n1415, div_DP_OP_279J39_124_314_n1414,
         div_DP_OP_279J39_124_314_n1413, div_DP_OP_279J39_124_314_n1412,
         div_DP_OP_279J39_124_314_n1411, div_DP_OP_279J39_124_314_n1410,
         div_DP_OP_279J39_124_314_n1409, div_DP_OP_279J39_124_314_n1408,
         div_DP_OP_279J39_124_314_n1407, div_DP_OP_279J39_124_314_n1406,
         div_DP_OP_279J39_124_314_n1405, div_DP_OP_279J39_124_314_n1404,
         div_DP_OP_279J39_124_314_n1403, div_DP_OP_279J39_124_314_n1402,
         div_DP_OP_279J39_124_314_n1401, div_DP_OP_279J39_124_314_n1400,
         div_DP_OP_279J39_124_314_n1399, div_DP_OP_279J39_124_314_n1398,
         div_DP_OP_279J39_124_314_n1397, div_DP_OP_279J39_124_314_n1396,
         div_DP_OP_279J39_124_314_n1395, div_DP_OP_279J39_124_314_n1394,
         div_DP_OP_279J39_124_314_n1393, div_DP_OP_279J39_124_314_n1392,
         div_DP_OP_279J39_124_314_n1391, div_DP_OP_279J39_124_314_n1390,
         div_DP_OP_279J39_124_314_n1389, div_DP_OP_279J39_124_314_n1388,
         div_DP_OP_279J39_124_314_n1387, div_DP_OP_279J39_124_314_n1386,
         div_DP_OP_279J39_124_314_n1385, div_DP_OP_279J39_124_314_n1384,
         div_DP_OP_279J39_124_314_n1383, div_DP_OP_279J39_124_314_n1382,
         div_DP_OP_279J39_124_314_n1381, div_DP_OP_279J39_124_314_n1380,
         div_DP_OP_279J39_124_314_n1379, div_DP_OP_279J39_124_314_n1378,
         div_DP_OP_279J39_124_314_n1377, div_DP_OP_279J39_124_314_n1376,
         div_DP_OP_279J39_124_314_n1375, div_DP_OP_279J39_124_314_n1374,
         div_DP_OP_279J39_124_314_n1373, div_DP_OP_279J39_124_314_n1372,
         div_DP_OP_279J39_124_314_n1371, div_DP_OP_279J39_124_314_n1370,
         div_DP_OP_279J39_124_314_n1369, div_DP_OP_279J39_124_314_n1368,
         div_DP_OP_279J39_124_314_n1367, div_DP_OP_279J39_124_314_n1366,
         div_DP_OP_279J39_124_314_n1365, div_DP_OP_279J39_124_314_n1364,
         div_DP_OP_279J39_124_314_n1363, div_DP_OP_279J39_124_314_n1362,
         div_DP_OP_279J39_124_314_n1361, div_DP_OP_279J39_124_314_n1360,
         div_DP_OP_279J39_124_314_n1359, div_DP_OP_279J39_124_314_n1358,
         div_DP_OP_279J39_124_314_n1357, div_DP_OP_279J39_124_314_n1356,
         div_DP_OP_279J39_124_314_n1355, div_DP_OP_279J39_124_314_n1354,
         div_DP_OP_279J39_124_314_n1353, div_DP_OP_279J39_124_314_n1352,
         div_DP_OP_279J39_124_314_n1351, div_DP_OP_279J39_124_314_n1350,
         div_DP_OP_279J39_124_314_n1349, div_DP_OP_279J39_124_314_n1348,
         div_DP_OP_279J39_124_314_n1347, div_DP_OP_279J39_124_314_n1346,
         div_DP_OP_279J39_124_314_n1345, div_DP_OP_279J39_124_314_n1344,
         div_DP_OP_279J39_124_314_n1343, div_DP_OP_279J39_124_314_n1342,
         div_DP_OP_279J39_124_314_n1341, div_DP_OP_279J39_124_314_n1340,
         div_DP_OP_279J39_124_314_n1339, div_DP_OP_279J39_124_314_n1338,
         div_DP_OP_279J39_124_314_n1337, div_DP_OP_279J39_124_314_n1336,
         div_DP_OP_279J39_124_314_n1335, div_DP_OP_279J39_124_314_n1334,
         div_DP_OP_279J39_124_314_n1333, div_DP_OP_279J39_124_314_n1332,
         div_DP_OP_279J39_124_314_n1331, div_DP_OP_279J39_124_314_n1330,
         div_DP_OP_279J39_124_314_n1329, div_DP_OP_279J39_124_314_n1328,
         div_DP_OP_279J39_124_314_n1327, div_DP_OP_279J39_124_314_n1326,
         div_DP_OP_279J39_124_314_n1325, div_DP_OP_279J39_124_314_n1324,
         div_DP_OP_279J39_124_314_n1323, div_DP_OP_279J39_124_314_n1322,
         div_DP_OP_279J39_124_314_n1321, div_DP_OP_279J39_124_314_n1320,
         div_DP_OP_279J39_124_314_n1319, div_DP_OP_279J39_124_314_n1318,
         div_DP_OP_279J39_124_314_n1317, div_DP_OP_279J39_124_314_n1316,
         div_DP_OP_279J39_124_314_n1315, div_DP_OP_279J39_124_314_n1314,
         div_DP_OP_279J39_124_314_n1313, div_DP_OP_279J39_124_314_n1312,
         div_DP_OP_279J39_124_314_n1311, div_DP_OP_279J39_124_314_n1310,
         div_DP_OP_279J39_124_314_n1309, div_DP_OP_279J39_124_314_n1308,
         div_DP_OP_279J39_124_314_n1307, div_DP_OP_279J39_124_314_n1306,
         div_DP_OP_279J39_124_314_n1305, div_DP_OP_279J39_124_314_n1304,
         div_DP_OP_279J39_124_314_n1303, div_DP_OP_279J39_124_314_n1302,
         div_DP_OP_279J39_124_314_n1301, div_DP_OP_279J39_124_314_n1300,
         div_DP_OP_279J39_124_314_n1299, div_DP_OP_279J39_124_314_n1298,
         div_DP_OP_279J39_124_314_n1297, div_DP_OP_279J39_124_314_n1296,
         div_DP_OP_279J39_124_314_n1295, div_DP_OP_279J39_124_314_n1294,
         div_DP_OP_279J39_124_314_n1293, div_DP_OP_279J39_124_314_n1292,
         div_DP_OP_279J39_124_314_n1291, div_DP_OP_279J39_124_314_n1290,
         div_DP_OP_279J39_124_314_n1289, div_DP_OP_279J39_124_314_n1288,
         div_DP_OP_279J39_124_314_n1287, div_DP_OP_279J39_124_314_n1286,
         div_DP_OP_279J39_124_314_n1285, div_DP_OP_279J39_124_314_n1284,
         div_DP_OP_279J39_124_314_n1283, div_DP_OP_279J39_124_314_n1282,
         div_DP_OP_279J39_124_314_n1281, div_DP_OP_279J39_124_314_n1280,
         div_DP_OP_279J39_124_314_n1279, div_DP_OP_279J39_124_314_n1278,
         div_DP_OP_279J39_124_314_n1277, div_DP_OP_279J39_124_314_n1276,
         div_DP_OP_279J39_124_314_n1275, div_DP_OP_279J39_124_314_n1274,
         div_DP_OP_279J39_124_314_n1273, div_DP_OP_279J39_124_314_n1272,
         div_DP_OP_279J39_124_314_n1271, div_DP_OP_279J39_124_314_n1270,
         div_DP_OP_279J39_124_314_n1269, div_DP_OP_279J39_124_314_n1268,
         div_DP_OP_279J39_124_314_n1267, div_DP_OP_279J39_124_314_n1266,
         div_DP_OP_279J39_124_314_n1265, div_DP_OP_279J39_124_314_n1264,
         div_DP_OP_279J39_124_314_n1263, div_DP_OP_279J39_124_314_n1262,
         div_DP_OP_279J39_124_314_n1261, div_DP_OP_279J39_124_314_n1260,
         div_DP_OP_279J39_124_314_n1259, div_DP_OP_279J39_124_314_n1258,
         div_DP_OP_279J39_124_314_n1257, div_DP_OP_279J39_124_314_n1256,
         div_DP_OP_279J39_124_314_n1255, div_DP_OP_279J39_124_314_n1254,
         div_DP_OP_279J39_124_314_n1253, div_DP_OP_279J39_124_314_n1252,
         div_DP_OP_279J39_124_314_n1251, div_DP_OP_279J39_124_314_n1250,
         div_DP_OP_279J39_124_314_n1249, div_DP_OP_279J39_124_314_n1248,
         div_DP_OP_279J39_124_314_n1247, div_DP_OP_279J39_124_314_n1246,
         div_DP_OP_279J39_124_314_n1245, div_DP_OP_279J39_124_314_n1244,
         div_DP_OP_279J39_124_314_n1243, div_DP_OP_279J39_124_314_n1242,
         div_DP_OP_279J39_124_314_n1241, div_DP_OP_279J39_124_314_n1240,
         div_DP_OP_279J39_124_314_n1239, div_DP_OP_279J39_124_314_n1238,
         div_DP_OP_279J39_124_314_n1237, div_DP_OP_279J39_124_314_n1236,
         div_DP_OP_279J39_124_314_n1235, div_DP_OP_279J39_124_314_n1234,
         div_DP_OP_279J39_124_314_n1233, div_DP_OP_279J39_124_314_n1232,
         div_DP_OP_279J39_124_314_n1231, div_DP_OP_279J39_124_314_n1230,
         div_DP_OP_279J39_124_314_n1229, div_DP_OP_279J39_124_314_n1228,
         div_DP_OP_279J39_124_314_n1227, div_DP_OP_279J39_124_314_n1226,
         div_DP_OP_279J39_124_314_n1225, div_DP_OP_279J39_124_314_n1224,
         div_DP_OP_279J39_124_314_n1223, div_DP_OP_279J39_124_314_n1222,
         div_DP_OP_279J39_124_314_n1221, div_DP_OP_279J39_124_314_n1220,
         div_DP_OP_279J39_124_314_n1219, div_DP_OP_279J39_124_314_n1218,
         div_DP_OP_279J39_124_314_n1217, div_DP_OP_279J39_124_314_n1216,
         div_DP_OP_279J39_124_314_n1215, div_DP_OP_279J39_124_314_n1214,
         div_DP_OP_279J39_124_314_n1213, div_DP_OP_279J39_124_314_n1212,
         div_DP_OP_279J39_124_314_n1211, div_DP_OP_279J39_124_314_n1210,
         div_DP_OP_279J39_124_314_n1209, div_DP_OP_279J39_124_314_n1208,
         div_DP_OP_279J39_124_314_n1207, div_DP_OP_279J39_124_314_n1206,
         div_DP_OP_279J39_124_314_n1205, div_DP_OP_279J39_124_314_n1204,
         div_DP_OP_279J39_124_314_n1203, div_DP_OP_279J39_124_314_n1202,
         div_DP_OP_279J39_124_314_n1201, div_DP_OP_279J39_124_314_n1200,
         div_DP_OP_279J39_124_314_n1199, div_DP_OP_279J39_124_314_n1198,
         div_DP_OP_279J39_124_314_n1197, div_DP_OP_279J39_124_314_n1196,
         div_DP_OP_279J39_124_314_n1195, div_DP_OP_279J39_124_314_n1194,
         div_DP_OP_279J39_124_314_n1193, div_DP_OP_279J39_124_314_n1192,
         div_DP_OP_279J39_124_314_n1191, div_DP_OP_279J39_124_314_n1190,
         div_DP_OP_279J39_124_314_n1189, div_DP_OP_279J39_124_314_n1188,
         div_DP_OP_279J39_124_314_n1187, div_DP_OP_279J39_124_314_n1186,
         div_DP_OP_279J39_124_314_n1185, div_DP_OP_279J39_124_314_n1184,
         div_DP_OP_279J39_124_314_n1183, div_DP_OP_279J39_124_314_n1182,
         div_DP_OP_279J39_124_314_n1181, div_DP_OP_279J39_124_314_n1180,
         div_DP_OP_279J39_124_314_n1179, div_DP_OP_279J39_124_314_n1178,
         div_DP_OP_279J39_124_314_n1177, div_DP_OP_279J39_124_314_n1176,
         div_DP_OP_279J39_124_314_n1175, div_DP_OP_279J39_124_314_n1174,
         div_DP_OP_279J39_124_314_n1173, div_DP_OP_279J39_124_314_n1172,
         div_DP_OP_279J39_124_314_n1171, div_DP_OP_279J39_124_314_n1170,
         div_DP_OP_279J39_124_314_n1169, div_DP_OP_279J39_124_314_n1168,
         div_DP_OP_279J39_124_314_n1167, div_DP_OP_279J39_124_314_n1166,
         div_DP_OP_279J39_124_314_n1165, div_DP_OP_279J39_124_314_n1164,
         div_DP_OP_279J39_124_314_n1163, div_DP_OP_279J39_124_314_n1162,
         div_DP_OP_279J39_124_314_n1161, div_DP_OP_279J39_124_314_n1160,
         div_DP_OP_279J39_124_314_n1159, div_DP_OP_279J39_124_314_n1158,
         div_DP_OP_279J39_124_314_n1157, div_DP_OP_279J39_124_314_n1156,
         div_DP_OP_279J39_124_314_n1155, div_DP_OP_279J39_124_314_n1154,
         div_DP_OP_279J39_124_314_n1153, div_DP_OP_279J39_124_314_n1152,
         div_DP_OP_279J39_124_314_n1151, div_DP_OP_279J39_124_314_n1150,
         div_DP_OP_279J39_124_314_n1149, div_DP_OP_279J39_124_314_n1148,
         div_DP_OP_279J39_124_314_n1147, div_DP_OP_279J39_124_314_n1146,
         div_DP_OP_279J39_124_314_n1145, div_DP_OP_279J39_124_314_n1144,
         div_DP_OP_279J39_124_314_n1143, div_DP_OP_279J39_124_314_n1142,
         div_DP_OP_279J39_124_314_n1141, div_DP_OP_279J39_124_314_n1140,
         div_DP_OP_279J39_124_314_n1139, div_DP_OP_279J39_124_314_n1138,
         div_DP_OP_279J39_124_314_n1137, div_DP_OP_279J39_124_314_n1136,
         div_DP_OP_279J39_124_314_n1135, div_DP_OP_279J39_124_314_n1134,
         div_DP_OP_279J39_124_314_n1133, div_DP_OP_279J39_124_314_n1132,
         div_DP_OP_279J39_124_314_n1131, div_DP_OP_279J39_124_314_n1130,
         div_DP_OP_279J39_124_314_n1129, div_DP_OP_279J39_124_314_n1128,
         div_DP_OP_279J39_124_314_n1127, div_DP_OP_279J39_124_314_n1126,
         div_DP_OP_279J39_124_314_n1125, div_DP_OP_279J39_124_314_n1124,
         div_DP_OP_279J39_124_314_n1123, div_DP_OP_279J39_124_314_n1122,
         div_DP_OP_279J39_124_314_n1121, div_DP_OP_279J39_124_314_n1120,
         div_DP_OP_279J39_124_314_n1119, div_DP_OP_279J39_124_314_n1118,
         div_DP_OP_279J39_124_314_n1117, div_DP_OP_279J39_124_314_n1116,
         div_DP_OP_279J39_124_314_n1115, div_DP_OP_279J39_124_314_n1114,
         div_DP_OP_279J39_124_314_n1113, div_DP_OP_279J39_124_314_n1112,
         div_DP_OP_279J39_124_314_n1111, div_DP_OP_279J39_124_314_n1110,
         div_DP_OP_279J39_124_314_n1109, div_DP_OP_279J39_124_314_n1108,
         div_DP_OP_279J39_124_314_n1107, div_DP_OP_279J39_124_314_n1106,
         div_DP_OP_279J39_124_314_n1105, div_DP_OP_279J39_124_314_n1104,
         div_DP_OP_279J39_124_314_n1103, div_DP_OP_279J39_124_314_n1102,
         div_DP_OP_279J39_124_314_n1101, div_DP_OP_279J39_124_314_n1100,
         div_DP_OP_279J39_124_314_n1099, div_DP_OP_279J39_124_314_n1098,
         div_DP_OP_279J39_124_314_n1097, div_DP_OP_279J39_124_314_n1096,
         div_DP_OP_279J39_124_314_n1095, div_DP_OP_279J39_124_314_n1094,
         div_DP_OP_279J39_124_314_n1093, div_DP_OP_279J39_124_314_n1092,
         div_DP_OP_279J39_124_314_n1091, div_DP_OP_279J39_124_314_n1090,
         div_DP_OP_279J39_124_314_n1089, div_DP_OP_279J39_124_314_n1088,
         div_DP_OP_279J39_124_314_n1087, div_DP_OP_279J39_124_314_n1086,
         div_DP_OP_279J39_124_314_n1085, div_DP_OP_279J39_124_314_n1084,
         div_DP_OP_279J39_124_314_n1083, div_DP_OP_279J39_124_314_n1082,
         div_DP_OP_279J39_124_314_n1081, div_DP_OP_279J39_124_314_n1080,
         div_DP_OP_279J39_124_314_n1079, div_DP_OP_279J39_124_314_n1078,
         div_DP_OP_279J39_124_314_n1077, div_DP_OP_279J39_124_314_n1076,
         div_DP_OP_279J39_124_314_n1075, div_DP_OP_279J39_124_314_n1074,
         div_DP_OP_279J39_124_314_n1073, div_DP_OP_279J39_124_314_n1072,
         div_DP_OP_279J39_124_314_n1071, div_DP_OP_279J39_124_314_n1070,
         div_DP_OP_279J39_124_314_n1069, div_DP_OP_279J39_124_314_n1068,
         div_DP_OP_279J39_124_314_n1067, div_DP_OP_279J39_124_314_n1066,
         div_DP_OP_279J39_124_314_n1065, div_DP_OP_279J39_124_314_n1064,
         div_DP_OP_279J39_124_314_n1063, div_DP_OP_279J39_124_314_n1062,
         div_DP_OP_279J39_124_314_n1061, div_DP_OP_279J39_124_314_n1060,
         div_DP_OP_279J39_124_314_n1059, div_DP_OP_279J39_124_314_n1058,
         div_DP_OP_279J39_124_314_n1057, div_DP_OP_279J39_124_314_n1056,
         div_DP_OP_279J39_124_314_n1055, div_DP_OP_279J39_124_314_n1054,
         div_DP_OP_279J39_124_314_n1053, div_DP_OP_279J39_124_314_n1052,
         div_DP_OP_279J39_124_314_n1051, div_DP_OP_279J39_124_314_n1050,
         div_DP_OP_279J39_124_314_n1049, div_DP_OP_279J39_124_314_n1048,
         div_DP_OP_279J39_124_314_n1047, div_DP_OP_279J39_124_314_n1046,
         div_DP_OP_279J39_124_314_n1045, div_DP_OP_279J39_124_314_n1044,
         div_DP_OP_279J39_124_314_n1043, div_DP_OP_279J39_124_314_n1042,
         div_DP_OP_279J39_124_314_n1041, div_DP_OP_279J39_124_314_n1040,
         div_DP_OP_279J39_124_314_n1039, div_DP_OP_279J39_124_314_n1038,
         div_DP_OP_279J39_124_314_n1037, div_DP_OP_279J39_124_314_n1036,
         div_DP_OP_279J39_124_314_n1035, div_DP_OP_279J39_124_314_n1034,
         div_DP_OP_279J39_124_314_n1033, div_DP_OP_279J39_124_314_n1032,
         div_DP_OP_279J39_124_314_n1031, div_DP_OP_279J39_124_314_n1030,
         div_DP_OP_279J39_124_314_n1029, div_DP_OP_279J39_124_314_n1028,
         div_DP_OP_279J39_124_314_n1027, div_DP_OP_279J39_124_314_n1026,
         div_DP_OP_279J39_124_314_n1025, div_DP_OP_279J39_124_314_n1024,
         div_DP_OP_279J39_124_314_n1023, div_DP_OP_279J39_124_314_n1022,
         div_DP_OP_279J39_124_314_n1021, div_DP_OP_279J39_124_314_n1020,
         div_DP_OP_279J39_124_314_n1019, div_DP_OP_279J39_124_314_n1018,
         div_DP_OP_279J39_124_314_n1017, div_DP_OP_279J39_124_314_n1016,
         div_DP_OP_279J39_124_314_n1015, div_DP_OP_279J39_124_314_n1014,
         div_DP_OP_279J39_124_314_n1013, div_DP_OP_279J39_124_314_n1012,
         div_DP_OP_279J39_124_314_n1011, div_DP_OP_279J39_124_314_n1010,
         div_DP_OP_279J39_124_314_n1009, div_DP_OP_279J39_124_314_n1008,
         div_DP_OP_279J39_124_314_n1007, div_DP_OP_279J39_124_314_n1006,
         div_DP_OP_279J39_124_314_n1005, div_DP_OP_279J39_124_314_n1004,
         div_DP_OP_279J39_124_314_n1003, div_DP_OP_279J39_124_314_n1002,
         div_DP_OP_279J39_124_314_n1001, div_DP_OP_279J39_124_314_n1000,
         div_DP_OP_279J39_124_314_n999, div_DP_OP_279J39_124_314_n998,
         div_DP_OP_279J39_124_314_n997, div_DP_OP_279J39_124_314_n996,
         div_DP_OP_279J39_124_314_n995, div_DP_OP_279J39_124_314_n994,
         div_DP_OP_279J39_124_314_n993, div_DP_OP_279J39_124_314_n992,
         div_DP_OP_279J39_124_314_n991, div_DP_OP_279J39_124_314_n990,
         div_DP_OP_279J39_124_314_n989, div_DP_OP_279J39_124_314_n988,
         div_DP_OP_279J39_124_314_n987, div_DP_OP_279J39_124_314_n986,
         div_DP_OP_279J39_124_314_n985, div_DP_OP_279J39_124_314_n984,
         div_DP_OP_279J39_124_314_n983, div_DP_OP_279J39_124_314_n982,
         div_DP_OP_279J39_124_314_n981, div_DP_OP_279J39_124_314_n980,
         div_DP_OP_279J39_124_314_n979, div_DP_OP_279J39_124_314_n978,
         div_DP_OP_279J39_124_314_n977, div_DP_OP_279J39_124_314_n976,
         div_DP_OP_279J39_124_314_n975, div_DP_OP_279J39_124_314_n974,
         div_DP_OP_279J39_124_314_n973, div_DP_OP_279J39_124_314_n972,
         div_DP_OP_279J39_124_314_n971, div_DP_OP_279J39_124_314_n970,
         div_DP_OP_279J39_124_314_n969, div_DP_OP_279J39_124_314_n968,
         div_DP_OP_279J39_124_314_n967, div_DP_OP_279J39_124_314_n966,
         div_DP_OP_279J39_124_314_n965, div_DP_OP_279J39_124_314_n964,
         div_DP_OP_279J39_124_314_n963, div_DP_OP_279J39_124_314_n962,
         div_DP_OP_279J39_124_314_n961, div_DP_OP_279J39_124_314_n960,
         div_DP_OP_279J39_124_314_n959, div_DP_OP_279J39_124_314_n958,
         div_DP_OP_279J39_124_314_n957, div_DP_OP_279J39_124_314_n956,
         div_DP_OP_279J39_124_314_n955, div_DP_OP_279J39_124_314_n954,
         div_DP_OP_279J39_124_314_n953, div_DP_OP_279J39_124_314_n952,
         div_DP_OP_279J39_124_314_n951, div_DP_OP_279J39_124_314_n950,
         div_DP_OP_279J39_124_314_n949, div_DP_OP_279J39_124_314_n948,
         div_DP_OP_279J39_124_314_n947, div_DP_OP_279J39_124_314_n946,
         div_DP_OP_279J39_124_314_n945, div_DP_OP_279J39_124_314_n944,
         div_DP_OP_279J39_124_314_n943, div_DP_OP_279J39_124_314_n942,
         div_DP_OP_279J39_124_314_n941, div_DP_OP_279J39_124_314_n940,
         div_DP_OP_279J39_124_314_n939, div_DP_OP_279J39_124_314_n938,
         div_DP_OP_279J39_124_314_n937, div_DP_OP_279J39_124_314_n936,
         div_DP_OP_279J39_124_314_n935, div_DP_OP_279J39_124_314_n934,
         div_DP_OP_279J39_124_314_n933, div_DP_OP_279J39_124_314_n932,
         div_DP_OP_279J39_124_314_n931, div_DP_OP_279J39_124_314_n930,
         div_DP_OP_279J39_124_314_n929, div_DP_OP_279J39_124_314_n928,
         div_DP_OP_279J39_124_314_n927, div_DP_OP_279J39_124_314_n926,
         div_DP_OP_279J39_124_314_n925, div_DP_OP_279J39_124_314_n924,
         div_DP_OP_279J39_124_314_n923, div_DP_OP_279J39_124_314_n922,
         div_DP_OP_279J39_124_314_n921, div_DP_OP_279J39_124_314_n920,
         div_DP_OP_279J39_124_314_n919, div_DP_OP_279J39_124_314_n918,
         div_DP_OP_279J39_124_314_n917, div_DP_OP_279J39_124_314_n916,
         div_DP_OP_279J39_124_314_n915, div_DP_OP_279J39_124_314_n914,
         div_DP_OP_279J39_124_314_n913, div_DP_OP_279J39_124_314_n912,
         div_DP_OP_279J39_124_314_n911, div_DP_OP_279J39_124_314_n910,
         div_DP_OP_279J39_124_314_n909, div_DP_OP_279J39_124_314_n908,
         div_DP_OP_279J39_124_314_n907, div_DP_OP_279J39_124_314_n906,
         div_DP_OP_279J39_124_314_n905, div_DP_OP_279J39_124_314_n904,
         div_DP_OP_279J39_124_314_n903, div_DP_OP_279J39_124_314_n902,
         div_DP_OP_279J39_124_314_n901, div_DP_OP_279J39_124_314_n900,
         div_DP_OP_279J39_124_314_n899, div_DP_OP_279J39_124_314_n898,
         div_DP_OP_279J39_124_314_n897, div_DP_OP_279J39_124_314_n896,
         div_DP_OP_279J39_124_314_n895, div_DP_OP_279J39_124_314_n894,
         div_DP_OP_279J39_124_314_n893, div_DP_OP_279J39_124_314_n892,
         div_DP_OP_279J39_124_314_n891, div_DP_OP_279J39_124_314_n890,
         div_DP_OP_279J39_124_314_n889, div_DP_OP_279J39_124_314_n888,
         div_DP_OP_279J39_124_314_n887, div_DP_OP_279J39_124_314_n886,
         div_DP_OP_279J39_124_314_n885, div_DP_OP_279J39_124_314_n884,
         div_DP_OP_279J39_124_314_n883, div_DP_OP_279J39_124_314_n882,
         div_DP_OP_279J39_124_314_n881, div_DP_OP_279J39_124_314_n880,
         div_DP_OP_279J39_124_314_n879, div_DP_OP_279J39_124_314_n878,
         div_DP_OP_279J39_124_314_n877, div_DP_OP_279J39_124_314_n876,
         div_DP_OP_279J39_124_314_n875, div_DP_OP_279J39_124_314_n874,
         div_DP_OP_279J39_124_314_n873, div_DP_OP_279J39_124_314_n872,
         div_DP_OP_279J39_124_314_n871, div_DP_OP_279J39_124_314_n870,
         div_DP_OP_279J39_124_314_n869, div_DP_OP_279J39_124_314_n868,
         div_DP_OP_279J39_124_314_n867, div_DP_OP_279J39_124_314_n866,
         div_DP_OP_279J39_124_314_n865, div_DP_OP_279J39_124_314_n864,
         div_DP_OP_279J39_124_314_n863, div_DP_OP_279J39_124_314_n862,
         div_DP_OP_279J39_124_314_n861, div_DP_OP_279J39_124_314_n860,
         div_DP_OP_279J39_124_314_n859, div_DP_OP_279J39_124_314_n858,
         div_DP_OP_279J39_124_314_n857, div_DP_OP_279J39_124_314_n856,
         div_DP_OP_279J39_124_314_n855, div_DP_OP_279J39_124_314_n854,
         div_DP_OP_279J39_124_314_n853, div_DP_OP_279J39_124_314_n852,
         div_DP_OP_279J39_124_314_n851, div_DP_OP_279J39_124_314_n850,
         div_DP_OP_279J39_124_314_n849, div_DP_OP_279J39_124_314_n848,
         div_DP_OP_279J39_124_314_n847, div_DP_OP_279J39_124_314_n846,
         div_DP_OP_279J39_124_314_n845, div_DP_OP_279J39_124_314_n844,
         div_DP_OP_279J39_124_314_n843, div_DP_OP_279J39_124_314_n842,
         div_DP_OP_279J39_124_314_n841, div_DP_OP_279J39_124_314_n840,
         div_DP_OP_279J39_124_314_n839, div_DP_OP_279J39_124_314_n838,
         div_DP_OP_279J39_124_314_n837, div_DP_OP_279J39_124_314_n836,
         div_DP_OP_279J39_124_314_n835, div_DP_OP_279J39_124_314_n834,
         div_DP_OP_279J39_124_314_n833, div_DP_OP_279J39_124_314_n832,
         div_DP_OP_279J39_124_314_n831, div_DP_OP_279J39_124_314_n830,
         div_DP_OP_279J39_124_314_n829, div_DP_OP_279J39_124_314_n828,
         div_DP_OP_279J39_124_314_n827, div_DP_OP_279J39_124_314_n826,
         div_DP_OP_279J39_124_314_n825, div_DP_OP_279J39_124_314_n824,
         div_DP_OP_279J39_124_314_n823, div_DP_OP_279J39_124_314_n822,
         div_DP_OP_279J39_124_314_n821, div_DP_OP_279J39_124_314_n820,
         div_DP_OP_279J39_124_314_n819, div_DP_OP_279J39_124_314_n818,
         div_DP_OP_279J39_124_314_n817, div_DP_OP_279J39_124_314_n816,
         div_DP_OP_279J39_124_314_n815, div_DP_OP_279J39_124_314_n814,
         div_DP_OP_279J39_124_314_n813, div_DP_OP_279J39_124_314_n812,
         div_DP_OP_279J39_124_314_n811, div_DP_OP_279J39_124_314_n810,
         div_DP_OP_279J39_124_314_n809, div_DP_OP_279J39_124_314_n808,
         div_DP_OP_279J39_124_314_n807, div_DP_OP_279J39_124_314_n806,
         div_DP_OP_279J39_124_314_n805, div_DP_OP_279J39_124_314_n804,
         div_DP_OP_279J39_124_314_n803, div_DP_OP_279J39_124_314_n802,
         div_DP_OP_279J39_124_314_n801, div_DP_OP_279J39_124_314_n800,
         div_DP_OP_279J39_124_314_n799, div_DP_OP_279J39_124_314_n798,
         div_DP_OP_279J39_124_314_n797, div_DP_OP_279J39_124_314_n796,
         div_DP_OP_279J39_124_314_n795, div_DP_OP_279J39_124_314_n794,
         div_DP_OP_279J39_124_314_n793, div_DP_OP_279J39_124_314_n792,
         div_DP_OP_279J39_124_314_n791, div_DP_OP_279J39_124_314_n790,
         div_DP_OP_279J39_124_314_n789, div_DP_OP_279J39_124_314_n788,
         div_DP_OP_279J39_124_314_n787, div_DP_OP_279J39_124_314_n786,
         div_DP_OP_279J39_124_314_n785, div_DP_OP_279J39_124_314_n784,
         div_DP_OP_279J39_124_314_n783, div_DP_OP_279J39_124_314_n782,
         div_DP_OP_279J39_124_314_n781, div_DP_OP_279J39_124_314_n780,
         div_DP_OP_279J39_124_314_n779, div_DP_OP_279J39_124_314_n778,
         div_DP_OP_279J39_124_314_n777, div_DP_OP_279J39_124_314_n776,
         div_DP_OP_279J39_124_314_n775, div_DP_OP_279J39_124_314_n774,
         div_DP_OP_279J39_124_314_n773, div_DP_OP_279J39_124_314_n772,
         div_DP_OP_279J39_124_314_n771, div_DP_OP_279J39_124_314_n770,
         div_DP_OP_279J39_124_314_n769, div_DP_OP_279J39_124_314_n768,
         div_DP_OP_279J39_124_314_n767, div_DP_OP_279J39_124_314_n766,
         div_DP_OP_279J39_124_314_n765, div_DP_OP_279J39_124_314_n764,
         div_DP_OP_279J39_124_314_n763, div_DP_OP_279J39_124_314_n762,
         div_DP_OP_279J39_124_314_n761, div_DP_OP_279J39_124_314_n760,
         div_DP_OP_279J39_124_314_n759, div_DP_OP_279J39_124_314_n758,
         div_DP_OP_279J39_124_314_n757, div_DP_OP_279J39_124_314_n756,
         div_DP_OP_279J39_124_314_n755, div_DP_OP_279J39_124_314_n754,
         div_DP_OP_279J39_124_314_n753, div_DP_OP_279J39_124_314_n752,
         div_DP_OP_279J39_124_314_n751, div_DP_OP_279J39_124_314_n750,
         div_DP_OP_279J39_124_314_n749, div_DP_OP_279J39_124_314_n748,
         div_DP_OP_279J39_124_314_n747, div_DP_OP_279J39_124_314_n746,
         div_DP_OP_279J39_124_314_n745, div_DP_OP_279J39_124_314_n744,
         div_DP_OP_279J39_124_314_n743, div_DP_OP_279J39_124_314_n742,
         div_DP_OP_279J39_124_314_n741, div_DP_OP_279J39_124_314_n740,
         div_DP_OP_279J39_124_314_n739, div_DP_OP_279J39_124_314_n738,
         div_DP_OP_279J39_124_314_n737, div_DP_OP_279J39_124_314_n736,
         div_DP_OP_279J39_124_314_n735, div_DP_OP_279J39_124_314_n734,
         div_DP_OP_279J39_124_314_n733, div_DP_OP_279J39_124_314_n732,
         div_DP_OP_279J39_124_314_n731, div_DP_OP_279J39_124_314_n730,
         div_DP_OP_279J39_124_314_n729, div_DP_OP_279J39_124_314_n728,
         div_DP_OP_279J39_124_314_n727, div_DP_OP_279J39_124_314_n726,
         div_DP_OP_279J39_124_314_n725, div_DP_OP_279J39_124_314_n724,
         div_DP_OP_279J39_124_314_n723, div_DP_OP_279J39_124_314_n722,
         div_DP_OP_279J39_124_314_n721, div_DP_OP_279J39_124_314_n720,
         div_DP_OP_279J39_124_314_n719, div_DP_OP_279J39_124_314_n718,
         div_DP_OP_279J39_124_314_n717, div_DP_OP_279J39_124_314_n716,
         div_DP_OP_279J39_124_314_n715, div_DP_OP_279J39_124_314_n714,
         div_DP_OP_279J39_124_314_n713, div_DP_OP_279J39_124_314_n712,
         div_DP_OP_279J39_124_314_n711, div_DP_OP_279J39_124_314_n710,
         div_DP_OP_279J39_124_314_n709, div_DP_OP_279J39_124_314_n708,
         div_DP_OP_279J39_124_314_n707, div_DP_OP_279J39_124_314_n706,
         div_DP_OP_279J39_124_314_n705, div_DP_OP_279J39_124_314_n704,
         div_DP_OP_279J39_124_314_n703, div_DP_OP_279J39_124_314_n702,
         div_DP_OP_279J39_124_314_n701, div_DP_OP_279J39_124_314_n700,
         div_DP_OP_279J39_124_314_n699, div_DP_OP_279J39_124_314_n698,
         div_DP_OP_279J39_124_314_n697, div_DP_OP_279J39_124_314_n696,
         div_DP_OP_279J39_124_314_n695, div_DP_OP_279J39_124_314_n694,
         div_DP_OP_279J39_124_314_n693, div_DP_OP_279J39_124_314_n692,
         div_DP_OP_279J39_124_314_n691, div_DP_OP_279J39_124_314_n690,
         div_DP_OP_279J39_124_314_n689, div_DP_OP_279J39_124_314_n688,
         div_DP_OP_279J39_124_314_n687, div_DP_OP_279J39_124_314_n686,
         div_DP_OP_279J39_124_314_n685, div_DP_OP_279J39_124_314_n684,
         div_DP_OP_279J39_124_314_n683, div_DP_OP_279J39_124_314_n682,
         div_DP_OP_279J39_124_314_n681, div_DP_OP_279J39_124_314_n680,
         div_DP_OP_279J39_124_314_n679, div_DP_OP_279J39_124_314_n678,
         div_DP_OP_279J39_124_314_n677, div_DP_OP_279J39_124_314_n676,
         div_DP_OP_279J39_124_314_n675, div_DP_OP_279J39_124_314_n674,
         div_DP_OP_279J39_124_314_n673, div_DP_OP_279J39_124_314_n672,
         div_DP_OP_279J39_124_314_n671, div_DP_OP_279J39_124_314_n670,
         div_DP_OP_279J39_124_314_n669, div_DP_OP_279J39_124_314_n668,
         div_DP_OP_279J39_124_314_n667, div_DP_OP_279J39_124_314_n666,
         div_DP_OP_279J39_124_314_n665, div_DP_OP_279J39_124_314_n664,
         div_DP_OP_279J39_124_314_n663, div_DP_OP_279J39_124_314_n662,
         div_DP_OP_279J39_124_314_n661, div_DP_OP_279J39_124_314_n660,
         div_DP_OP_279J39_124_314_n659, div_DP_OP_279J39_124_314_n658,
         div_DP_OP_279J39_124_314_n657, div_DP_OP_279J39_124_314_n656,
         div_DP_OP_279J39_124_314_n655, div_DP_OP_279J39_124_314_n654,
         div_DP_OP_279J39_124_314_n653, div_DP_OP_279J39_124_314_n652,
         div_DP_OP_279J39_124_314_n651, div_DP_OP_279J39_124_314_n650,
         div_DP_OP_279J39_124_314_n649, div_DP_OP_279J39_124_314_n648,
         div_DP_OP_279J39_124_314_n647, div_DP_OP_279J39_124_314_n646,
         div_DP_OP_279J39_124_314_n645, div_DP_OP_279J39_124_314_n644,
         div_DP_OP_279J39_124_314_n643, div_DP_OP_279J39_124_314_n642,
         div_DP_OP_279J39_124_314_n641, div_DP_OP_279J39_124_314_n640,
         div_DP_OP_279J39_124_314_n639, div_DP_OP_279J39_124_314_n638,
         div_DP_OP_279J39_124_314_n637, div_DP_OP_279J39_124_314_n636,
         div_DP_OP_279J39_124_314_n635, div_DP_OP_279J39_124_314_n634,
         div_DP_OP_279J39_124_314_n633, div_DP_OP_279J39_124_314_n632,
         div_DP_OP_279J39_124_314_n631, div_DP_OP_279J39_124_314_n630,
         div_DP_OP_279J39_124_314_n629, div_DP_OP_279J39_124_314_n628,
         div_DP_OP_279J39_124_314_n627, div_DP_OP_279J39_124_314_n551,
         div_ash_111_n1038, div_ash_111_n1037, div_ash_111_n1036,
         div_ash_111_n1035, div_ash_111_n1034, div_ash_111_n1033,
         div_ash_111_n1032, div_ash_111_n1031, div_ash_111_n1030,
         div_ash_111_n1029, div_ash_111_n1028, div_ash_111_n1027,
         div_ash_111_n1026, div_ash_111_n1025, div_ash_111_n1024,
         div_ash_111_n1023, div_ash_111_n1022, div_ash_111_n1021,
         div_ash_111_n1020, div_ash_111_n1019, div_ash_111_n1018,
         div_ash_111_n1017, div_ash_111_n1016, div_ash_111_n1015,
         div_ash_111_n1014, div_ash_111_n1013, div_ash_111_n1012,
         div_ash_111_n1011, div_ash_111_n1010, div_ash_111_n1009,
         div_ash_111_n1008, div_ash_111_n1007, div_ash_111_n1006,
         div_ash_111_n1005, div_ash_111_n1004, div_ash_111_n1003,
         div_ash_111_n1002, div_ash_111_n1001, div_ash_111_n1000,
         div_ash_111_n999, div_ash_111_n998, div_ash_111_n997,
         div_ash_111_n996, div_ash_111_n995, div_ash_111_n994,
         div_ash_111_n993, div_ash_111_n992, div_ash_111_n991,
         div_ash_111_n990, div_ash_111_n989, div_ash_111_n988,
         div_ash_111_n987, div_ash_111_n986, div_ash_111_n985,
         div_ash_111_n984, div_ash_111_n983, div_ash_111_n982,
         div_ash_111_n981, div_ash_111_n980, div_ash_111_n979,
         div_ash_111_n978, div_ash_111_n977, div_ash_111_n976,
         div_ash_111_n975, div_ash_111_n974, div_ash_111_n973,
         div_ash_111_n972, div_ash_111_n971, div_ash_111_n970,
         div_ash_111_n969, div_ash_111_n968, div_ash_111_n967,
         div_ash_111_n966, div_ash_111_n965, div_ash_111_n964,
         div_ash_111_n963, div_ash_111_n962, div_ash_111_n961,
         div_ash_111_n960, div_ash_111_n959, div_ash_111_n958,
         div_ash_111_n957, div_ash_111_n956, div_ash_111_n955,
         div_ash_111_n954, div_ash_111_n953, div_ash_111_n952,
         div_ash_111_n951, div_ash_111_n950, div_ash_111_n949,
         div_ash_111_n948, div_ash_111_n947, div_ash_111_n946,
         div_ash_111_n945, div_ash_111_n944, div_ash_111_n943,
         div_ash_111_n942, div_ash_111_n941, div_ash_111_n940,
         div_ash_111_n939, div_ash_111_n938, div_ash_111_n937,
         div_ash_111_n936, div_ash_111_n935, div_ash_111_n934,
         div_ash_111_n933, div_ash_111_n932, div_ash_111_n931,
         div_ash_111_n930, div_ash_111_n929, div_ash_111_n928,
         div_ash_111_n927, div_ash_111_n926, div_ash_111_n925,
         div_ash_111_n924, div_ash_111_n923, div_ash_111_n922,
         div_ash_111_n921, div_ash_111_n920, div_ash_111_n919,
         div_ash_111_n918, div_ash_111_n917, div_ash_111_n916,
         div_ash_111_n915, div_ash_111_n914, div_ash_111_n913,
         div_ash_111_n912, div_ash_111_n911, div_ash_111_n910,
         div_ash_111_n909, div_ash_111_n908, div_ash_111_n907,
         div_ash_111_n906, div_ash_111_n905, div_ash_111_n904,
         div_ash_111_n903, div_ash_111_n902, div_ash_111_n901,
         div_ash_111_n900, div_ash_111_n899, div_ash_111_n898,
         div_ash_111_n897, div_ash_111_n896, div_ash_111_n895,
         div_ash_111_n894, div_ash_111_n893, div_ash_111_n892,
         div_ash_111_n891, div_ash_111_n890, div_ash_111_n889,
         div_ash_111_n888, div_ash_111_n887, div_ash_111_n886,
         div_ash_111_n885, div_ash_111_n884, div_ash_111_n883,
         div_ash_111_n882, div_ash_111_n881, div_ash_111_n880,
         div_ash_111_n879, div_ash_111_n878, div_ash_111_n877,
         div_ash_111_n876, div_ash_111_n875, div_ash_111_n874,
         div_ash_111_n873, div_ash_111_n872, div_ash_111_n871,
         div_ash_111_n870, div_ash_111_n869, div_ash_111_n868,
         div_ash_111_n867, div_ash_111_n866, div_ash_111_n865,
         div_ash_111_n864, div_ash_111_n863, div_ash_111_n862,
         div_ash_111_n861, div_ash_111_n860, div_ash_111_n859,
         div_ash_111_n858, div_ash_111_n857, div_ash_111_n856,
         div_ash_111_n855, div_ash_111_n854, div_ash_111_n853,
         div_ash_111_n852, div_ash_111_n851, div_ash_111_n850,
         div_ash_111_n849, div_ash_111_n848, div_ash_111_n847,
         div_ash_111_n846, div_ash_111_n845, div_ash_111_n844,
         div_ash_111_n843, div_ash_111_n842, div_ash_111_n841,
         div_ash_111_n840, div_ash_111_n839, div_ash_111_n838,
         div_ash_111_n837, div_ash_111_n836, div_ash_111_n835,
         div_ash_111_n834, div_ash_111_n833, div_ash_111_n832,
         div_ash_111_n831, div_ash_111_n830, div_ash_111_n829,
         div_ash_111_n828, div_ash_111_n827, div_ash_111_n826,
         div_ash_111_n825, div_ash_111_n824, div_ash_111_n823,
         div_ash_111_n822, div_ash_111_n821, div_ash_111_n820,
         div_ash_111_n819, div_ash_111_n818, div_ash_111_n817,
         div_ash_111_n816, div_ash_111_n815, div_ash_111_n814,
         div_ash_111_n813, div_ash_111_n812, div_ash_111_n811,
         div_ash_111_n810, div_ash_111_n809, div_ash_111_n808,
         div_ash_111_n807, div_ash_111_n806, div_ash_111_n805,
         div_ash_111_n804, div_ash_111_n803, div_ash_111_n802,
         div_ash_111_n801, div_ash_111_n800, div_ash_111_n799,
         div_ash_111_n798, div_ash_111_n797, div_ash_111_n796,
         div_ash_111_n795, div_ash_111_n794, div_ash_111_n793,
         div_ash_111_n792, div_ash_111_n791, div_ash_111_n790,
         div_ash_111_n789, div_ash_111_n788, div_ash_111_n787,
         div_ash_111_n786, div_ash_111_n785, div_ash_111_n784,
         div_ash_111_n783, div_ash_111_n782, div_ash_111_n781,
         div_ash_111_n780, div_ash_111_n779, div_ash_111_n778,
         div_ash_111_n777, div_ash_111_n776, div_ash_111_n775,
         div_ash_111_n774, div_ash_111_n773, div_ash_111_n772,
         div_ash_111_n771, div_ash_111_n770, div_ash_111_n769,
         div_ash_111_n768, div_ash_111_n767, div_ash_111_n766,
         div_ash_111_n765, div_ash_111_n764, div_ash_111_n763,
         div_ash_111_n762, div_ash_111_n761, div_ash_111_n760,
         div_ash_111_n759, div_ash_111_n758, div_ash_111_n757,
         div_ash_111_n756, div_ash_111_n755, div_ash_111_n754,
         div_ash_111_n753, div_ash_111_n752, div_ash_111_n751,
         div_ash_111_n750, div_ash_111_n749, div_ash_111_n748,
         div_ash_111_n747, div_ash_111_n746, div_ash_111_n745,
         div_ash_111_n744, div_ash_111_n743, div_ash_111_n742,
         div_ash_111_n741, div_ash_111_n740, div_ash_111_n739,
         div_ash_111_n738, div_ash_111_n737, div_ash_111_n736,
         div_ash_111_n735, div_ash_111_n734, div_ash_111_n733,
         div_ash_111_n732, div_ash_111_n731, div_ash_111_n730,
         div_ash_111_n729, div_ash_111_n728, div_ash_111_n727,
         div_ash_111_n726, div_ash_111_n725, div_ash_111_n724,
         div_ash_111_n723, div_ash_111_n722, div_ash_111_n721,
         div_ash_111_n720, div_ash_111_n719, div_ash_111_n718,
         div_ash_111_n717, div_ash_111_n716, div_ash_111_n715,
         div_ash_111_n714, div_ash_111_n713, div_ash_111_n712,
         div_ash_111_n711, div_ash_111_n710, div_ash_111_n709,
         div_ash_111_n708, div_ash_111_n707, div_ash_111_n706,
         div_ash_111_n705, div_ash_111_n704, div_ash_111_n703,
         div_ash_111_n702, div_ash_111_n701, div_ash_111_n700,
         div_ash_111_n699, div_ash_111_n698, div_ash_111_n697,
         div_ash_111_n696, div_ash_111_n695, div_ash_111_n694,
         div_ash_111_n693, div_ash_111_n692, div_ash_111_n691,
         div_ash_111_n690, div_ash_111_n689, div_ash_111_n688,
         div_ash_111_n687, div_ash_111_n686, div_ash_111_n685,
         div_ash_111_n684, div_ash_111_n683, div_ash_111_n682,
         div_ash_111_n681, div_ash_111_n680, div_ash_111_n679,
         div_sub_x_110_n85, div_sub_x_110_n84, div_sub_x_110_n83,
         div_sub_x_110_n82, div_sub_x_110_n81, div_sub_x_110_n80,
         div_sub_x_110_n79, div_sub_x_110_n78, div_sub_x_110_n77,
         div_sub_x_110_n76, div_sub_x_110_n75, div_sub_x_110_n74,
         div_sub_x_110_n73, div_sub_x_110_n72, div_sub_x_110_n71,
         div_sub_x_110_n70, div_sub_x_110_n69, div_sub_x_110_n68,
         div_sub_x_110_n67, div_sub_x_110_n66, div_sub_x_110_n65,
         div_sub_x_110_n64, div_ashr_12_n1043, div_ashr_12_n1042,
         div_ashr_12_n1041, div_ashr_12_n1040, div_ashr_12_n1039,
         div_ashr_12_n1038, div_ashr_12_n1037, div_ashr_12_n1036,
         div_ashr_12_n1035, div_ashr_12_n1034, div_ashr_12_n1033,
         div_ashr_12_n1032, div_ashr_12_n1031, div_ashr_12_n1030,
         div_ashr_12_n1029, div_ashr_12_n1028, div_ashr_12_n1027,
         div_ashr_12_n1026, div_ashr_12_n1025, div_ashr_12_n1024,
         div_ashr_12_n1023, div_ashr_12_n1022, div_ashr_12_n1021,
         div_ashr_12_n1020, div_ashr_12_n1019, div_ashr_12_n1018,
         div_ashr_12_n1017, div_ashr_12_n1016, div_ashr_12_n1015,
         div_ashr_12_n1014, div_ashr_12_n1013, div_ashr_12_n1012,
         div_ashr_12_n1011, div_ashr_12_n1010, div_ashr_12_n1009,
         div_ashr_12_n1008, div_ashr_12_n1007, div_ashr_12_n1006,
         div_ashr_12_n1005, div_ashr_12_n1004, div_ashr_12_n1003,
         div_ashr_12_n1002, div_ashr_12_n1001, div_ashr_12_n1000,
         div_ashr_12_n999, div_ashr_12_n998, div_ashr_12_n997,
         div_ashr_12_n996, div_ashr_12_n995, div_ashr_12_n994,
         div_ashr_12_n993, div_ashr_12_n992, div_ashr_12_n991,
         div_ashr_12_n990, div_ashr_12_n989, div_ashr_12_n988,
         div_ashr_12_n987, div_ashr_12_n986, div_ashr_12_n985,
         div_ashr_12_n984, div_ashr_12_n983, div_ashr_12_n982,
         div_ashr_12_n981, div_ashr_12_n980, div_ashr_12_n979,
         div_ashr_12_n978, div_ashr_12_n977, div_ashr_12_n976,
         div_ashr_12_n975, div_ashr_12_n974, div_ashr_12_n973,
         div_ashr_12_n972, div_ashr_12_n971, div_ashr_12_n970,
         div_ashr_12_n969, div_ashr_12_n968, div_ashr_12_n967,
         div_ashr_12_n966, div_ashr_12_n965, div_ashr_12_n964,
         div_ashr_12_n963, div_ashr_12_n962, div_ashr_12_n961,
         div_ashr_12_n960, div_ashr_12_n959, div_ashr_12_n958,
         div_ashr_12_n957, div_ashr_12_n956, div_ashr_12_n955,
         div_ashr_12_n954, div_ashr_12_n953, div_ashr_12_n952,
         div_ashr_12_n951, div_ashr_12_n950, div_ashr_12_n949,
         div_ashr_12_n948, div_ashr_12_n947, div_ashr_12_n946,
         div_ashr_12_n945, div_ashr_12_n944, div_ashr_12_n943,
         div_ashr_12_n942, div_ashr_12_n941, div_ashr_12_n940,
         div_ashr_12_n939, div_ashr_12_n938, div_ashr_12_n937,
         div_ashr_12_n936, div_ashr_12_n935, div_ashr_12_n934,
         div_ashr_12_n933, div_ashr_12_n932, div_ashr_12_n931,
         div_ashr_12_n930, div_ashr_12_n929, div_ashr_12_n928,
         div_ashr_12_n927, div_ashr_12_n926, div_ashr_12_n925,
         div_ashr_12_n924, div_ashr_12_n923, div_ashr_12_n922,
         div_ashr_12_n921, div_ashr_12_n920, div_ashr_12_n919,
         div_ashr_12_n918, div_ashr_12_n917, div_ashr_12_n916,
         div_ashr_12_n915, div_ashr_12_n914, div_ashr_12_n913,
         div_ashr_12_n912, div_ashr_12_n911, div_ashr_12_n910,
         div_ashr_12_n909, div_ashr_12_n908, div_ashr_12_n907,
         div_ashr_12_n906, div_ashr_12_n905, div_ashr_12_n904,
         div_ashr_12_n903, div_ashr_12_n902, div_ashr_12_n901,
         div_ashr_12_n900, div_ashr_12_n899, div_ashr_12_n898,
         div_ashr_12_n897, div_ashr_12_n896, div_ashr_12_n895,
         div_ashr_12_n894, div_ashr_12_n893, div_ashr_12_n892,
         div_ashr_12_n891, div_ashr_12_n890, div_ashr_12_n889,
         div_ashr_12_n888, div_ashr_12_n887, div_ashr_12_n886,
         div_ashr_12_n885, div_ashr_12_n884, div_ashr_12_n883,
         div_ashr_12_n882, div_ashr_12_n881, div_ashr_12_n880,
         div_ashr_12_n879, div_ashr_12_n878, div_ashr_12_n877,
         div_ashr_12_n876, div_ashr_12_n875, div_ashr_12_n874,
         div_ashr_12_n873, div_ashr_12_n872, div_ashr_12_n871,
         div_ashr_12_n870, div_ashr_12_n869, div_ashr_12_n868,
         div_ashr_12_n867, div_ashr_12_n866, div_ashr_12_n865,
         div_ashr_12_n864, div_ashr_12_n863, div_ashr_12_n862,
         div_ashr_12_n861, div_ashr_12_n860, div_ashr_12_n859,
         div_ashr_12_n858, div_ashr_12_n857, div_ashr_12_n856,
         div_ashr_12_n855, div_ashr_12_n854, div_ashr_12_n853,
         div_ashr_12_n852, div_ashr_12_n851, div_ashr_12_n850,
         div_ashr_12_n849, div_ashr_12_n848, div_ashr_12_n847,
         div_ashr_12_n846, div_ashr_12_n845, div_ashr_12_n844,
         div_ashr_12_n843, div_ashr_12_n842, div_ashr_12_n841,
         div_ashr_12_n840, div_ashr_12_n839, div_ashr_12_n838,
         div_ashr_12_n837, div_ashr_12_n836, div_ashr_12_n835,
         div_ashr_12_n834, div_ashr_12_n833, div_ashr_12_n832,
         div_sub_x_9_n465, div_sub_x_9_n464, div_sub_x_9_n463,
         div_sub_x_9_n462, div_sub_x_9_n461, div_sub_x_9_n460,
         div_sub_x_9_n459, div_sub_x_9_n458, div_sub_x_9_n457,
         div_sub_x_9_n456, div_sub_x_9_n455, div_sub_x_9_n454,
         div_sub_x_9_n453, div_sub_x_9_n452, div_sub_x_9_n451,
         div_sub_x_9_n450, div_sub_x_9_n449, div_sub_x_9_n448,
         div_sub_x_9_n447, div_sub_x_9_n446, div_sub_x_9_n445,
         div_sub_x_9_n444, div_sub_x_9_n443, div_sub_x_9_n442,
         div_sub_x_9_n441, div_sub_x_9_n440, div_sub_x_9_n439,
         div_sub_x_9_n438, div_sub_x_9_n437, div_sub_x_9_n436,
         div_sub_x_9_n435, div_sub_x_9_n434, div_sub_x_9_n433,
         div_sub_x_9_n432, div_sub_x_9_n431, div_sub_x_9_n430,
         div_sub_x_9_n429, div_sub_x_9_n428, div_sub_x_9_n427,
         div_sub_x_9_n426, div_sub_x_9_n425, div_sub_x_9_n424,
         div_sub_x_9_n423, div_sub_x_9_n422, div_sub_x_9_n421,
         div_sub_x_9_n420, div_sub_x_9_n419, div_sub_x_9_n418,
         div_sub_x_9_n417, div_sub_x_9_n416, div_sub_x_9_n415,
         div_sub_x_9_n414, div_sub_x_9_n413, div_sub_x_9_n412,
         div_sub_x_9_n411, div_sub_x_9_n410, div_sub_x_9_n409,
         div_sub_x_9_n408, div_sub_x_9_n407, div_sub_x_9_n406,
         div_sub_x_9_n405, div_sub_x_9_n404, div_sub_x_9_n403,
         div_sub_x_9_n402, div_sub_x_9_n401, div_sub_x_9_n400,
         div_sub_x_9_n399, div_sub_x_9_n398, div_sub_x_9_n397,
         div_sub_x_9_n396, div_sub_x_9_n395, div_sub_x_9_n394,
         div_sub_x_9_n393, div_sub_x_9_n392, div_sub_x_9_n391,
         div_sub_x_9_n390, div_sub_x_9_n389, div_sub_x_9_n388,
         div_sub_x_9_n387, div_sub_x_9_n386, div_sub_x_9_n385,
         div_sub_x_9_n384, div_sub_x_9_n383, div_sub_x_9_n382,
         div_sub_x_9_n381, div_sub_x_9_n380, div_sub_x_9_n379,
         div_sub_x_9_n378, div_sub_x_9_n377, div_sub_x_9_n376,
         div_sub_x_9_n375, div_sub_x_9_n374, div_sub_x_9_n373,
         div_sub_x_9_n372, div_sub_x_9_n371, div_sub_x_9_n370,
         div_sub_x_9_n369, div_sub_x_9_n368, div_sub_x_9_n367,
         div_sub_x_9_n366, div_sub_x_9_n365, div_sub_x_9_n364,
         div_sub_x_9_n363, div_sub_x_9_n362, div_sub_x_9_n361,
         div_sub_x_9_n161, div_sub_x_7_n1116, div_sub_x_7_n1115,
         div_sub_x_7_n1114, div_sub_x_7_n1113, div_sub_x_7_n1112,
         div_sub_x_7_n1111, div_sub_x_7_n1110, div_sub_x_7_n1109,
         div_sub_x_7_n1108, div_sub_x_7_n1107, div_sub_x_7_n1106,
         div_sub_x_7_n1105, div_sub_x_7_n1104, div_sub_x_7_n1103,
         div_sub_x_7_n1102, div_sub_x_7_n1101, div_sub_x_7_n1100,
         div_sub_x_7_n1099, div_sub_x_7_n1098, div_sub_x_7_n1097,
         div_sub_x_7_n1096, div_sub_x_7_n1095, div_sub_x_7_n1094,
         div_sub_x_7_n1093, div_sub_x_7_n1092, div_sub_x_7_n1091,
         div_sub_x_7_n1090, div_sub_x_7_n1089, div_sub_x_7_n1088,
         div_sub_x_7_n1087, div_sub_x_7_n1086, div_sub_x_7_n1085,
         div_sub_x_7_n1084, div_sub_x_7_n1083, div_sub_x_7_n1082,
         div_sub_x_7_n1081, div_sub_x_7_n1080, div_sub_x_7_n1079,
         div_sub_x_7_n1078, div_sub_x_7_n1077, div_sub_x_7_n1076,
         div_sub_x_7_n1075, div_sub_x_7_n1074, div_sub_x_7_n1073,
         div_sub_x_7_n1072, div_sub_x_7_n1071, div_sub_x_7_n1070,
         div_sub_x_7_n1069, div_sub_x_7_n1068, div_sub_x_7_n1067,
         div_sub_x_7_n1066, div_sub_x_7_n1065, div_sub_x_7_n1064,
         div_sub_x_7_n1063, div_sub_x_7_n1062, div_sub_x_7_n1061,
         div_sub_x_7_n1060, div_sub_x_7_n1059, div_sub_x_7_n1058,
         div_sub_x_7_n1057, div_sub_x_7_n1056, div_sub_x_7_n1055,
         div_sub_x_7_n1054, div_sub_x_7_n1053, div_sub_x_7_n1052,
         div_sub_x_7_n1051, div_sub_x_7_n1050, div_sub_x_7_n1049,
         div_sub_x_7_n1048, div_sub_x_7_n1047, div_sub_x_7_n1046,
         div_sub_x_7_n1045, div_sub_x_7_n1044, div_sub_x_7_n1043,
         div_sub_x_7_n1042, div_sub_x_7_n1041, div_sub_x_7_n1040,
         div_sub_x_7_n1039, div_sub_x_7_n1038, div_sub_x_7_n1037,
         div_sub_x_7_n1036, div_sub_x_7_n1035, div_sub_x_7_n1034,
         div_sub_x_7_n1033, div_sub_x_7_n1032, div_sub_x_7_n1031,
         div_sub_x_7_n1030, div_sub_x_7_n1029, div_sub_x_7_n1028,
         div_sub_x_7_n1027, div_sub_x_7_n1026, div_sub_x_7_n1025,
         div_sub_x_7_n1024, div_sub_x_7_n1023, div_sub_x_7_n1022,
         div_sub_x_7_n1021, div_sub_x_7_n1020, div_sub_x_7_n1019,
         div_sub_x_7_n1018, div_sub_x_7_n1017, div_sub_x_7_n1016,
         div_sub_x_7_n1015, div_sub_x_7_n1014, div_sub_x_7_n1013,
         div_sub_x_7_n1012, div_sub_x_7_n1011, div_sub_x_7_n1010,
         div_sub_x_7_n1009, div_sub_x_7_n1008, div_sub_x_7_n1007,
         div_sub_x_7_n1006, div_sub_x_7_n1005, div_sub_x_7_n1004,
         div_sub_x_7_n1003, div_sub_x_7_n1002, div_sub_x_7_n1001,
         div_sub_x_7_n1000, div_sub_x_7_n999, div_sub_x_7_n998,
         div_sub_x_7_n997, div_sub_x_7_n996, div_sub_x_7_n995,
         div_sub_x_7_n994, div_sub_x_7_n993, div_sub_x_7_n992,
         div_sub_x_7_n991, div_sub_x_7_n990, div_sub_x_7_n989,
         div_sub_x_7_n988, div_sub_x_7_n987, div_sub_x_7_n986,
         div_sub_x_7_n985, div_sub_x_7_n984, div_sub_x_7_n983,
         div_sub_x_7_n982, div_sub_x_7_n981, div_sub_x_7_n980,
         div_sub_x_7_n979, div_sub_x_7_n978, div_sub_x_7_n977,
         div_sub_x_7_n976, div_sub_x_7_n975, div_sub_x_7_n974,
         div_sub_x_7_n973, div_sub_x_7_n972, div_sub_x_7_n971,
         div_sub_x_7_n970, div_sub_x_7_n969, div_sub_x_7_n968,
         div_sub_x_7_n967, div_sub_x_7_n966, div_sub_x_7_n965,
         div_sub_x_7_n964, div_sub_x_7_n963, div_sub_x_7_n962,
         div_sub_x_7_n961, div_sub_x_7_n960, div_sub_x_7_n959,
         div_sub_x_7_n958, div_sub_x_7_n957, div_sub_x_7_n956,
         div_sub_x_7_n955, div_sub_x_7_n954, div_sub_x_7_n953,
         div_sub_x_7_n952, div_sub_x_7_n951, div_sub_x_7_n950,
         div_sub_x_7_n949, div_sub_x_7_n948, div_sub_x_7_n947,
         div_sub_x_7_n946, div_sub_x_7_n945, div_sub_x_7_n944,
         div_sub_x_7_n943, div_sub_x_7_n942, div_sub_x_7_n941,
         div_sub_x_7_n940, div_sub_x_7_n939, div_sub_x_7_n938,
         div_sub_x_7_n937, div_sub_x_7_n936, div_sub_x_7_n935,
         div_sub_x_7_n934, div_sub_x_7_n933, div_sub_x_7_n932,
         div_sub_x_7_n931, div_sub_x_7_n930, div_sub_x_7_n929,
         div_sub_x_7_n928, div_sub_x_7_n927, div_sub_x_7_n926,
         div_sub_x_7_n925, div_sub_x_7_n924, div_sub_x_7_n923,
         div_sub_x_7_n922, div_sub_x_7_n921, div_sub_x_7_n920,
         div_sub_x_7_n919, div_sub_x_7_n918, div_sub_x_7_n917,
         div_sub_x_7_n916, div_sub_x_7_n915, div_sub_x_7_n914,
         div_sub_x_7_n913, div_sub_x_7_n912, div_sub_x_7_n911,
         div_sub_x_7_n910, div_sub_x_7_n909, div_sub_x_7_n908,
         div_sub_x_7_n907, div_sub_x_7_n906, div_sub_x_7_n905,
         div_sub_x_7_n904, div_sub_x_7_n903, div_sub_x_7_n902,
         div_sub_x_7_n901, div_sub_x_7_n900, div_sub_x_7_n899,
         div_sub_x_7_n898, div_sub_x_7_n897, div_sub_x_7_n896,
         div_sub_x_7_n895, div_sub_x_7_n894, div_sub_x_7_n893,
         div_sub_x_7_n892, div_sub_x_7_n891, div_sub_x_7_n890,
         div_sub_x_7_n889, div_sub_x_7_n888, div_sub_x_7_n887,
         div_sub_x_7_n886, div_sub_x_7_n885, div_sub_x_7_n884,
         div_sub_x_7_n883, div_sub_x_7_n882, div_sub_x_7_n881,
         div_sub_x_7_n880, div_sub_x_7_n879, div_sub_x_7_n878,
         div_sub_x_7_n877, div_sub_x_7_n876, div_sub_x_7_n875,
         div_sub_x_7_n874, div_sub_x_7_n873, div_sub_x_7_n872,
         div_sub_x_7_n871, div_sub_x_7_n870, div_sub_x_7_n869,
         div_sub_x_7_n868, div_sub_x_7_n867, div_sub_x_7_n866,
         div_sub_x_7_n865, div_sub_x_7_n864, div_sub_x_7_n863,
         div_sub_x_7_n862, div_sub_x_7_n861, div_sub_x_7_n860,
         div_sub_x_7_n859, div_sub_x_7_n858, div_sub_x_7_n857,
         div_sub_x_7_n856, div_sub_x_7_n855, div_sub_x_7_n854,
         div_sub_x_7_n853, div_sub_x_7_n852, div_sub_x_7_n851,
         div_sub_x_7_n850, div_sub_x_7_n849, div_sub_x_7_n848,
         div_sub_x_7_n847, div_sub_x_7_n846, div_sub_x_7_n845,
         div_sub_x_7_n844, div_sub_x_7_n843, div_sub_x_7_n842,
         div_sub_x_7_n841, div_sub_x_7_n840, div_sub_x_7_n839,
         div_sub_x_7_n838, div_sub_x_7_n837, div_sub_x_7_n836,
         div_sub_x_7_n835, div_sub_x_7_n834, div_sub_x_7_n833,
         div_sub_x_7_n832, div_sub_x_7_n831, div_sub_x_7_n830,
         div_sub_x_7_n829, div_sub_x_7_n828, div_sub_x_7_n827,
         div_sub_x_7_n825, div_sub_x_7_n824, div_sub_x_7_n823,
         div_sub_x_7_n822, div_sub_x_7_n820, div_sub_x_7_n819,
         div_sub_x_7_n818, div_sub_x_7_n817, div_sub_x_7_n816,
         div_sub_x_7_n815, div_sub_x_7_n813, div_sub_x_7_n812,
         div_sub_x_7_n811, div_sub_x_7_n810, div_sub_x_7_n808,
         div_sub_x_7_n807, div_sub_x_7_n806, div_sub_x_7_n805,
         div_sub_x_7_n804, div_sub_x_7_n803, div_sub_x_7_n802,
         div_sub_x_7_n801, div_sub_x_7_n800, div_sub_x_7_n799,
         div_sub_x_7_n798, div_sub_x_7_n796, div_sub_x_7_n795,
         div_sub_x_7_n794, div_sub_x_7_n793, div_sub_x_7_n792,
         div_sub_x_7_n791, div_sub_x_7_n790, div_sub_x_7_n789,
         div_sub_x_7_n788, div_sub_x_7_n787, div_sub_x_7_n786,
         div_sub_x_7_n784, div_sub_x_7_n783, div_sub_x_7_n782, add_x_94_n309,
         add_x_94_n308, add_x_94_n307, add_x_94_n306, add_x_94_n305,
         add_x_94_n304, add_x_94_n303, add_x_94_n302, add_x_94_n301,
         add_x_94_n300, add_x_94_n299, add_x_94_n298, add_x_94_n297,
         add_x_94_n296, add_x_94_n295, add_x_94_n294, add_x_94_n293,
         add_x_94_n292, add_x_94_n291, add_x_94_n290, add_x_94_n289,
         add_x_94_n288, add_x_94_n287, add_x_94_n286, add_x_94_n285,
         add_x_94_n284, add_x_94_n283, add_x_94_n282, add_x_94_n281,
         add_x_94_n280, add_x_94_n279, add_x_94_n278, add_x_94_n277,
         add_x_94_n276, add_x_94_n275, add_x_94_n274, add_x_94_n273,
         add_x_94_n272, add_x_94_n271, add_x_94_n270, add_x_94_n269,
         add_x_94_n268, add_x_94_n267, add_x_94_n266, add_x_94_n265,
         add_x_94_n264, add_x_94_n263, add_x_94_n262, add_x_94_n261,
         add_x_94_n260, add_x_94_n259, add_x_94_n258, add_x_94_n257,
         add_x_94_n256, add_x_94_n255, add_x_94_n254, add_x_94_n253,
         add_x_94_n252, add_x_94_n125, add_x_5_n504, add_x_5_n503,
         add_x_5_n502, add_x_5_n501, add_x_5_n500, add_x_5_n499, add_x_5_n498,
         add_x_5_n497, add_x_5_n496, add_x_5_n495, add_x_5_n494, add_x_5_n493,
         add_x_5_n492, add_x_5_n491, add_x_5_n490, add_x_5_n489, add_x_5_n488,
         add_x_5_n487, add_x_5_n486, add_x_5_n485, add_x_5_n484, add_x_5_n483,
         add_x_5_n482, add_x_5_n481, add_x_5_n480, add_x_5_n479, add_x_5_n478,
         add_x_5_n477, add_x_5_n476, add_x_5_n475, add_x_5_n474, add_x_5_n473,
         add_x_5_n472, add_x_5_n471, add_x_5_n470, add_x_5_n469, add_x_5_n468,
         add_x_5_n467, add_x_5_n466, add_x_5_n465, add_x_5_n464, add_x_5_n463,
         add_x_5_n462, add_x_5_n461, add_x_5_n460, add_x_5_n459, add_x_5_n458,
         add_x_5_n457, add_x_5_n456, add_x_5_n455, add_x_5_n454, add_x_5_n453,
         add_x_5_n452, add_x_5_n451, add_x_5_n450, add_x_5_n449, add_x_5_n448,
         add_x_5_n447, add_x_5_n446, add_x_5_n445, add_x_5_n444, add_x_5_n443,
         add_x_5_n442, add_x_5_n441, add_x_5_n440, add_x_5_n439, add_x_5_n438,
         add_x_5_n437, add_x_5_n436, add_x_5_n435, add_x_5_n434, add_x_5_n433,
         add_x_5_n432, add_x_5_n431, add_x_5_n430, add_x_5_n429, add_x_5_n428,
         add_x_5_n427, add_x_5_n426, add_x_5_n425, add_x_5_n424, add_x_5_n423,
         add_x_5_n422, add_x_5_n421, add_x_5_n420, add_x_5_n419, add_x_5_n418,
         add_x_5_n417, add_x_5_n416, add_x_5_n415, add_x_5_n414, add_x_5_n413,
         add_x_5_n412, add_x_5_n411, add_x_5_n410, add_x_5_n409, add_x_5_n408,
         add_x_5_n407, add_x_5_n406, add_x_5_n405, add_x_5_n404, add_x_5_n403,
         add_x_5_n402, add_x_5_n401, add_x_5_n400, add_x_5_n399, add_x_5_n398,
         add_x_5_n397, add_x_5_n396, add_x_5_n395, add_x_5_n394, add_x_5_n246;
  wire   [39:0] ibuf_io_pc;
  wire   [4:0] ibuf_io_btb_resp_entry;
  wire   [7:0] ibuf_io_btb_resp_bht_history;
  wire   [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire   [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire   [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire   [30:0] ibuf_io_inst_0_bits_raw;
  wire   [11:0] csr_io_rw_addr;
  wire   [63:0] csr_io_rw_rdata;
  wire   [12:0] csr_io_status_isa;
  wire   [39:1] csr_io_evec;
  wire   [39:0] csr_io_pc;
  wire   [39:0] csr_io_tval;
  wire   [31:0] csr_io_time;
  wire   [3:0] csr_io_interrupt_cause;
  wire   [1:0] csr_io_bp_0_control_tmatch;
  wire   [38:0] csr_io_bp_0_address;
  wire   [3:0] alu_io_fn;
  wire   [63:0] alu_io_in2;
  wire   [63:0] alu_io_in1;
  wire   [63:0] alu_io_out;
  wire   [63:0] div_io_resp_bits_data;
  wire   [4:0] div_io_resp_bits_tag;
  wire   [1942:0] n_T_427;
  wire   [63:0] n_T_427__T_1136_data;
  wire   [63:0] n_T_918;
  wire   [11:1] n_T_849;
  wire   [7:0] n_T_904;
  wire   [4:1] n_T_911;
  wire   [19:1] n_T_914;
  wire   [39:1] mem_reg_pc;
  wire   [2:0] id_ctrl_sel_imm;
  wire   [4:1] wb_waddr;
  wire   [63:1] n_T_628;
  wire   [63:1] n_T_635;
  wire   [2:0] ex_ctrl_sel_imm;
  wire   [10:0] n_T_642;
  wire   [7:0] n_T_648;
  wire   [39:0] n_T_698;
  wire   [63:0] n_T_702;
  wire   [1:0] ex_ctrl_sel_alu2;
  wire   [2:0] ex_ctrl_csr;
  wire   [2:0] mem_ctrl_csr;
  wire   [31:1] n_T_1187;
  wire   [31:0] n_T_1298;
  wire   [1:0] n_T_726;
  wire   [1:0] n_T_728;
  wire   [2:0] wb_ctrl_csr;
  wire   [63:2] id_rs_1;
  wire   [63:0] wb_cause;
  wire   [63:0] wb_reg_cause;
  wire   [63:39] n_T_1165;
  wire   [63:0] mem_reg_rs2;
  wire   [63:0] mem_reg_cause;
  wire   [7:0] ibuf_ibufBTBResp_bht_history;
  wire   [4:0] ibuf_ibufBTBResp_entry;
  wire   [39:0] ibuf_buf__pc;
  wire   [15:0] ibuf_buf__data;
  wire   [15:0] ibuf_n_T_34;
  wire   [4:0] csr_n_GEN_345;
  wire   [29:0] csr_n_GEN_307;
  wire   [29:0] csr_n_GEN_300;
  wire   [29:0] csr_n_GEN_293;
  wire   [29:0] csr_n_GEN_286;
  wire   [29:0] csr_n_GEN_279;
  wire   [29:0] csr_n_GEN_272;
  wire   [29:0] csr_n_GEN_265;
  wire   [29:0] csr_n_GEN_258;
  wire   [2:0] csr_n_GEN_155;
  wire   [63:0] csr_reg_scause;
  wire   [63:0] csr_reg_sscratch;
  wire   [63:0] csr_reg_dscratch;
  wire   [63:0] csr_reg_mcause;
  wire   [63:0] csr_reg_mscratch;
  wire   [39:0] csr_n_T_444;
  wire   [8:6] csr_n_T_389;
  wire   [39:0] csr_n_T_383;
  wire   [29:1] csr_n_T_304;
  wire   [29:1] csr_n_T_295;
  wire   [29:1] csr_n_T_286;
  wire   [29:1] csr_n_T_277;
  wire   [29:1] csr_n_T_268;
  wire   [29:1] csr_n_T_259;
  wire   [29:1] csr_n_T_250;
  wire   [29:1] csr_n_T_241;
  wire   [57:1] csr_n_T_52;
  wire   [57:1] csr_n_T_44;
  wire   [126:0] div_n_T_442;
  wire   [4:0] div_n_T_429;
  wire   [4:0] div_n_T_272;
  wire   [63:0] div_n_T_87;
  wire   [72:0] div_n_T_65;
  wire   [63:1] div_negated_remainder;
  assign io_ptw_sfence_valid = io_imem_sfence_valid;
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1;
  assign io_ptw_sfence_bits_rs2 = io_imem_sfence_bits_rs2;
  assign io_ptw_sfence_bits_addr[38] = io_imem_sfence_bits_addr[38];
  assign io_ptw_sfence_bits_addr[37] = io_imem_sfence_bits_addr[37];
  assign io_ptw_sfence_bits_addr[36] = io_imem_sfence_bits_addr[36];
  assign io_ptw_sfence_bits_addr[35] = io_imem_sfence_bits_addr[35];
  assign io_ptw_sfence_bits_addr[34] = io_imem_sfence_bits_addr[34];
  assign io_ptw_sfence_bits_addr[33] = io_imem_sfence_bits_addr[33];
  assign io_ptw_sfence_bits_addr[32] = io_imem_sfence_bits_addr[32];
  assign io_ptw_sfence_bits_addr[31] = io_imem_sfence_bits_addr[31];
  assign io_ptw_sfence_bits_addr[30] = io_imem_sfence_bits_addr[30];
  assign io_ptw_sfence_bits_addr[29] = io_imem_sfence_bits_addr[29];
  assign io_ptw_sfence_bits_addr[28] = io_imem_sfence_bits_addr[28];
  assign io_ptw_sfence_bits_addr[27] = io_imem_sfence_bits_addr[27];
  assign io_ptw_sfence_bits_addr[26] = io_imem_sfence_bits_addr[26];
  assign io_ptw_sfence_bits_addr[25] = io_imem_sfence_bits_addr[25];
  assign io_ptw_sfence_bits_addr[24] = io_imem_sfence_bits_addr[24];
  assign io_ptw_sfence_bits_addr[23] = io_imem_sfence_bits_addr[23];
  assign io_ptw_sfence_bits_addr[22] = io_imem_sfence_bits_addr[22];
  assign io_ptw_sfence_bits_addr[21] = io_imem_sfence_bits_addr[21];
  assign io_ptw_sfence_bits_addr[20] = io_imem_sfence_bits_addr[20];
  assign io_ptw_sfence_bits_addr[19] = io_imem_sfence_bits_addr[19];
  assign io_ptw_sfence_bits_addr[18] = io_imem_sfence_bits_addr[18];
  assign io_ptw_sfence_bits_addr[17] = io_imem_sfence_bits_addr[17];
  assign io_ptw_sfence_bits_addr[16] = io_imem_sfence_bits_addr[16];
  assign io_ptw_sfence_bits_addr[15] = io_imem_sfence_bits_addr[15];
  assign io_ptw_sfence_bits_addr[14] = io_imem_sfence_bits_addr[14];
  assign io_ptw_sfence_bits_addr[13] = io_imem_sfence_bits_addr[13];
  assign io_ptw_sfence_bits_addr[12] = io_imem_sfence_bits_addr[12];
  assign io_ptw_sfence_bits_addr[11] = io_imem_sfence_bits_addr[11];
  assign io_ptw_sfence_bits_addr[10] = io_imem_sfence_bits_addr[10];
  assign io_ptw_sfence_bits_addr[9] = io_imem_sfence_bits_addr[9];
  assign io_ptw_sfence_bits_addr[8] = io_imem_sfence_bits_addr[8];
  assign io_ptw_sfence_bits_addr[7] = io_imem_sfence_bits_addr[7];
  assign io_ptw_sfence_bits_addr[6] = io_imem_sfence_bits_addr[6];
  assign io_ptw_sfence_bits_addr[5] = io_imem_sfence_bits_addr[5];
  assign io_ptw_sfence_bits_addr[4] = io_imem_sfence_bits_addr[4];
  assign io_ptw_sfence_bits_addr[3] = io_imem_sfence_bits_addr[3];
  assign io_ptw_sfence_bits_addr[2] = io_imem_sfence_bits_addr[2];
  assign io_ptw_sfence_bits_addr[1] = io_imem_sfence_bits_addr[1];
  assign io_ptw_sfence_bits_addr[0] = io_imem_sfence_bits_addr[0];
  assign io_imem_bht_update_bits_pc[38] = io_imem_btb_update_bits_br_pc[38];
  assign io_imem_btb_update_bits_pc[38] = io_imem_btb_update_bits_br_pc[38];
  assign io_imem_bht_update_bits_pc[37] = io_imem_btb_update_bits_br_pc[37];
  assign io_imem_btb_update_bits_pc[37] = io_imem_btb_update_bits_br_pc[37];
  assign io_imem_bht_update_bits_pc[36] = io_imem_btb_update_bits_br_pc[36];
  assign io_imem_btb_update_bits_pc[36] = io_imem_btb_update_bits_br_pc[36];
  assign io_imem_bht_update_bits_pc[35] = io_imem_btb_update_bits_br_pc[35];
  assign io_imem_btb_update_bits_pc[35] = io_imem_btb_update_bits_br_pc[35];
  assign io_imem_bht_update_bits_pc[34] = io_imem_btb_update_bits_br_pc[34];
  assign io_imem_btb_update_bits_pc[34] = io_imem_btb_update_bits_br_pc[34];
  assign io_imem_bht_update_bits_pc[33] = io_imem_btb_update_bits_br_pc[33];
  assign io_imem_btb_update_bits_pc[33] = io_imem_btb_update_bits_br_pc[33];
  assign io_imem_bht_update_bits_pc[32] = io_imem_btb_update_bits_br_pc[32];
  assign io_imem_btb_update_bits_pc[32] = io_imem_btb_update_bits_br_pc[32];
  assign io_imem_bht_update_bits_pc[31] = io_imem_btb_update_bits_br_pc[31];
  assign io_imem_btb_update_bits_pc[31] = io_imem_btb_update_bits_br_pc[31];
  assign io_imem_bht_update_bits_pc[30] = io_imem_btb_update_bits_br_pc[30];
  assign io_imem_btb_update_bits_pc[30] = io_imem_btb_update_bits_br_pc[30];
  assign io_imem_bht_update_bits_pc[29] = io_imem_btb_update_bits_br_pc[29];
  assign io_imem_btb_update_bits_pc[29] = io_imem_btb_update_bits_br_pc[29];
  assign io_imem_bht_update_bits_pc[28] = io_imem_btb_update_bits_br_pc[28];
  assign io_imem_btb_update_bits_pc[28] = io_imem_btb_update_bits_br_pc[28];
  assign io_imem_bht_update_bits_pc[27] = io_imem_btb_update_bits_br_pc[27];
  assign io_imem_btb_update_bits_pc[27] = io_imem_btb_update_bits_br_pc[27];
  assign io_imem_bht_update_bits_pc[26] = io_imem_btb_update_bits_br_pc[26];
  assign io_imem_btb_update_bits_pc[26] = io_imem_btb_update_bits_br_pc[26];
  assign io_imem_bht_update_bits_pc[25] = io_imem_btb_update_bits_br_pc[25];
  assign io_imem_btb_update_bits_pc[25] = io_imem_btb_update_bits_br_pc[25];
  assign io_imem_bht_update_bits_pc[24] = io_imem_btb_update_bits_br_pc[24];
  assign io_imem_btb_update_bits_pc[24] = io_imem_btb_update_bits_br_pc[24];
  assign io_imem_bht_update_bits_pc[23] = io_imem_btb_update_bits_br_pc[23];
  assign io_imem_btb_update_bits_pc[23] = io_imem_btb_update_bits_br_pc[23];
  assign io_imem_bht_update_bits_pc[22] = io_imem_btb_update_bits_br_pc[22];
  assign io_imem_btb_update_bits_pc[22] = io_imem_btb_update_bits_br_pc[22];
  assign io_imem_bht_update_bits_pc[21] = io_imem_btb_update_bits_br_pc[21];
  assign io_imem_btb_update_bits_pc[21] = io_imem_btb_update_bits_br_pc[21];
  assign io_imem_bht_update_bits_pc[20] = io_imem_btb_update_bits_br_pc[20];
  assign io_imem_btb_update_bits_pc[20] = io_imem_btb_update_bits_br_pc[20];
  assign io_imem_bht_update_bits_pc[19] = io_imem_btb_update_bits_br_pc[19];
  assign io_imem_btb_update_bits_pc[19] = io_imem_btb_update_bits_br_pc[19];
  assign io_imem_bht_update_bits_pc[18] = io_imem_btb_update_bits_br_pc[18];
  assign io_imem_btb_update_bits_pc[18] = io_imem_btb_update_bits_br_pc[18];
  assign io_imem_bht_update_bits_pc[17] = io_imem_btb_update_bits_br_pc[17];
  assign io_imem_btb_update_bits_pc[17] = io_imem_btb_update_bits_br_pc[17];
  assign io_imem_bht_update_bits_pc[16] = io_imem_btb_update_bits_br_pc[16];
  assign io_imem_btb_update_bits_pc[16] = io_imem_btb_update_bits_br_pc[16];
  assign io_imem_bht_update_bits_pc[15] = io_imem_btb_update_bits_br_pc[15];
  assign io_imem_btb_update_bits_pc[15] = io_imem_btb_update_bits_br_pc[15];
  assign io_imem_bht_update_bits_pc[14] = io_imem_btb_update_bits_br_pc[14];
  assign io_imem_btb_update_bits_pc[14] = io_imem_btb_update_bits_br_pc[14];
  assign io_imem_bht_update_bits_pc[13] = io_imem_btb_update_bits_br_pc[13];
  assign io_imem_btb_update_bits_pc[13] = io_imem_btb_update_bits_br_pc[13];
  assign io_imem_bht_update_bits_pc[12] = io_imem_btb_update_bits_br_pc[12];
  assign io_imem_btb_update_bits_pc[12] = io_imem_btb_update_bits_br_pc[12];
  assign io_imem_bht_update_bits_pc[11] = io_imem_btb_update_bits_br_pc[11];
  assign io_imem_btb_update_bits_pc[11] = io_imem_btb_update_bits_br_pc[11];
  assign io_imem_bht_update_bits_pc[10] = io_imem_btb_update_bits_br_pc[10];
  assign io_imem_btb_update_bits_pc[10] = io_imem_btb_update_bits_br_pc[10];
  assign io_imem_bht_update_bits_pc[9] = io_imem_btb_update_bits_br_pc[9];
  assign io_imem_btb_update_bits_pc[9] = io_imem_btb_update_bits_br_pc[9];
  assign io_imem_bht_update_bits_pc[8] = io_imem_btb_update_bits_br_pc[8];
  assign io_imem_btb_update_bits_pc[8] = io_imem_btb_update_bits_br_pc[8];
  assign io_imem_bht_update_bits_pc[7] = io_imem_btb_update_bits_br_pc[7];
  assign io_imem_btb_update_bits_pc[7] = io_imem_btb_update_bits_br_pc[7];
  assign io_imem_bht_update_bits_pc[6] = io_imem_btb_update_bits_br_pc[6];
  assign io_imem_btb_update_bits_pc[6] = io_imem_btb_update_bits_br_pc[6];
  assign io_imem_bht_update_bits_pc[5] = io_imem_btb_update_bits_br_pc[5];
  assign io_imem_btb_update_bits_pc[5] = io_imem_btb_update_bits_br_pc[5];
  assign io_imem_bht_update_bits_pc[4] = io_imem_btb_update_bits_br_pc[4];
  assign io_imem_btb_update_bits_pc[4] = io_imem_btb_update_bits_br_pc[4];
  assign io_imem_bht_update_bits_pc[3] = io_imem_btb_update_bits_br_pc[3];
  assign io_imem_btb_update_bits_pc[3] = io_imem_btb_update_bits_br_pc[3];
  assign io_imem_bht_update_bits_pc[2] = io_imem_btb_update_bits_br_pc[2];
  assign io_imem_btb_update_bits_pc[2] = io_imem_btb_update_bits_br_pc[2];
  assign io_ptw_status_dprv[1] = io_dmem_req_bits_dprv[1];
  assign io_ptw_status_dprv[0] = io_dmem_req_bits_dprv[0];
  assign io_ptw_pmp_0_mask[2] = io_ptw_pmp_0_cfg_a[0];
  assign io_ptw_pmp_1_mask[2] = io_ptw_pmp_1_cfg_a[0];
  assign io_ptw_pmp_2_mask[2] = io_ptw_pmp_2_cfg_a[0];
  assign io_ptw_pmp_3_mask[2] = io_ptw_pmp_3_cfg_a[0];
  assign io_ptw_pmp_4_mask[2] = io_ptw_pmp_4_cfg_a[0];
  assign io_ptw_pmp_5_mask[2] = io_ptw_pmp_5_cfg_a[0];
  assign io_ptw_pmp_6_mask[2] = io_ptw_pmp_6_cfg_a[0];
  assign io_ptw_pmp_7_mask[2] = io_ptw_pmp_7_cfg_a[0];
  assign io_dmem_req_bits_tag[6] = 1'b0;
  assign io_fpu_dmem_resp_type[2] = 1'b0;
  assign io_imem_btb_update_bits_pc[1] = 1'b0;
  assign io_imem_btb_update_bits_pc[0] = 1'b0;
  assign io_imem_bht_update_bits_pc[1] = 1'b0;
  assign io_imem_bht_update_bits_pc[0] = 1'b0;
  assign io_ptw_ptbr_mode[0] = 1'b0;
  assign io_ptw_ptbr_mode[1] = 1'b0;
  assign io_ptw_ptbr_mode[2] = 1'b0;
  assign io_ptw_ptbr_ppn[20] = 1'b0;
  assign io_ptw_ptbr_ppn[21] = 1'b0;
  assign io_ptw_ptbr_ppn[22] = 1'b0;
  assign io_ptw_ptbr_ppn[23] = 1'b0;
  assign io_ptw_ptbr_ppn[24] = 1'b0;
  assign io_ptw_ptbr_ppn[25] = 1'b0;
  assign io_ptw_ptbr_ppn[26] = 1'b0;
  assign io_ptw_ptbr_ppn[27] = 1'b0;
  assign io_ptw_ptbr_ppn[28] = 1'b0;
  assign io_ptw_ptbr_ppn[29] = 1'b0;
  assign io_ptw_ptbr_ppn[30] = 1'b0;
  assign io_ptw_ptbr_ppn[31] = 1'b0;
  assign io_ptw_ptbr_ppn[32] = 1'b0;
  assign io_ptw_ptbr_ppn[33] = 1'b0;
  assign io_ptw_ptbr_ppn[34] = 1'b0;
  assign io_ptw_ptbr_ppn[35] = 1'b0;
  assign io_ptw_ptbr_ppn[36] = 1'b0;
  assign io_ptw_ptbr_ppn[37] = 1'b0;
  assign io_ptw_ptbr_ppn[38] = 1'b0;
  assign io_ptw_ptbr_ppn[39] = 1'b0;
  assign io_ptw_ptbr_ppn[40] = 1'b0;
  assign io_ptw_ptbr_ppn[41] = 1'b0;
  assign io_ptw_ptbr_ppn[42] = 1'b0;
  assign io_ptw_ptbr_ppn[43] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[0] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[1] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[2] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[4] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[5] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[6] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[7] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[8] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[10] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[11] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[12] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[13] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[14] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[15] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[16] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[17] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[18] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[19] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[20] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[21] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[22] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[23] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[24] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[25] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[26] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[27] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[28] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[29] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[30] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[31] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[32] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[33] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[34] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[35] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[36] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[37] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[38] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[39] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[40] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[41] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[42] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[43] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[44] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[45] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[46] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[47] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[48] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[49] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[50] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[51] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[52] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[53] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[54] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[55] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[56] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[57] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[58] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[59] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[60] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[61] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[62] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[63] = 1'b0;
  assign io_ptw_pmp_0_mask[1] = 1'b1;
  assign io_ptw_pmp_0_mask[0] = 1'b1;
  assign io_ptw_pmp_1_mask[1] = 1'b1;
  assign io_ptw_pmp_1_mask[0] = 1'b1;
  assign io_ptw_pmp_2_mask[1] = 1'b1;
  assign io_ptw_pmp_2_mask[0] = 1'b1;
  assign io_ptw_pmp_3_mask[1] = 1'b1;
  assign io_ptw_pmp_3_mask[0] = 1'b1;
  assign io_ptw_pmp_4_mask[1] = 1'b1;
  assign io_ptw_pmp_4_mask[0] = 1'b1;
  assign io_ptw_pmp_5_mask[1] = 1'b1;
  assign io_ptw_pmp_5_mask[0] = 1'b1;
  assign io_ptw_pmp_6_mask[1] = 1'b1;
  assign io_ptw_pmp_6_mask[0] = 1'b1;
  assign io_ptw_pmp_7_mask[1] = 1'b1;
  assign io_ptw_pmp_7_mask[0] = 1'b1;
  assign io_fpu_inst[1] = 1'b1;
  assign io_fpu_inst[0] = 1'b1;
  assign io_fpu_dmem_resp_type[1] = io_dmem_resp_bits_size[1];
  assign io_fpu_dmem_resp_type[0] = io_dmem_resp_bits_size[0];
  assign io_fpu_dmem_resp_tag[4] = io_dmem_resp_bits_tag[5];
  assign io_fpu_dmem_resp_tag[3] = io_dmem_resp_bits_tag[4];
  assign io_fpu_dmem_resp_tag[2] = io_dmem_resp_bits_tag[3];
  assign io_fpu_dmem_resp_tag[1] = io_dmem_resp_bits_tag[2];
  assign io_fpu_dmem_resp_tag[0] = io_dmem_resp_bits_tag[1];
  assign io_fpu_dmem_resp_data[63] = io_dmem_resp_bits_data_word_bypass[63];
  assign io_fpu_dmem_resp_data[62] = io_dmem_resp_bits_data_word_bypass[62];
  assign io_fpu_dmem_resp_data[61] = io_dmem_resp_bits_data_word_bypass[61];
  assign io_fpu_dmem_resp_data[60] = io_dmem_resp_bits_data_word_bypass[60];
  assign io_fpu_dmem_resp_data[59] = io_dmem_resp_bits_data_word_bypass[59];
  assign io_fpu_dmem_resp_data[58] = io_dmem_resp_bits_data_word_bypass[58];
  assign io_fpu_dmem_resp_data[57] = io_dmem_resp_bits_data_word_bypass[57];
  assign io_fpu_dmem_resp_data[56] = io_dmem_resp_bits_data_word_bypass[56];
  assign io_fpu_dmem_resp_data[55] = io_dmem_resp_bits_data_word_bypass[55];
  assign io_fpu_dmem_resp_data[54] = io_dmem_resp_bits_data_word_bypass[54];
  assign io_fpu_dmem_resp_data[53] = io_dmem_resp_bits_data_word_bypass[53];
  assign io_fpu_dmem_resp_data[52] = io_dmem_resp_bits_data_word_bypass[52];
  assign io_fpu_dmem_resp_data[51] = io_dmem_resp_bits_data_word_bypass[51];
  assign io_fpu_dmem_resp_data[50] = io_dmem_resp_bits_data_word_bypass[50];
  assign io_fpu_dmem_resp_data[49] = io_dmem_resp_bits_data_word_bypass[49];
  assign io_fpu_dmem_resp_data[48] = io_dmem_resp_bits_data_word_bypass[48];
  assign io_fpu_dmem_resp_data[47] = io_dmem_resp_bits_data_word_bypass[47];
  assign io_fpu_dmem_resp_data[46] = io_dmem_resp_bits_data_word_bypass[46];
  assign io_fpu_dmem_resp_data[45] = io_dmem_resp_bits_data_word_bypass[45];
  assign io_fpu_dmem_resp_data[44] = io_dmem_resp_bits_data_word_bypass[44];
  assign io_fpu_dmem_resp_data[43] = io_dmem_resp_bits_data_word_bypass[43];
  assign io_fpu_dmem_resp_data[42] = io_dmem_resp_bits_data_word_bypass[42];
  assign io_fpu_dmem_resp_data[41] = io_dmem_resp_bits_data_word_bypass[41];
  assign io_fpu_dmem_resp_data[40] = io_dmem_resp_bits_data_word_bypass[40];
  assign io_fpu_dmem_resp_data[39] = io_dmem_resp_bits_data_word_bypass[39];
  assign io_fpu_dmem_resp_data[38] = io_dmem_resp_bits_data_word_bypass[38];
  assign io_fpu_dmem_resp_data[37] = io_dmem_resp_bits_data_word_bypass[37];
  assign io_fpu_dmem_resp_data[36] = io_dmem_resp_bits_data_word_bypass[36];
  assign io_fpu_dmem_resp_data[35] = io_dmem_resp_bits_data_word_bypass[35];
  assign io_fpu_dmem_resp_data[34] = io_dmem_resp_bits_data_word_bypass[34];
  assign io_fpu_dmem_resp_data[33] = io_dmem_resp_bits_data_word_bypass[33];
  assign io_fpu_dmem_resp_data[32] = io_dmem_resp_bits_data_word_bypass[32];
  assign io_fpu_dmem_resp_data[31] = io_dmem_resp_bits_data_word_bypass[31];
  assign io_fpu_dmem_resp_data[30] = io_dmem_resp_bits_data_word_bypass[30];
  assign io_fpu_dmem_resp_data[29] = io_dmem_resp_bits_data_word_bypass[29];
  assign io_fpu_dmem_resp_data[28] = io_dmem_resp_bits_data_word_bypass[28];
  assign io_fpu_dmem_resp_data[27] = io_dmem_resp_bits_data_word_bypass[27];
  assign io_fpu_dmem_resp_data[26] = io_dmem_resp_bits_data_word_bypass[26];
  assign io_fpu_dmem_resp_data[25] = io_dmem_resp_bits_data_word_bypass[25];
  assign io_fpu_dmem_resp_data[24] = io_dmem_resp_bits_data_word_bypass[24];
  assign io_fpu_dmem_resp_data[23] = io_dmem_resp_bits_data_word_bypass[23];
  assign io_fpu_dmem_resp_data[22] = io_dmem_resp_bits_data_word_bypass[22];
  assign io_fpu_dmem_resp_data[21] = io_dmem_resp_bits_data_word_bypass[21];
  assign io_fpu_dmem_resp_data[20] = io_dmem_resp_bits_data_word_bypass[20];
  assign io_fpu_dmem_resp_data[19] = io_dmem_resp_bits_data_word_bypass[19];
  assign io_fpu_dmem_resp_data[18] = io_dmem_resp_bits_data_word_bypass[18];
  assign io_fpu_dmem_resp_data[17] = io_dmem_resp_bits_data_word_bypass[17];
  assign io_fpu_dmem_resp_data[16] = io_dmem_resp_bits_data_word_bypass[16];
  assign io_fpu_dmem_resp_data[15] = io_dmem_resp_bits_data_word_bypass[15];
  assign io_fpu_dmem_resp_data[14] = io_dmem_resp_bits_data_word_bypass[14];
  assign io_fpu_dmem_resp_data[13] = io_dmem_resp_bits_data_word_bypass[13];
  assign io_fpu_dmem_resp_data[12] = io_dmem_resp_bits_data_word_bypass[12];
  assign io_fpu_dmem_resp_data[11] = io_dmem_resp_bits_data_word_bypass[11];
  assign io_fpu_dmem_resp_data[10] = io_dmem_resp_bits_data_word_bypass[10];
  assign io_fpu_dmem_resp_data[9] = io_dmem_resp_bits_data_word_bypass[9];
  assign io_fpu_dmem_resp_data[8] = io_dmem_resp_bits_data_word_bypass[8];
  assign io_fpu_dmem_resp_data[7] = io_dmem_resp_bits_data_word_bypass[7];
  assign io_fpu_dmem_resp_data[6] = io_dmem_resp_bits_data_word_bypass[6];
  assign io_fpu_dmem_resp_data[5] = io_dmem_resp_bits_data_word_bypass[5];
  assign io_fpu_dmem_resp_data[4] = io_dmem_resp_bits_data_word_bypass[4];
  assign io_fpu_dmem_resp_data[3] = io_dmem_resp_bits_data_word_bypass[3];
  assign io_fpu_dmem_resp_data[2] = io_dmem_resp_bits_data_word_bypass[2];
  assign io_fpu_dmem_resp_data[1] = io_dmem_resp_bits_data_word_bypass[1];
  assign io_fpu_dmem_resp_data[0] = io_dmem_resp_bits_data_word_bypass[0];

  PlusArgTimeout PlusArgTimeout ( .clock(n3595), .reset(reset), .io_count(
        csr_io_time) );
  SNPS_CLOCK_GATE_HIGH_Rocket_0 clk_gate_ex_reg_rs_bypass_1_reg ( .CLK(n3595), 
        .EN(n406), .ENCLK(net34469), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_39 clk_gate_wb_ctrl_wxd_reg ( .CLK(n4499), .EN(
        mem_pc_valid), .ENCLK(net34475), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_38 clk_gate_mem_ctrl_branch_reg ( .CLK(n4499), 
        .EN(N290), .ENCLK(net34480), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_37 clk_gate__T_427_reg_0_ ( .CLK(n3595), .EN(
        N268), .ENCLK(net34485), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_36 clk_gate__T_427_reg_1_ ( .CLK(n3595), .EN(
        N267), .ENCLK(net34490), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_35 clk_gate__T_427_reg_2_ ( .CLK(n3595), .EN(
        N266), .ENCLK(net34495), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_34 clk_gate__T_427_reg_3_ ( .CLK(n3595), .EN(
        N265), .ENCLK(net34500), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_33 clk_gate__T_427_reg_4_ ( .CLK(n3595), .EN(
        N264), .ENCLK(net34505), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_32 clk_gate__T_427_reg_5_ ( .CLK(n3595), .EN(
        N263), .ENCLK(net34510), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_31 clk_gate__T_427_reg_6_ ( .CLK(n3595), .EN(
        N262), .ENCLK(net34515), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_30 clk_gate__T_427_reg_7_ ( .CLK(n3785), .EN(
        N261), .ENCLK(net34520), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_29 clk_gate__T_427_reg_8_ ( .CLK(n3594), .EN(
        N260), .ENCLK(net34525), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_28 clk_gate__T_427_reg_9_ ( .CLK(n3785), .EN(
        N259), .ENCLK(net34530), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_27 clk_gate__T_427_reg_10_ ( .CLK(n4499), .EN(
        N258), .ENCLK(net34535), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_26 clk_gate__T_427_reg_11_ ( .CLK(n3785), .EN(
        N257), .ENCLK(net34540), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_25 clk_gate__T_427_reg_12_ ( .CLK(n4499), .EN(
        N256), .ENCLK(net34545), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_24 clk_gate__T_427_reg_13_ ( .CLK(n3785), .EN(
        N255), .ENCLK(net34550), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_23 clk_gate__T_427_reg_14_ ( .CLK(n4499), .EN(
        N254), .ENCLK(net34555), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_22 clk_gate__T_427_reg_15_ ( .CLK(n3785), .EN(
        N253), .ENCLK(net34560), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_21 clk_gate__T_427_reg_16_ ( .CLK(n4499), .EN(
        N252), .ENCLK(net34565), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_20 clk_gate__T_427_reg_17_ ( .CLK(n3595), .EN(
        N251), .ENCLK(net34570), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_19 clk_gate__T_427_reg_18_ ( .CLK(n3594), .EN(
        N250), .ENCLK(net34575), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_18 clk_gate__T_427_reg_19_ ( .CLK(n3785), .EN(
        N249), .ENCLK(net34580), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_17 clk_gate__T_427_reg_20_ ( .CLK(n4499), .EN(
        N248), .ENCLK(net34585), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_16 clk_gate__T_427_reg_21_ ( .CLK(n3785), .EN(
        N247), .ENCLK(net34590), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_15 clk_gate__T_427_reg_22_ ( .CLK(n4499), .EN(
        N246), .ENCLK(net34595), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_14 clk_gate__T_427_reg_23_ ( .CLK(n3785), .EN(
        N245), .ENCLK(net34600), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_13 clk_gate__T_427_reg_24_ ( .CLK(n4499), .EN(
        N244), .ENCLK(net34605), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_12 clk_gate__T_427_reg_25_ ( .CLK(n3785), .EN(
        N243), .ENCLK(net34610), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_11 clk_gate__T_427_reg_26_ ( .CLK(n4499), .EN(
        N242), .ENCLK(net34615), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_10 clk_gate__T_427_reg_27_ ( .CLK(n3785), .EN(
        N241), .ENCLK(net34620), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_9 clk_gate__T_427_reg_28_ ( .CLK(n4499), .EN(
        N240), .ENCLK(net34625), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_8 clk_gate__T_427_reg_29_ ( .CLK(n3785), .EN(
        N239), .ENCLK(net34630), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_7 clk_gate__T_427_reg_30_ ( .CLK(n4499), .EN(
        N238), .ENCLK(net34635), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_6 clk_gate_ex_reg_btb_resp_bht_history_reg ( 
        .CLK(n3785), .EN(n_T_760), .ENCLK(net34640), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_5 clk_gate_mem_reg_rs2_reg ( .CLK(n4499), .EN(
        N526), .ENCLK(net34645), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_4 clk_gate_ex_reg_rs_msb_0_reg ( .CLK(n3594), 
        .EN(N744), .ENCLK(net34650), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_3 clk_gate_ex_reg_rs_msb_1_reg ( .CLK(n3785), 
        .EN(N745), .ENCLK(net34655), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_2 clk_gate__T_1185_reg ( .CLK(clock), .EN(N746), 
        .ENCLK(net34660), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_1 clk_gate__T_1298_reg ( .CLK(n3595), .EN(N778), 
        .ENCLK(net34665), .TE(1'b0) );
  DFFX1_LVT mem_reg_inst_reg_7_ ( .D(n592), .CLK(n4286), .Q(n3202), .QN(
        n_T_849[11]) );
  DFFX1_LVT ex_reg_valid_reg ( .D(n2874), .CLK(n3594), .QN(ex_reg_valid) );
  DFFX1_LVT mem_reg_valid_reg ( .D(io_fpu_killx), .CLK(n3594), .Q(n3206), .QN(
        mem_reg_valid) );
  DFFX1_LVT wb_reg_wdata_reg_0_ ( .D(N598), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[0]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_61_ ( .D(id_rs_1[63]), .CLK(n4079), .Q(
        n_T_635[63]) );
  DFFX1_LVT mem_reg_wdata_reg_63_ ( .D(alu_io_out[63]), .CLK(n4293), .Q(
        n_T_918[63]) );
  DFFSSRX1_LVT mem_reg_replay_reg ( .D(n9421), .SETB(n9418), .RSTB(1'b1), 
        .CLK(n3594), .QN(mem_reg_replay) );
  DFFX1_LVT wb_reg_replay_reg ( .D(N530), .CLK(n3594), .Q(wb_reg_replay) );
  DFFX1_LVT ex_ctrl_sel_imm_reg_1_ ( .D(id_ctrl_sel_imm[1]), .CLK(n4312), .QN(
        n546) );
  DFFX1_LVT ex_ctrl_mem_cmd_reg_4_ ( .D(n1891), .CLK(n4315), .Q(
        io_dmem_req_bits_cmd[4]), .QN(n3245) );
  DFFX1_LVT ex_ctrl_jal_reg ( .D(n9428), .CLK(n4315), .Q(ex_ctrl_jal) );
  DFFX1_LVT ex_ctrl_branch_reg ( .D(n9429), .CLK(n4315), .QN(n323) );
  DFFX1_LVT ex_ctrl_sel_imm_reg_0_ ( .D(id_ctrl_sel_imm[0]), .CLK(n4315), .Q(
        ex_ctrl_sel_imm[0]) );
  DFFX1_LVT ex_ctrl_csr_reg_0_ ( .D(N286), .CLK(n4315), .Q(ex_ctrl_csr[0]), 
        .QN(n320) );
  DFFX1_LVT ex_ctrl_csr_reg_1_ ( .D(n1628), .CLK(n4314), .Q(n319), .QN(
        ex_ctrl_csr[1]) );
  DFFX1_LVT ex_ctrl_fence_i_reg ( .D(n1828), .CLK(n4314), .QN(n318) );
  DFFX1_LVT ex_ctrl_sel_imm_reg_2_ ( .D(id_ctrl_sel_imm[2]), .CLK(n4314), .Q(
        ex_ctrl_sel_imm[2]), .QN(n3231) );
  DFFX1_LVT ex_ctrl_jalr_reg ( .D(n1823), .CLK(n4314), .Q(ex_ctrl_jalr), .QN(
        n2495) );
  DFFX1_LVT id_reg_pause_reg ( .D(n1820), .CLK(n3594), .Q(id_reg_pause) );
  DFFX1_LVT ex_ctrl_div_reg ( .D(n9413), .CLK(n4314), .Q(n317), .QN(
        ex_ctrl_div) );
  DFFX1_LVT ex_ctrl_mem_cmd_reg_0_ ( .D(n9431), .CLK(n4314), .Q(
        io_dmem_req_bits_cmd[0]), .QN(n560) );
  DFFSSRX1_LVT ex_ctrl_rxs2_reg ( .D(n1531), .SETB(1'b1), .RSTB(n1532), .CLK(
        n4312), .QN(ex_ctrl_rxs2) );
  DFFX1_LVT ex_ctrl_wfd_reg ( .D(id_ctrl_wfd), .CLK(n4314), .Q(ex_ctrl_wfd), 
        .QN(n315) );
  DFFX1_LVT ex_ctrl_wxd_reg ( .D(id_ctrl_wxd), .CLK(n4314), .Q(ex_ctrl_wxd), 
        .QN(n314) );
  DFFX1_LVT ex_ctrl_mem_cmd_reg_2_ ( .D(id_ctrl_mem_cmd_2_), .CLK(n4314), .Q(
        io_dmem_req_bits_cmd[2]), .QN(n3244) );
  DFFX1_LVT ex_reg_mem_size_reg_0_ ( .D(N369), .CLK(n4314), .Q(
        io_dmem_req_bits_size[0]), .QN(n313) );
  DFFX1_LVT id_reg_fence_reg ( .D(n1821), .CLK(n3595), .Q(id_reg_fence) );
  DFFX1_LVT blocked_reg ( .D(N811), .CLK(n3594), .Q(blocked) );
  DFFSSRX1_LVT ex_ctrl_csr_reg_2_ ( .D(n1628), .SETB(n2569), .RSTB(n2131), 
        .CLK(n4312), .Q(ex_ctrl_csr[2]), .QN(n310) );
  DFFX1_LVT ex_reg_flush_pipe_reg ( .D(n_T_731), .CLK(n4313), .QN(n309) );
  DFFX1_LVT ex_reg_inst_reg_31_ ( .D(n9434), .CLK(n4098), .Q(n172), .QN(
        ex_reg_inst_31_) );
  DFFX1_LVT ex_reg_inst_reg_30_ ( .D(n9435), .CLK(n4098), .Q(n171), .QN(
        n_T_642[10]) );
  DFFX1_LVT ex_reg_inst_reg_29_ ( .D(n9436), .CLK(n4098), .Q(n170), .QN(
        n_T_642[9]) );
  DFFX1_LVT ex_reg_inst_reg_28_ ( .D(n9437), .CLK(n4098), .Q(n169), .QN(
        n_T_642[8]) );
  DFFX1_LVT ex_reg_inst_reg_27_ ( .D(n9438), .CLK(n4098), .Q(n168), .QN(
        n_T_642[7]) );
  DFFX1_LVT ex_reg_inst_reg_26_ ( .D(n9439), .CLK(n4098), .Q(n167), .QN(
        n_T_642[6]) );
  DFFX1_LVT ex_reg_inst_reg_25_ ( .D(n9440), .CLK(n4098), .Q(n166), .QN(
        n_T_642[5]) );
  DFFX1_LVT ex_reg_inst_reg_24_ ( .D(io_fpu_inst[24]), .CLK(n4098), .Q(
        n_T_642[4]), .QN(n165) );
  DFFX1_LVT ex_reg_inst_reg_23_ ( .D(n9441), .CLK(n4098), .Q(n164), .QN(
        n_T_642[3]) );
  DFFX1_LVT ex_reg_inst_reg_22_ ( .D(n9442), .CLK(n4098), .Q(n163), .QN(
        n_T_642[2]) );
  DFFX1_LVT ex_reg_inst_reg_21_ ( .D(n9443), .CLK(n4098), .Q(n162), .QN(
        n_T_642[1]) );
  DFFX1_LVT ex_reg_inst_reg_20_ ( .D(n9444), .CLK(n4097), .Q(n161), .QN(
        n_T_642[0]) );
  DFFX1_LVT ex_reg_inst_reg_19_ ( .D(io_fpu_inst[19]), .CLK(n4097), .Q(
        n_T_648[7]), .QN(n160) );
  DFFX1_LVT ex_reg_inst_reg_18_ ( .D(io_fpu_inst[18]), .CLK(n4097), .Q(
        n_T_648[6]), .QN(n159) );
  DFFX1_LVT ex_reg_inst_reg_17_ ( .D(io_fpu_inst[17]), .CLK(n4097), .Q(
        n_T_648[5]), .QN(n158) );
  DFFX1_LVT ex_reg_inst_reg_16_ ( .D(io_fpu_inst[16]), .CLK(n4097), .Q(
        n_T_648[4]), .QN(n157) );
  DFFX1_LVT ex_reg_inst_reg_15_ ( .D(io_fpu_inst[15]), .CLK(n4097), .Q(
        n_T_648[3]), .QN(n156) );
  DFFX1_LVT ex_reg_inst_reg_14_ ( .D(n9445), .CLK(n4097), .Q(
        io_dmem_req_bits_signed), .QN(n_T_648[2]) );
  DFFX1_LVT ex_reg_inst_reg_13_ ( .D(n9446), .CLK(n4097), .Q(n155), .QN(
        n_T_648[1]) );
  DFFX1_LVT ex_reg_inst_reg_12_ ( .D(n3583), .CLK(n4097), .Q(n154), .QN(
        n_T_648[0]) );
  DFFX1_LVT ex_reg_inst_reg_11_ ( .D(io_fpu_inst[11]), .CLK(n4097), .Q(
        io_dmem_req_bits_tag[5]), .QN(n588) );
  DFFX1_LVT ex_reg_inst_reg_10_ ( .D(n9447), .CLK(n4097), .Q(n589), .QN(
        io_dmem_req_bits_tag[4]) );
  DFFX1_LVT ex_reg_inst_reg_9_ ( .D(io_fpu_inst[9]), .CLK(n4097), .Q(
        io_dmem_req_bits_tag[3]), .QN(n590) );
  DFFX1_LVT ex_reg_inst_reg_8_ ( .D(io_fpu_inst[8]), .CLK(n4096), .Q(
        io_dmem_req_bits_tag[2]), .QN(n591) );
  DFFX1_LVT ex_reg_inst_reg_7_ ( .D(io_fpu_inst[7]), .CLK(n4096), .Q(
        io_dmem_req_bits_tag[1]), .QN(n592) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_0_ ( .D(
        ibuf_io_btb_resp_bht_history[0]), .CLK(n4096), .QN(n152) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_1_ ( .D(
        ibuf_io_btb_resp_bht_history[1]), .CLK(n4096), .QN(n151) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_2_ ( .D(
        ibuf_io_btb_resp_bht_history[2]), .CLK(n4096), .QN(n150) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_3_ ( .D(
        ibuf_io_btb_resp_bht_history[3]), .CLK(n4096), .QN(n149) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_4_ ( .D(
        ibuf_io_btb_resp_bht_history[4]), .CLK(n4096), .QN(n148) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_5_ ( .D(
        ibuf_io_btb_resp_bht_history[5]), .CLK(n4096), .QN(n147) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_6_ ( .D(
        ibuf_io_btb_resp_bht_history[6]), .CLK(n4096), .QN(n146) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_7_ ( .D(
        ibuf_io_btb_resp_bht_history[7]), .CLK(n4096), .QN(n145) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_0_ ( .D(ibuf_io_btb_resp_entry[0]), 
        .CLK(n4096), .QN(n144) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_1_ ( .D(ibuf_io_btb_resp_entry[1]), 
        .CLK(n4096), .QN(n143) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_2_ ( .D(ibuf_io_btb_resp_entry[2]), 
        .CLK(n4095), .QN(n142) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_3_ ( .D(ibuf_io_btb_resp_entry[3]), 
        .CLK(n4095), .QN(n141) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_4_ ( .D(ibuf_io_btb_resp_entry[4]), 
        .CLK(n4095), .QN(n140) );
  DFFX1_LVT ex_reg_pc_reg_0_ ( .D(ibuf_io_pc[0]), .CLK(n4095), .Q(n_T_698[0]), 
        .QN(n139) );
  DFFX1_LVT ex_reg_pc_reg_1_ ( .D(ibuf_io_pc[1]), .CLK(n4095), .Q(n_T_698[1]), 
        .QN(n138) );
  DFFX1_LVT ex_reg_pc_reg_2_ ( .D(ibuf_io_pc[2]), .CLK(n4095), .Q(n_T_698[2]), 
        .QN(n137) );
  DFFX1_LVT ex_reg_pc_reg_3_ ( .D(ibuf_io_pc[3]), .CLK(n4095), .Q(n_T_698[3]), 
        .QN(n136) );
  DFFX1_LVT ex_reg_pc_reg_4_ ( .D(ibuf_io_pc[4]), .CLK(n4095), .Q(n_T_698[4]), 
        .QN(n135) );
  DFFX1_LVT ex_reg_pc_reg_5_ ( .D(ibuf_io_pc[5]), .CLK(n4095), .Q(n_T_698[5]), 
        .QN(n134) );
  DFFX1_LVT ex_reg_pc_reg_6_ ( .D(ibuf_io_pc[6]), .CLK(n4095), .Q(n_T_698[6]), 
        .QN(n133) );
  DFFX1_LVT ex_reg_pc_reg_7_ ( .D(ibuf_io_pc[7]), .CLK(n4095), .Q(n_T_698[7]), 
        .QN(n132) );
  DFFX1_LVT ex_reg_pc_reg_8_ ( .D(ibuf_io_pc[8]), .CLK(n4095), .Q(n_T_698[8]), 
        .QN(n131) );
  DFFX1_LVT ex_reg_pc_reg_9_ ( .D(ibuf_io_pc[9]), .CLK(n4094), .Q(n_T_698[9]), 
        .QN(n130) );
  DFFX1_LVT ex_reg_pc_reg_10_ ( .D(ibuf_io_pc[10]), .CLK(n4094), .Q(
        n_T_698[10]), .QN(n129) );
  DFFX1_LVT ex_reg_pc_reg_11_ ( .D(ibuf_io_pc[11]), .CLK(n4094), .Q(
        n_T_698[11]), .QN(n128) );
  DFFX1_LVT ex_reg_pc_reg_12_ ( .D(ibuf_io_pc[12]), .CLK(n4094), .Q(
        n_T_698[12]), .QN(n127) );
  DFFX1_LVT ex_reg_pc_reg_13_ ( .D(ibuf_io_pc[13]), .CLK(n4094), .Q(
        n_T_698[13]), .QN(n126) );
  DFFX1_LVT ex_reg_pc_reg_14_ ( .D(ibuf_io_pc[14]), .CLK(n4094), .Q(
        n_T_698[14]), .QN(n125) );
  DFFX1_LVT ex_reg_pc_reg_15_ ( .D(ibuf_io_pc[15]), .CLK(n4094), .Q(
        n_T_698[15]), .QN(n124) );
  DFFX1_LVT ex_reg_pc_reg_16_ ( .D(ibuf_io_pc[16]), .CLK(n4094), .Q(
        n_T_698[16]), .QN(n123) );
  DFFX1_LVT ex_reg_pc_reg_17_ ( .D(ibuf_io_pc[17]), .CLK(n4094), .Q(
        n_T_698[17]), .QN(n122) );
  DFFX1_LVT ex_reg_pc_reg_18_ ( .D(ibuf_io_pc[18]), .CLK(n4094), .Q(
        n_T_698[18]), .QN(n121) );
  DFFX1_LVT ex_reg_pc_reg_19_ ( .D(ibuf_io_pc[19]), .CLK(n4094), .Q(
        n_T_698[19]), .QN(n120) );
  DFFX1_LVT ex_reg_pc_reg_20_ ( .D(ibuf_io_pc[20]), .CLK(n4094), .Q(
        n_T_698[20]), .QN(n119) );
  DFFX1_LVT ex_reg_pc_reg_21_ ( .D(ibuf_io_pc[21]), .CLK(n4093), .Q(
        n_T_698[21]), .QN(n118) );
  DFFX1_LVT ex_reg_pc_reg_22_ ( .D(ibuf_io_pc[22]), .CLK(n4093), .Q(
        n_T_698[22]), .QN(n117) );
  DFFX1_LVT ex_reg_pc_reg_23_ ( .D(ibuf_io_pc[23]), .CLK(n4093), .Q(
        n_T_698[23]), .QN(n116) );
  DFFX1_LVT ex_reg_pc_reg_24_ ( .D(ibuf_io_pc[24]), .CLK(n4093), .Q(
        n_T_698[24]), .QN(n115) );
  DFFX1_LVT ex_reg_pc_reg_25_ ( .D(ibuf_io_pc[25]), .CLK(n4093), .Q(
        n_T_698[25]), .QN(n114) );
  DFFX1_LVT ex_reg_pc_reg_26_ ( .D(ibuf_io_pc[26]), .CLK(n4093), .Q(
        n_T_698[26]), .QN(n113) );
  DFFX1_LVT ex_reg_pc_reg_27_ ( .D(ibuf_io_pc[27]), .CLK(n4093), .Q(
        n_T_698[27]), .QN(n112) );
  DFFX1_LVT ex_reg_pc_reg_28_ ( .D(ibuf_io_pc[28]), .CLK(n4093), .Q(
        n_T_698[28]), .QN(n111) );
  DFFX1_LVT ex_reg_pc_reg_29_ ( .D(ibuf_io_pc[29]), .CLK(n4093), .Q(
        n_T_698[29]), .QN(n110) );
  DFFX1_LVT ex_reg_pc_reg_30_ ( .D(ibuf_io_pc[30]), .CLK(n4093), .Q(
        n_T_698[30]), .QN(n109) );
  DFFX1_LVT ex_reg_pc_reg_31_ ( .D(ibuf_io_pc[31]), .CLK(n4093), .Q(
        n_T_698[31]), .QN(n108) );
  DFFX1_LVT ex_reg_pc_reg_32_ ( .D(ibuf_io_pc[32]), .CLK(n4093), .Q(
        n_T_698[32]), .QN(n107) );
  DFFX1_LVT ex_reg_pc_reg_33_ ( .D(ibuf_io_pc[33]), .CLK(n4092), .Q(
        n_T_698[33]), .QN(n106) );
  DFFX1_LVT ex_reg_pc_reg_34_ ( .D(ibuf_io_pc[34]), .CLK(n4092), .Q(
        n_T_698[34]), .QN(n105) );
  DFFX1_LVT ex_reg_pc_reg_35_ ( .D(ibuf_io_pc[35]), .CLK(n4092), .Q(
        n_T_698[35]), .QN(n104) );
  DFFX1_LVT ex_reg_pc_reg_36_ ( .D(ibuf_io_pc[36]), .CLK(n4092), .Q(
        n_T_698[36]), .QN(n103) );
  DFFX1_LVT ex_reg_pc_reg_37_ ( .D(ibuf_io_pc[37]), .CLK(n4092), .Q(
        n_T_698[37]), .QN(n102) );
  DFFX1_LVT ex_reg_pc_reg_38_ ( .D(ibuf_io_pc[38]), .CLK(n4092), .Q(
        n_T_698[38]), .QN(n101) );
  DFFX1_LVT ex_reg_pc_reg_39_ ( .D(ibuf_io_pc[39]), .CLK(n4092), .Q(
        n_T_698[39]), .QN(n100) );
  DFFSSRX1_LVT ex_reg_replay_reg ( .D(n9433), .SETB(n9417), .RSTB(1'b1), .CLK(
        n3594), .Q(n3233), .QN(ex_reg_replay) );
  DFFSSRX1_LVT ex_reg_xcpt_interrupt_reg ( .D(n9448), .SETB(n9417), .RSTB(1'b1), .CLK(n3594), .Q(n98), .QN(ex_reg_xcpt_interrupt) );
  DFFX1_LVT mem_ctrl_branch_reg ( .D(n323), .CLK(n4286), .QN(
        io_imem_bht_update_bits_branch) );
  DFFX1_LVT mem_ctrl_fp_reg ( .D(n322), .CLK(n4286), .Q(n3246), .QN(n2492) );
  DFFX1_LVT mem_ctrl_jalr_reg ( .D(ex_ctrl_jalr), .CLK(n4286), .Q(
        mem_ctrl_jalr), .QN(n3104) );
  DFFX1_LVT mem_reg_wdata_reg_62_ ( .D(alu_io_out[62]), .CLK(n4286), .Q(
        n_T_918[62]) );
  DFFX1_LVT mem_reg_wdata_reg_61_ ( .D(alu_io_out[61]), .CLK(n4286), .Q(
        n_T_918[61]) );
  DFFX1_LVT mem_reg_wdata_reg_60_ ( .D(alu_io_out[60]), .CLK(n4286), .Q(
        n_T_918[60]) );
  DFFX1_LVT mem_reg_wdata_reg_59_ ( .D(alu_io_out[59]), .CLK(n4287), .Q(
        n_T_918[59]) );
  DFFX1_LVT mem_reg_wdata_reg_58_ ( .D(alu_io_out[58]), .CLK(n4287), .Q(
        n_T_918[58]) );
  DFFX1_LVT mem_reg_wdata_reg_57_ ( .D(alu_io_out[57]), .CLK(n4287), .Q(
        n_T_918[57]) );
  DFFX1_LVT mem_reg_wdata_reg_56_ ( .D(alu_io_out[56]), .CLK(n4287), .Q(
        n_T_918[56]) );
  DFFX1_LVT mem_reg_wdata_reg_55_ ( .D(alu_io_out[55]), .CLK(n4287), .Q(
        n_T_918[55]) );
  DFFX1_LVT mem_reg_wdata_reg_54_ ( .D(alu_io_out[54]), .CLK(n4287), .Q(
        n_T_918[54]) );
  DFFX1_LVT mem_reg_wdata_reg_53_ ( .D(alu_io_out[53]), .CLK(n4287), .Q(
        n_T_918[53]) );
  DFFX1_LVT mem_reg_wdata_reg_52_ ( .D(alu_io_out[52]), .CLK(n4287), .Q(
        n_T_918[52]) );
  DFFX1_LVT mem_reg_wdata_reg_51_ ( .D(alu_io_out[51]), .CLK(n4288), .Q(
        n_T_918[51]), .QN(n3249) );
  DFFX1_LVT mem_reg_wdata_reg_50_ ( .D(alu_io_out[50]), .CLK(n4287), .Q(
        n_T_918[50]) );
  DFFX1_LVT mem_reg_wdata_reg_49_ ( .D(alu_io_out[49]), .CLK(n4287), .Q(
        n_T_918[49]) );
  DFFX1_LVT mem_reg_wdata_reg_48_ ( .D(alu_io_out[48]), .CLK(n4287), .Q(
        n_T_918[48]) );
  DFFX1_LVT mem_reg_wdata_reg_47_ ( .D(alu_io_out[47]), .CLK(n4288), .Q(
        n_T_918[47]) );
  DFFX1_LVT mem_reg_wdata_reg_46_ ( .D(alu_io_out[46]), .CLK(n4287), .Q(
        n_T_918[46]) );
  DFFX1_LVT mem_reg_wdata_reg_45_ ( .D(alu_io_out[45]), .CLK(n4288), .Q(
        n_T_918[45]) );
  DFFX1_LVT mem_reg_wdata_reg_44_ ( .D(alu_io_out[44]), .CLK(n4288), .Q(
        n_T_918[44]) );
  DFFX1_LVT mem_reg_wdata_reg_43_ ( .D(alu_io_out[43]), .CLK(n4288), .Q(
        n_T_918[43]) );
  DFFX1_LVT mem_reg_wdata_reg_42_ ( .D(alu_io_out[42]), .CLK(n4288), .Q(
        n_T_918[42]) );
  DFFX1_LVT mem_reg_wdata_reg_41_ ( .D(alu_io_out[41]), .CLK(n4288), .Q(
        n_T_918[41]) );
  DFFX1_LVT mem_reg_wdata_reg_40_ ( .D(alu_io_out[40]), .CLK(n4288), .Q(
        n_T_918[40]) );
  DFFX1_LVT mem_reg_wdata_reg_39_ ( .D(alu_io_out[39]), .CLK(n4288), .Q(
        n_T_918[39]) );
  DFFX1_LVT mem_reg_wdata_reg_38_ ( .D(alu_io_out[38]), .CLK(n4288), .Q(
        n_T_918[38]), .QN(n3205) );
  DFFX1_LVT mem_reg_wdata_reg_37_ ( .D(alu_io_out[37]), .CLK(n4289), .Q(
        n_T_918[37]), .QN(n3528) );
  DFFX1_LVT mem_reg_wdata_reg_36_ ( .D(alu_io_out[36]), .CLK(n4288), .Q(
        n_T_918[36]), .QN(n3227) );
  DFFX1_LVT mem_reg_wdata_reg_35_ ( .D(alu_io_out[35]), .CLK(n4289), .Q(
        n_T_918[35]) );
  DFFX1_LVT mem_reg_wdata_reg_34_ ( .D(alu_io_out[34]), .CLK(n4288), .Q(
        n_T_918[34]) );
  DFFX1_LVT mem_reg_wdata_reg_33_ ( .D(alu_io_out[33]), .CLK(n4289), .Q(
        n_T_918[33]), .QN(n3210) );
  DFFX1_LVT mem_reg_wdata_reg_32_ ( .D(alu_io_out[32]), .CLK(n4289), .Q(
        n_T_918[32]), .QN(n3226) );
  DFFX1_LVT mem_reg_wdata_reg_31_ ( .D(alu_io_out[31]), .CLK(n4289), .Q(
        n_T_918[31]), .QN(n3105) );
  DFFX1_LVT mem_reg_wdata_reg_30_ ( .D(alu_io_out[30]), .CLK(n4290), .Q(
        n_T_918[30]), .QN(n3219) );
  DFFX1_LVT mem_reg_wdata_reg_29_ ( .D(alu_io_out[29]), .CLK(n4289), .Q(
        n_T_918[29]), .QN(n3111) );
  DFFX1_LVT mem_reg_wdata_reg_28_ ( .D(alu_io_out[28]), .CLK(n4289), .Q(
        n_T_918[28]) );
  DFFX1_LVT mem_reg_wdata_reg_27_ ( .D(alu_io_out[27]), .CLK(n4289), .Q(
        n_T_918[27]), .QN(n3209) );
  DFFX1_LVT mem_reg_wdata_reg_26_ ( .D(alu_io_out[26]), .CLK(n4289), .Q(
        n_T_918[26]), .QN(n3218) );
  DFFX1_LVT mem_reg_wdata_reg_25_ ( .D(alu_io_out[25]), .CLK(n4289), .Q(
        n_T_918[25]), .QN(n3110) );
  DFFX1_LVT mem_reg_wdata_reg_24_ ( .D(alu_io_out[24]), .CLK(n4289), .Q(
        n_T_918[24]) );
  DFFX1_LVT mem_reg_wdata_reg_23_ ( .D(alu_io_out[23]), .CLK(n4290), .Q(
        n_T_918[23]), .QN(n3213) );
  DFFX1_LVT mem_reg_wdata_reg_22_ ( .D(alu_io_out[22]), .CLK(n4289), .Q(
        n_T_918[22]), .QN(n3216) );
  DFFX1_LVT mem_reg_wdata_reg_21_ ( .D(alu_io_out[21]), .CLK(n4290), .Q(
        n_T_918[21]) );
  DFFX1_LVT mem_reg_wdata_reg_20_ ( .D(alu_io_out[20]), .CLK(n4290), .Q(
        n_T_918[20]), .QN(n3224) );
  DFFX1_LVT mem_reg_wdata_reg_19_ ( .D(alu_io_out[19]), .CLK(n4290), .Q(
        n_T_918[19]), .QN(n3212) );
  DFFX1_LVT mem_reg_wdata_reg_18_ ( .D(alu_io_out[18]), .CLK(n4290), .Q(
        n_T_918[18]), .QN(n3220) );
  DFFX1_LVT mem_reg_wdata_reg_17_ ( .D(alu_io_out[17]), .CLK(n4290), .Q(
        n_T_918[17]), .QN(n3107) );
  DFFX1_LVT mem_reg_wdata_reg_16_ ( .D(alu_io_out[16]), .CLK(n4291), .Q(
        n_T_918[16]) );
  DFFX1_LVT mem_reg_wdata_reg_15_ ( .D(alu_io_out[15]), .CLK(n4290), .Q(
        n_T_918[15]) );
  DFFX1_LVT mem_reg_wdata_reg_14_ ( .D(alu_io_out[14]), .CLK(n4290), .Q(
        n_T_918[14]), .QN(n3223) );
  DFFX1_LVT mem_reg_wdata_reg_13_ ( .D(alu_io_out[13]), .CLK(n4290), .Q(
        n_T_918[13]), .QN(n3106) );
  DFFX1_LVT mem_reg_wdata_reg_12_ ( .D(alu_io_out[12]), .CLK(n4290), .Q(
        n_T_918[12]), .QN(n3221) );
  DFFX1_LVT mem_reg_wdata_reg_11_ ( .D(alu_io_out[11]), .CLK(n4291), .Q(
        n_T_918[11]), .QN(n3211) );
  DFFX1_LVT mem_reg_wdata_reg_10_ ( .D(alu_io_out[10]), .CLK(n4290), .Q(
        n_T_918[10]), .QN(n3225) );
  DFFX1_LVT mem_reg_wdata_reg_9_ ( .D(alu_io_out[9]), .CLK(n4291), .Q(
        n_T_918[9]), .QN(n3108) );
  DFFX1_LVT mem_reg_wdata_reg_8_ ( .D(alu_io_out[8]), .CLK(n4291), .Q(
        n_T_918[8]), .QN(n3222) );
  DFFX1_LVT mem_reg_wdata_reg_7_ ( .D(alu_io_out[7]), .CLK(n4291), .Q(
        n_T_918[7]), .QN(n3214) );
  DFFX1_LVT mem_reg_wdata_reg_6_ ( .D(alu_io_out[6]), .CLK(n4291), .Q(
        n_T_918[6]), .QN(n3217) );
  DFFX1_LVT mem_reg_wdata_reg_5_ ( .D(alu_io_out[5]), .CLK(n4291), .Q(
        n_T_918[5]), .QN(n3109) );
  DFFX1_LVT mem_reg_wdata_reg_4_ ( .D(alu_io_out[4]), .CLK(n4291), .Q(
        n_T_918[4]), .QN(n3112) );
  DFFX1_LVT mem_reg_wdata_reg_3_ ( .D(alu_io_out[3]), .CLK(n4291), .Q(
        n_T_918[3]), .QN(n3208) );
  DFFX1_LVT mem_reg_wdata_reg_2_ ( .D(alu_io_out[2]), .CLK(n4292), .Q(
        n_T_918[2]) );
  DFFX1_LVT mem_reg_wdata_reg_1_ ( .D(alu_io_out[1]), .CLK(n4291), .Q(
        n_T_918[1]), .QN(n3207) );
  DFFX1_LVT mem_reg_wdata_reg_0_ ( .D(alu_io_out[0]), .CLK(n4291), .Q(
        n_T_918[0]) );
  DFFX1_LVT ex_reg_cause_reg_0_ ( .D(N303), .CLK(n4092), .QN(n80) );
  DFFX1_LVT ex_ctrl_sel_alu2_reg_1_ ( .D(N275), .CLK(n4313), .Q(
        ex_ctrl_sel_alu2[1]), .QN(n3278) );
  DFFX1_LVT ex_ctrl_sel_alu1_reg_0_ ( .D(N279), .CLK(n4313), .Q(
        ex_ctrl_sel_alu1_0_) );
  DFFSSRX1_LVT ex_ctrl_alu_fn_reg_0_ ( .D(n3583), .SETB(n1589), .RSTB(1'b1), 
        .CLK(n4312), .QN(alu_io_fn[0]) );
  DFFX1_LVT ex_ctrl_alu_fn_reg_1_ ( .D(N282), .CLK(n4313), .Q(alu_io_fn[1]) );
  DFFX1_LVT ex_ctrl_alu_fn_reg_3_ ( .D(N284), .CLK(n4313), .Q(alu_io_fn[3]) );
  DFFX1_LVT ex_ctrl_alu_dw_reg ( .D(n_GEN_9), .CLK(n4313), .Q(alu_io_dw) );
  DFFX1_LVT ex_ctrl_sel_alu2_reg_0_ ( .D(N274), .CLK(n4313), .Q(
        ex_ctrl_sel_alu2[0]) );
  DFFX1_LVT ex_reg_cause_reg_1_ ( .D(N304), .CLK(n4092), .QN(n76) );
  DFFSSRX1_LVT ex_reg_cause_reg_2_ ( .D(n9448), .SETB(
        csr_io_interrupt_cause[2]), .RSTB(n74), .CLK(n4092), .Q(n73) );
  DFFX1_LVT mem_reg_mem_size_reg_1_ ( .D(n586), .CLK(n4292), .Q(n72) );
  DFFX1_LVT mem_reg_mem_size_reg_0_ ( .D(n313), .CLK(n4291), .Q(n71) );
  DFFX1_LVT mem_ctrl_jal_reg ( .D(ex_ctrl_jal), .CLK(n4292), .Q(n3230), .QN(
        n555) );
  DFFX1_LVT mem_reg_rvc_reg ( .D(ex_reg_rvc), .CLK(n4292), .Q(mem_reg_rvc), 
        .QN(n570) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_4_ ( .D(n140), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[4]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_3_ ( .D(n141), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[3]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_2_ ( .D(n142), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[2]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_1_ ( .D(n143), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[1]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_0_ ( .D(n144), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[0]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_7_ ( .D(n145), .CLK(n4292), .QN(
        io_imem_bht_update_bits_prediction_history[7]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_6_ ( .D(n146), .CLK(n4292), .QN(
        io_imem_bht_update_bits_prediction_history[6]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_5_ ( .D(n147), .CLK(n4292), .QN(
        io_imem_bht_update_bits_prediction_history[5]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_4_ ( .D(n148), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[4]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_3_ ( .D(n149), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[3]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_2_ ( .D(n150), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[2]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_1_ ( .D(n151), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[1]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_0_ ( .D(n152), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[0]) );
  DFFSSRX1_LVT mem_reg_load_reg ( .D(n312), .SETB(n997), .RSTB(n882), .CLK(
        n4286), .QN(mem_reg_load) );
  DFFSSRX1_LVT mem_reg_store_reg ( .D(n312), .SETB(n997), .RSTB(n996), .CLK(
        n4286), .QN(mem_reg_store) );
  DFFX1_LVT mem_ctrl_mem_reg ( .D(n312), .CLK(n4293), .Q(n572), .QN(
        mem_ctrl_mem) );
  DFFX1_LVT mem_br_taken_reg ( .D(alu_io_cmp_out), .CLK(n4293), .Q(
        io_imem_bht_update_bits_taken), .QN(n3310) );
  DFFX1_LVT mem_ctrl_wfd_reg ( .D(n315), .CLK(n4293), .Q(n69), .QN(
        mem_ctrl_wfd) );
  DFFX1_LVT mem_ctrl_div_reg ( .D(n317), .CLK(n4293), .Q(n370) );
  DFFX1_LVT mem_ctrl_wxd_reg ( .D(n314), .CLK(n4293), .QN(mem_ctrl_wxd) );
  DFFX1_LVT mem_ctrl_csr_reg_2_ ( .D(n310), .CLK(n4293), .Q(n68), .QN(
        mem_ctrl_csr[2]) );
  DFFX1_LVT mem_ctrl_csr_reg_1_ ( .D(n319), .CLK(n4294), .Q(n369), .QN(n3279)
         );
  DFFX1_LVT mem_ctrl_csr_reg_0_ ( .D(n320), .CLK(n4294), .Q(n67), .QN(
        mem_ctrl_csr[0]) );
  DFFSSRX1_LVT mem_ctrl_fence_i_reg ( .D(n9516), .SETB(ex_ctrl_jalr), .RSTB(
        n318), .CLK(n4286), .Q(n66) );
  DFFX1_LVT mem_reg_cause_reg_3_ ( .D(n75), .CLK(n4294), .QN(mem_reg_cause[3])
         );
  DFFX1_LVT mem_reg_cause_reg_2_ ( .D(n73), .CLK(n4294), .QN(mem_reg_cause[2])
         );
  DFFX1_LVT mem_reg_cause_reg_1_ ( .D(n76), .CLK(n4294), .Q(n63) );
  DFFX1_LVT mem_reg_cause_reg_0_ ( .D(n80), .CLK(n4294), .QN(mem_reg_cause[0])
         );
  DFFX1_LVT mem_reg_pc_reg_39_ ( .D(n100), .CLK(n4294), .Q(n62), .QN(
        mem_reg_pc[39]) );
  DFFX1_LVT mem_reg_pc_reg_38_ ( .D(n101), .CLK(n4294), .Q(n61), .QN(
        mem_reg_pc[38]) );
  DFFX1_LVT mem_reg_pc_reg_37_ ( .D(n102), .CLK(n4294), .Q(n60), .QN(
        mem_reg_pc[37]) );
  DFFX1_LVT mem_reg_pc_reg_36_ ( .D(n103), .CLK(n4294), .Q(n59), .QN(
        mem_reg_pc[36]) );
  DFFX1_LVT mem_reg_pc_reg_35_ ( .D(n104), .CLK(n4295), .Q(n58), .QN(
        mem_reg_pc[35]) );
  DFFX1_LVT mem_reg_pc_reg_34_ ( .D(n105), .CLK(n4295), .Q(n57), .QN(
        mem_reg_pc[34]) );
  DFFX1_LVT mem_reg_pc_reg_33_ ( .D(n106), .CLK(n4295), .Q(n56), .QN(
        mem_reg_pc[33]) );
  DFFX1_LVT mem_reg_pc_reg_32_ ( .D(n107), .CLK(n4295), .Q(n55), .QN(
        mem_reg_pc[32]) );
  DFFX1_LVT mem_reg_pc_reg_31_ ( .D(n108), .CLK(n4295), .Q(n54), .QN(
        mem_reg_pc[31]) );
  DFFX1_LVT mem_reg_pc_reg_30_ ( .D(n109), .CLK(n4295), .Q(n53), .QN(
        mem_reg_pc[30]) );
  DFFX1_LVT mem_reg_pc_reg_29_ ( .D(n110), .CLK(n4295), .Q(n52), .QN(
        mem_reg_pc[29]) );
  DFFX1_LVT mem_reg_pc_reg_28_ ( .D(n111), .CLK(n4295), .Q(n51), .QN(
        mem_reg_pc[28]) );
  DFFX1_LVT mem_reg_pc_reg_27_ ( .D(n112), .CLK(n4295), .Q(n50), .QN(
        mem_reg_pc[27]) );
  DFFX1_LVT mem_reg_pc_reg_26_ ( .D(n113), .CLK(n4295), .Q(n49), .QN(
        mem_reg_pc[26]) );
  DFFX1_LVT mem_reg_pc_reg_25_ ( .D(n114), .CLK(n4295), .Q(n48), .QN(
        mem_reg_pc[25]) );
  DFFX1_LVT mem_reg_pc_reg_24_ ( .D(n115), .CLK(n4295), .Q(n47), .QN(
        mem_reg_pc[24]) );
  DFFX1_LVT mem_reg_pc_reg_23_ ( .D(n116), .CLK(n4296), .Q(n46), .QN(
        mem_reg_pc[23]) );
  DFFX1_LVT mem_reg_pc_reg_22_ ( .D(n117), .CLK(n4296), .Q(n45), .QN(
        mem_reg_pc[22]) );
  DFFX1_LVT mem_reg_pc_reg_21_ ( .D(n118), .CLK(n4296), .Q(n44), .QN(
        mem_reg_pc[21]) );
  DFFX1_LVT mem_reg_pc_reg_20_ ( .D(n119), .CLK(n4296), .Q(n43), .QN(
        mem_reg_pc[20]) );
  DFFX1_LVT mem_reg_pc_reg_19_ ( .D(n120), .CLK(n4296), .Q(n42), .QN(
        mem_reg_pc[19]) );
  DFFX1_LVT mem_reg_pc_reg_18_ ( .D(n121), .CLK(n4296), .Q(n41), .QN(
        mem_reg_pc[18]) );
  DFFX1_LVT mem_reg_pc_reg_17_ ( .D(n122), .CLK(n4296), .Q(n40), .QN(
        mem_reg_pc[17]) );
  DFFX1_LVT mem_reg_pc_reg_16_ ( .D(n123), .CLK(n4296), .Q(n39), .QN(
        mem_reg_pc[16]) );
  DFFX1_LVT mem_reg_pc_reg_15_ ( .D(n124), .CLK(n4296), .Q(n38), .QN(
        mem_reg_pc[15]) );
  DFFX1_LVT mem_reg_pc_reg_14_ ( .D(n125), .CLK(n4296), .Q(n37), .QN(
        mem_reg_pc[14]) );
  DFFX1_LVT mem_reg_pc_reg_13_ ( .D(n126), .CLK(n4296), .Q(n36), .QN(
        mem_reg_pc[13]) );
  DFFX1_LVT mem_reg_pc_reg_12_ ( .D(n127), .CLK(n4296), .Q(n35), .QN(
        mem_reg_pc[12]) );
  DFFX1_LVT mem_reg_pc_reg_11_ ( .D(n128), .CLK(n4297), .Q(n34), .QN(
        mem_reg_pc[11]) );
  DFFX1_LVT mem_reg_pc_reg_10_ ( .D(n129), .CLK(n4297), .Q(n33), .QN(
        mem_reg_pc[10]) );
  DFFX1_LVT mem_reg_pc_reg_9_ ( .D(n130), .CLK(n4297), .Q(n32), .QN(
        mem_reg_pc[9]) );
  DFFX1_LVT mem_reg_pc_reg_8_ ( .D(n131), .CLK(n4297), .Q(n31), .QN(
        mem_reg_pc[8]) );
  DFFX1_LVT mem_reg_pc_reg_7_ ( .D(n132), .CLK(n4297), .Q(n30), .QN(
        mem_reg_pc[7]) );
  DFFX1_LVT mem_reg_pc_reg_6_ ( .D(n133), .CLK(n4297), .Q(n29), .QN(
        mem_reg_pc[6]) );
  DFFX1_LVT mem_reg_pc_reg_5_ ( .D(n134), .CLK(n4297), .Q(n28), .QN(
        mem_reg_pc[5]) );
  DFFX1_LVT mem_reg_pc_reg_4_ ( .D(n135), .CLK(n4297), .Q(n27), .QN(
        mem_reg_pc[4]) );
  DFFX1_LVT mem_reg_pc_reg_3_ ( .D(n136), .CLK(n4297), .Q(n26), .QN(
        mem_reg_pc[3]) );
  DFFX1_LVT mem_reg_pc_reg_2_ ( .D(n137), .CLK(n4297), .Q(n25), .QN(
        mem_reg_pc[2]) );
  DFFX1_LVT mem_reg_pc_reg_1_ ( .D(n138), .CLK(n4297), .Q(n24), .QN(
        mem_reg_pc[1]) );
  DFFX1_LVT mem_reg_pc_reg_0_ ( .D(n139), .CLK(n4297), .Q(n23), .QN(
        io_imem_btb_update_bits_br_pc[0]) );
  DFFX1_LVT mem_reg_inst_reg_31_ ( .D(n172), .CLK(n4298), .Q(n22), .QN(
        n_T_844_10_) );
  DFFX1_LVT mem_reg_inst_reg_30_ ( .D(n171), .CLK(n4298), .Q(n21), .QN(
        n_T_849[10]) );
  DFFX1_LVT mem_reg_inst_reg_29_ ( .D(n170), .CLK(n4298), .Q(n20), .QN(
        n_T_849[9]) );
  DFFX1_LVT mem_reg_inst_reg_28_ ( .D(n169), .CLK(n4298), .Q(n19), .QN(
        n_T_849[8]) );
  DFFX1_LVT mem_reg_inst_reg_27_ ( .D(n168), .CLK(n4298), .Q(n18), .QN(
        n_T_849[7]) );
  DFFX1_LVT mem_reg_inst_reg_26_ ( .D(n167), .CLK(n4298), .Q(n17), .QN(
        n_T_849[6]) );
  DFFX1_LVT mem_reg_inst_reg_25_ ( .D(n166), .CLK(n4298), .Q(n16), .QN(
        n_T_849[5]) );
  DFFX1_LVT mem_reg_inst_reg_24_ ( .D(n165), .CLK(n4298), .Q(n15), .QN(
        n_T_911[4]) );
  DFFX1_LVT mem_reg_inst_reg_23_ ( .D(n164), .CLK(n4298), .Q(n14), .QN(
        n_T_911[3]) );
  DFFX1_LVT mem_reg_inst_reg_22_ ( .D(n163), .CLK(n4298), .Q(n13), .QN(
        n_T_911[2]) );
  DFFX1_LVT mem_reg_inst_reg_21_ ( .D(n162), .CLK(n4298), .Q(n12), .QN(
        n_T_911[1]) );
  DFFX1_LVT mem_reg_inst_reg_20_ ( .D(n161), .CLK(n4298), .Q(n11), .QN(
        n_T_911_11) );
  DFFX1_LVT mem_reg_inst_reg_19_ ( .D(n160), .CLK(n4299), .QN(n_T_904[7]) );
  DFFX1_LVT mem_reg_inst_reg_18_ ( .D(n159), .CLK(n4299), .QN(n_T_904[6]) );
  DFFX1_LVT mem_reg_inst_reg_17_ ( .D(n158), .CLK(n4299), .QN(n_T_904[5]) );
  DFFX1_LVT mem_reg_inst_reg_16_ ( .D(n157), .CLK(n4299), .QN(n_T_904[4]) );
  DFFX1_LVT mem_reg_inst_reg_15_ ( .D(n156), .CLK(n4299), .QN(n_T_904[3]) );
  DFFX1_LVT mem_reg_inst_reg_14_ ( .D(io_dmem_req_bits_signed), .CLK(n4299), 
        .QN(n_T_904[2]) );
  DFFX1_LVT mem_reg_inst_reg_13_ ( .D(n155), .CLK(n4299), .QN(n_T_904[1]) );
  DFFX1_LVT mem_reg_inst_reg_12_ ( .D(n154), .CLK(n4299), .QN(n_T_904[0]) );
  DFFX1_LVT mem_reg_inst_reg_11_ ( .D(n588), .CLK(n4299), .Q(n595), .QN(
        n_T_849[4]) );
  DFFX1_LVT mem_reg_inst_reg_10_ ( .D(n589), .CLK(n4299), .Q(n596), .QN(n2566)
         );
  DFFX1_LVT mem_reg_inst_reg_9_ ( .D(n590), .CLK(n4299), .Q(n3200), .QN(
        n_T_849[2]) );
  DFFX1_LVT mem_reg_inst_reg_8_ ( .D(n591), .CLK(n4299), .Q(n598), .QN(
        n_T_849[1]) );
  DFFX1_LVT ex_reg_rs_bypass_1_reg ( .D(do_bypass_1), .CLK(n4313), .Q(
        ex_reg_rs_bypass_1), .QN(n3243) );
  DFFX1_LVT ex_reg_load_use_reg ( .D(n9424), .CLK(n4312), .Q(ex_reg_load_use)
         );
  DFFSSRX1_LVT mem_reg_xcpt_interrupt_reg ( .D(n98), .SETB(n9418), .RSTB(1'b1), 
        .CLK(n3594), .QN(mem_reg_xcpt_interrupt) );
  DFFX1_LVT wb_ctrl_wxd_reg ( .D(mem_ctrl_wxd), .CLK(n4300), .Q(wb_ctrl_wxd)
         );
  DFFX1_LVT wb_ctrl_csr_reg_2_ ( .D(n68), .CLK(n4300), .QN(wb_ctrl_csr[2]) );
  DFFX1_LVT wb_ctrl_csr_reg_1_ ( .D(n369), .CLK(n4300), .QN(wb_ctrl_csr[1]) );
  DFFX1_LVT wb_ctrl_csr_reg_0_ ( .D(n67), .CLK(n4300), .QN(wb_ctrl_csr[0]) );
  DFFX1_LVT wb_ctrl_wfd_reg ( .D(n69), .CLK(n4300), .Q(n3229), .QN(wb_ctrl_wfd) );
  DFFX1_LVT wb_ctrl_div_reg ( .D(n370), .CLK(n4300), .QN(wb_ctrl_div) );
  DFFX1_LVT wb_ctrl_mem_reg ( .D(n572), .CLK(n4300), .QN(wb_ctrl_mem) );
  DFFX1_LVT wb_reg_wdata_reg_63_ ( .D(N661), .CLK(n4300), .Q(n_T_1165[63]) );
  DFFX1_LVT wb_reg_wdata_reg_62_ ( .D(N660), .CLK(n4300), .Q(n_T_1165[62]) );
  DFFX1_LVT wb_reg_wdata_reg_61_ ( .D(N659), .CLK(n4300), .Q(n_T_1165[61]) );
  DFFX1_LVT wb_reg_wdata_reg_60_ ( .D(N658), .CLK(n4301), .Q(n_T_1165[60]) );
  DFFX1_LVT wb_reg_wdata_reg_59_ ( .D(N657), .CLK(n4301), .Q(n_T_1165[59]) );
  DFFX1_LVT wb_reg_wdata_reg_58_ ( .D(N656), .CLK(n4301), .Q(n_T_1165[58]) );
  DFFX1_LVT wb_reg_wdata_reg_57_ ( .D(N655), .CLK(n4301), .Q(n_T_1165[57]) );
  DFFX1_LVT wb_reg_wdata_reg_56_ ( .D(N654), .CLK(n4301), .Q(n_T_1165[56]) );
  DFFX1_LVT wb_reg_wdata_reg_55_ ( .D(N653), .CLK(n4301), .Q(n_T_1165[55]) );
  DFFX1_LVT wb_reg_wdata_reg_54_ ( .D(N652), .CLK(n4301), .Q(n_T_1165[54]) );
  DFFX1_LVT wb_reg_wdata_reg_53_ ( .D(N651), .CLK(n4301), .Q(n_T_1165[53]) );
  DFFX1_LVT wb_reg_wdata_reg_52_ ( .D(N650), .CLK(n4301), .Q(n_T_1165[52]) );
  DFFX1_LVT wb_reg_wdata_reg_51_ ( .D(N649), .CLK(n4301), .Q(n_T_1165[51]) );
  DFFX1_LVT wb_reg_wdata_reg_50_ ( .D(N648), .CLK(n4301), .Q(n_T_1165[50]) );
  DFFX1_LVT wb_reg_wdata_reg_49_ ( .D(N647), .CLK(n4301), .Q(n_T_1165[49]) );
  DFFX1_LVT wb_reg_wdata_reg_48_ ( .D(N646), .CLK(n4302), .Q(n_T_1165[48]) );
  DFFX1_LVT wb_reg_wdata_reg_47_ ( .D(N645), .CLK(n4302), .Q(n_T_1165[47]) );
  DFFX1_LVT wb_reg_wdata_reg_46_ ( .D(N644), .CLK(n4302), .Q(n_T_1165[46]) );
  DFFX1_LVT wb_reg_wdata_reg_45_ ( .D(N643), .CLK(n4302), .Q(n_T_1165[45]) );
  DFFX1_LVT wb_reg_wdata_reg_44_ ( .D(N642), .CLK(n4302), .Q(n_T_1165[44]) );
  DFFX1_LVT wb_reg_wdata_reg_43_ ( .D(N641), .CLK(n4302), .Q(n_T_1165[43]) );
  DFFX1_LVT wb_reg_wdata_reg_42_ ( .D(N640), .CLK(n4302), .Q(n_T_1165[42]) );
  DFFX1_LVT wb_reg_wdata_reg_41_ ( .D(N639), .CLK(n4302), .Q(n_T_1165[41]) );
  DFFX1_LVT wb_reg_wdata_reg_40_ ( .D(N638), .CLK(n4302), .Q(n_T_1165[40]) );
  DFFX1_LVT wb_reg_wdata_reg_39_ ( .D(N637), .CLK(n4302), .Q(n_T_1165[39]) );
  DFFX1_LVT wb_reg_wdata_reg_38_ ( .D(N636), .CLK(n4302), .Q(
        io_imem_sfence_bits_addr[38]), .QN(n3228) );
  DFFX1_LVT wb_reg_wdata_reg_37_ ( .D(N635), .CLK(n4302), .Q(
        io_imem_sfence_bits_addr[37]) );
  DFFX1_LVT wb_reg_wdata_reg_36_ ( .D(N634), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[36]) );
  DFFX1_LVT wb_reg_wdata_reg_35_ ( .D(N633), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[35]) );
  DFFX1_LVT wb_reg_wdata_reg_34_ ( .D(N632), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[34]) );
  DFFX1_LVT wb_reg_wdata_reg_33_ ( .D(N631), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[33]) );
  DFFX1_LVT wb_reg_wdata_reg_32_ ( .D(N630), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[32]) );
  DFFX1_LVT wb_reg_wdata_reg_31_ ( .D(N629), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[31]) );
  DFFX1_LVT wb_reg_wdata_reg_30_ ( .D(N628), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[30]) );
  DFFX1_LVT wb_reg_wdata_reg_29_ ( .D(N627), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[29]) );
  DFFX1_LVT wb_reg_wdata_reg_28_ ( .D(N626), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[28]) );
  DFFX1_LVT wb_reg_wdata_reg_27_ ( .D(N625), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[27]) );
  DFFX1_LVT wb_reg_wdata_reg_26_ ( .D(N624), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[26]) );
  DFFX1_LVT wb_reg_wdata_reg_25_ ( .D(N623), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[25]) );
  DFFX1_LVT wb_reg_wdata_reg_24_ ( .D(N622), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[24]) );
  DFFX1_LVT wb_reg_wdata_reg_23_ ( .D(N621), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[23]) );
  DFFX1_LVT wb_reg_wdata_reg_22_ ( .D(N620), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[22]) );
  DFFX1_LVT wb_reg_wdata_reg_21_ ( .D(N619), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[21]) );
  DFFX1_LVT wb_reg_wdata_reg_20_ ( .D(N618), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[20]) );
  DFFX1_LVT wb_reg_wdata_reg_19_ ( .D(N617), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[19]) );
  DFFX1_LVT wb_reg_wdata_reg_18_ ( .D(N616), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[18]) );
  DFFX1_LVT wb_reg_wdata_reg_17_ ( .D(N615), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[17]) );
  DFFX1_LVT wb_reg_wdata_reg_16_ ( .D(N614), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[16]) );
  DFFX1_LVT wb_reg_wdata_reg_15_ ( .D(N613), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[15]) );
  DFFX1_LVT wb_reg_wdata_reg_14_ ( .D(N612), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[14]) );
  DFFX1_LVT wb_reg_wdata_reg_13_ ( .D(N611), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[13]) );
  DFFX1_LVT wb_reg_wdata_reg_12_ ( .D(N610), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[12]) );
  DFFX1_LVT wb_reg_wdata_reg_11_ ( .D(N609), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[11]) );
  DFFX1_LVT wb_reg_wdata_reg_10_ ( .D(N608), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[10]) );
  DFFX1_LVT wb_reg_wdata_reg_9_ ( .D(N607), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[9]) );
  DFFX1_LVT wb_reg_wdata_reg_8_ ( .D(N606), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[8]) );
  DFFX1_LVT wb_reg_wdata_reg_7_ ( .D(N605), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[7]) );
  DFFX1_LVT wb_reg_wdata_reg_6_ ( .D(N604), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[6]) );
  DFFX1_LVT wb_reg_wdata_reg_5_ ( .D(N603), .CLK(n4300), .Q(
        io_imem_sfence_bits_addr[5]) );
  DFFX1_LVT wb_reg_wdata_reg_4_ ( .D(N602), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[4]) );
  DFFX1_LVT wb_reg_wdata_reg_3_ ( .D(N601), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[3]) );
  DFFX1_LVT wb_reg_wdata_reg_2_ ( .D(N600), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[2]) );
  DFFX1_LVT wb_reg_wdata_reg_1_ ( .D(N599), .CLK(n4306), .Q(
        io_imem_sfence_bits_addr[1]) );
  DFFX1_LVT wb_ctrl_fence_i_reg ( .D(n66), .CLK(n4306), .QN(wb_ctrl_fence_i)
         );
  DFFX1_LVT wb_reg_sfence_reg ( .D(n326), .CLK(n4306), .QN(wb_reg_sfence) );
  DFFX1_LVT wb_reg_pc_reg_39_ ( .D(n62), .CLK(n4306), .QN(csr_io_pc[39]) );
  DFFX1_LVT wb_reg_pc_reg_38_ ( .D(n61), .CLK(n4306), .QN(csr_io_pc[38]) );
  DFFX1_LVT wb_reg_pc_reg_37_ ( .D(n60), .CLK(n4306), .QN(csr_io_pc[37]) );
  DFFX1_LVT wb_reg_pc_reg_36_ ( .D(n59), .CLK(n4306), .QN(csr_io_pc[36]) );
  DFFX1_LVT wb_reg_pc_reg_35_ ( .D(n58), .CLK(n4306), .QN(csr_io_pc[35]) );
  DFFX1_LVT wb_reg_pc_reg_34_ ( .D(n57), .CLK(n4306), .QN(csr_io_pc[34]) );
  DFFX1_LVT wb_reg_pc_reg_33_ ( .D(n56), .CLK(n4306), .QN(csr_io_pc[33]) );
  DFFX1_LVT wb_reg_pc_reg_32_ ( .D(n55), .CLK(n4306), .QN(csr_io_pc[32]) );
  DFFX1_LVT wb_reg_pc_reg_31_ ( .D(n54), .CLK(n4306), .QN(csr_io_pc[31]) );
  DFFX1_LVT wb_reg_pc_reg_30_ ( .D(n53), .CLK(n4307), .QN(csr_io_pc[30]) );
  DFFX1_LVT wb_reg_pc_reg_29_ ( .D(n52), .CLK(n4307), .QN(csr_io_pc[29]) );
  DFFX1_LVT wb_reg_pc_reg_28_ ( .D(n51), .CLK(n4307), .QN(csr_io_pc[28]) );
  DFFX1_LVT wb_reg_pc_reg_27_ ( .D(n50), .CLK(n4307), .QN(csr_io_pc[27]) );
  DFFX1_LVT wb_reg_pc_reg_26_ ( .D(n49), .CLK(n4307), .QN(csr_io_pc[26]) );
  DFFX1_LVT wb_reg_pc_reg_25_ ( .D(n48), .CLK(n4307), .QN(csr_io_pc[25]) );
  DFFX1_LVT wb_reg_pc_reg_24_ ( .D(n47), .CLK(n4307), .QN(csr_io_pc[24]) );
  DFFX1_LVT wb_reg_pc_reg_23_ ( .D(n46), .CLK(n4307), .QN(csr_io_pc[23]) );
  DFFX1_LVT wb_reg_pc_reg_22_ ( .D(n45), .CLK(n4307), .QN(csr_io_pc[22]) );
  DFFX1_LVT wb_reg_pc_reg_21_ ( .D(n44), .CLK(n4307), .QN(csr_io_pc[21]) );
  DFFX1_LVT wb_reg_pc_reg_20_ ( .D(n43), .CLK(n4307), .QN(csr_io_pc[20]) );
  DFFX1_LVT wb_reg_pc_reg_19_ ( .D(n42), .CLK(n4307), .QN(csr_io_pc[19]) );
  DFFX1_LVT wb_reg_pc_reg_18_ ( .D(n41), .CLK(n4308), .QN(csr_io_pc[18]) );
  DFFX1_LVT wb_reg_pc_reg_17_ ( .D(n40), .CLK(n4308), .QN(csr_io_pc[17]) );
  DFFX1_LVT wb_reg_pc_reg_16_ ( .D(n39), .CLK(n4308), .QN(csr_io_pc[16]) );
  DFFX1_LVT wb_reg_pc_reg_15_ ( .D(n38), .CLK(n4308), .QN(csr_io_pc[15]) );
  DFFX1_LVT wb_reg_pc_reg_14_ ( .D(n37), .CLK(n4308), .QN(csr_io_pc[14]) );
  DFFX1_LVT wb_reg_pc_reg_13_ ( .D(n36), .CLK(n4308), .QN(csr_io_pc[13]) );
  DFFX1_LVT wb_reg_pc_reg_12_ ( .D(n35), .CLK(n4308), .QN(csr_io_pc[12]) );
  DFFX1_LVT wb_reg_pc_reg_11_ ( .D(n34), .CLK(n4308), .QN(csr_io_pc[11]) );
  DFFX1_LVT wb_reg_pc_reg_10_ ( .D(n33), .CLK(n4308), .QN(csr_io_pc[10]) );
  DFFX1_LVT wb_reg_pc_reg_9_ ( .D(n32), .CLK(n4308), .QN(csr_io_pc[9]) );
  DFFX1_LVT wb_reg_pc_reg_8_ ( .D(n31), .CLK(n4308), .QN(csr_io_pc[8]) );
  DFFX1_LVT wb_reg_pc_reg_7_ ( .D(n30), .CLK(n4308), .QN(csr_io_pc[7]) );
  DFFX1_LVT wb_reg_pc_reg_6_ ( .D(n29), .CLK(n4309), .QN(csr_io_pc[6]) );
  DFFX1_LVT wb_reg_pc_reg_5_ ( .D(n28), .CLK(n4309), .QN(csr_io_pc[5]) );
  DFFX1_LVT wb_reg_pc_reg_4_ ( .D(n27), .CLK(n4309), .QN(csr_io_pc[4]) );
  DFFX1_LVT wb_reg_pc_reg_3_ ( .D(n26), .CLK(n4309), .QN(csr_io_pc[3]) );
  DFFX1_LVT wb_reg_pc_reg_2_ ( .D(n25), .CLK(n4309), .QN(csr_io_pc[2]) );
  DFFX1_LVT wb_reg_pc_reg_1_ ( .D(n24), .CLK(n4309), .QN(csr_io_pc[1]) );
  DFFX1_LVT wb_reg_pc_reg_0_ ( .D(n23), .CLK(n4309), .QN(csr_io_pc[0]) );
  DFFX1_LVT wb_reg_mem_size_reg_1_ ( .D(n72), .CLK(n4309), .QN(
        io_imem_sfence_bits_rs2) );
  DFFX1_LVT wb_reg_mem_size_reg_0_ ( .D(n71), .CLK(n4309), .QN(
        io_imem_sfence_bits_rs1) );
  DFFX1_LVT wb_reg_inst_reg_31_ ( .D(n22), .CLK(n4309), .QN(csr_io_rw_addr[11]) );
  DFFX1_LVT wb_reg_inst_reg_30_ ( .D(n21), .CLK(n4309), .QN(csr_io_rw_addr[10]) );
  DFFX1_LVT wb_reg_inst_reg_29_ ( .D(n20), .CLK(n4309), .QN(csr_io_rw_addr[9])
         );
  DFFX1_LVT wb_reg_inst_reg_28_ ( .D(n19), .CLK(n4310), .QN(csr_io_rw_addr[8])
         );
  DFFX1_LVT wb_reg_inst_reg_27_ ( .D(n18), .CLK(n4310), .QN(csr_io_rw_addr[7])
         );
  DFFX1_LVT wb_reg_inst_reg_26_ ( .D(n17), .CLK(n4310), .QN(csr_io_rw_addr[6])
         );
  DFFX1_LVT wb_reg_inst_reg_25_ ( .D(n16), .CLK(n4310), .QN(csr_io_rw_addr[5])
         );
  DFFX1_LVT wb_reg_inst_reg_24_ ( .D(n15), .CLK(n4310), .QN(csr_io_rw_addr[4])
         );
  DFFX1_LVT wb_reg_inst_reg_23_ ( .D(n14), .CLK(n4310), .QN(csr_io_rw_addr[3])
         );
  DFFX1_LVT wb_reg_inst_reg_22_ ( .D(n13), .CLK(n4310), .QN(csr_io_rw_addr[2])
         );
  DFFX1_LVT wb_reg_inst_reg_21_ ( .D(n12), .CLK(n4310), .QN(csr_io_rw_addr[1])
         );
  DFFX1_LVT wb_reg_inst_reg_20_ ( .D(n11), .CLK(n4310), .QN(csr_io_rw_addr[0])
         );
  DFFX1_LVT wb_reg_inst_reg_11_ ( .D(n_T_849[4]), .CLK(n4310), .Q(wb_waddr[4]), 
        .QN(n3198) );
  DFFX1_LVT wb_reg_inst_reg_10_ ( .D(n2566), .CLK(n4310), .Q(wb_waddr[3]), 
        .QN(n3199) );
  DFFX1_LVT wb_reg_inst_reg_9_ ( .D(n_T_849[2]), .CLK(n4310), .Q(n3043), .QN(
        n3102) );
  DFFX1_LVT wb_reg_inst_reg_7_ ( .D(n_T_849[11]), .CLK(n4311), .Q(n3041), .QN(
        n3201) );
  DFFX1_LVT wb_reg_cause_reg_0_ ( .D(N533), .CLK(n4311), .Q(wb_reg_cause[0])
         );
  DFFX1_LVT wb_reg_cause_reg_2_ ( .D(N535), .CLK(n4311), .Q(wb_reg_cause[2])
         );
  DFFX1_LVT wb_reg_cause_reg_3_ ( .D(N536), .CLK(n4305), .QN(n3565) );
  DFFX1_LVT wb_reg_xcpt_reg ( .D(N529), .CLK(n3594), .Q(n3262), .QN(n576) );
  DFFX1_LVT ex_reg_rs_lsb_1_reg_0_ ( .D(N678), .CLK(n4312), .Q(n5481), .QN(
        n594) );
  DFFX1_LVT ex_reg_rs_lsb_1_reg_1_ ( .D(N679), .CLK(n4313), .Q(n_T_635[1]) );
  DFFX1_LVT mem_reg_rs2_reg_0_ ( .D(n_T_702[0]), .CLK(n4091), .Q(
        mem_reg_rs2[0]) );
  DFFX1_LVT mem_reg_rs2_reg_1_ ( .D(n_T_702[1]), .CLK(n4091), .Q(
        mem_reg_rs2[1]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_8_ ( .D(id_rs_1[10]), .CLK(n4079), .Q(
        n_T_635[10]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_9_ ( .D(id_rs_1[11]), .CLK(n4078), .Q(
        n_T_635[11]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_10_ ( .D(id_rs_1[12]), .CLK(n4078), .Q(
        n_T_635[12]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_11_ ( .D(id_rs_1[13]), .CLK(n4078), .Q(
        n_T_635[13]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_12_ ( .D(id_rs_1[14]), .CLK(n4078), .Q(
        n_T_635[14]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_13_ ( .D(id_rs_1[15]), .CLK(n4078), .Q(
        n_T_635[15]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_14_ ( .D(id_rs_1[16]), .CLK(n4078), .Q(
        n_T_635[16]) );
  DFFX1_LVT mem_reg_rs2_reg_16_ ( .D(N477), .CLK(n4091), .Q(mem_reg_rs2[16])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_15_ ( .D(id_rs_1[17]), .CLK(n4078), .Q(
        n_T_635[17]) );
  DFFX1_LVT mem_reg_rs2_reg_17_ ( .D(N478), .CLK(n4091), .Q(mem_reg_rs2[17])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_16_ ( .D(id_rs_1[18]), .CLK(n4078), .Q(
        n_T_635[18]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_17_ ( .D(id_rs_1[19]), .CLK(n4078), .Q(
        n_T_635[19]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_18_ ( .D(id_rs_1[20]), .CLK(n4078), .Q(
        n_T_635[20]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_19_ ( .D(id_rs_1[21]), .CLK(n4078), .Q(
        n_T_635[21]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_20_ ( .D(id_rs_1[22]), .CLK(n4078), .Q(
        n_T_635[22]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_21_ ( .D(id_rs_1[23]), .CLK(n4077), .Q(
        n_T_635[23]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_22_ ( .D(id_rs_1[24]), .CLK(n4077), .Q(
        n_T_635[24]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_23_ ( .D(id_rs_1[25]), .CLK(n4077), .Q(
        n_T_635[25]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_24_ ( .D(id_rs_1[26]), .CLK(n4077), .Q(
        n_T_635[26]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_25_ ( .D(id_rs_1[27]), .CLK(n4077), .Q(
        n_T_635[27]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_26_ ( .D(id_rs_1[28]), .CLK(n4077), .Q(
        n_T_635[28]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_27_ ( .D(id_rs_1[29]), .CLK(n4077), .Q(
        n_T_635[29]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_0_ ( .D(id_rs_1[2]), .CLK(n4077), .Q(
        n_T_635[2]) );
  DFFX1_LVT mem_reg_rs2_reg_26_ ( .D(N487), .CLK(n4090), .Q(mem_reg_rs2[26])
         );
  DFFX1_LVT mem_reg_rs2_reg_18_ ( .D(N479), .CLK(n4090), .Q(mem_reg_rs2[18])
         );
  DFFX1_LVT mem_reg_rs2_reg_10_ ( .D(N471), .CLK(n4090), .Q(mem_reg_rs2[10])
         );
  DFFX1_LVT mem_reg_rs2_reg_2_ ( .D(n_T_702[2]), .CLK(n4090), .Q(
        mem_reg_rs2[2]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_28_ ( .D(id_rs_1[30]), .CLK(n4077), .Q(
        n_T_635[30]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_29_ ( .D(id_rs_1[31]), .CLK(n4077), .Q(
        n_T_635[31]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_30_ ( .D(id_rs_1[32]), .CLK(n4077), .Q(
        n_T_635[32]) );
  DFFX1_LVT mem_reg_rs2_reg_32_ ( .D(N493), .CLK(n4090), .Q(mem_reg_rs2[32])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_31_ ( .D(id_rs_1[33]), .CLK(n4077), .Q(
        n_T_635[33]) );
  DFFX1_LVT mem_reg_rs2_reg_33_ ( .D(N494), .CLK(n4090), .Q(mem_reg_rs2[33])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_32_ ( .D(id_rs_1[34]), .CLK(n4076), .Q(
        n_T_635[34]) );
  DFFX1_LVT mem_reg_rs2_reg_34_ ( .D(N495), .CLK(n4090), .Q(mem_reg_rs2[34])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_33_ ( .D(id_rs_1[35]), .CLK(n4076), .Q(
        n_T_635[35]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_34_ ( .D(id_rs_1[36]), .CLK(n4076), .Q(
        n_T_635[36]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_35_ ( .D(id_rs_1[37]), .CLK(n4076), .Q(
        n_T_635[37]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_36_ ( .D(id_rs_1[38]), .CLK(n4076), .Q(
        n_T_635[38]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_37_ ( .D(id_rs_1[39]), .CLK(n4076), .Q(
        n_T_635[39]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_1_ ( .D(id_rs_1[3]), .CLK(n4076), .Q(
        n_T_635[3]) );
  DFFX1_LVT mem_reg_rs2_reg_35_ ( .D(N496), .CLK(n4090), .Q(mem_reg_rs2[35])
         );
  DFFX1_LVT mem_reg_rs2_reg_27_ ( .D(N488), .CLK(n4090), .Q(mem_reg_rs2[27])
         );
  DFFX1_LVT mem_reg_rs2_reg_19_ ( .D(N480), .CLK(n4090), .Q(mem_reg_rs2[19])
         );
  DFFX1_LVT mem_reg_rs2_reg_11_ ( .D(N472), .CLK(n4090), .Q(mem_reg_rs2[11])
         );
  DFFX1_LVT mem_reg_rs2_reg_3_ ( .D(n_T_702[3]), .CLK(n4090), .Q(
        mem_reg_rs2[3]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_38_ ( .D(id_rs_1[40]), .CLK(n4076), .Q(
        n_T_635[40]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_39_ ( .D(id_rs_1[41]), .CLK(n4076), .Q(
        n_T_635[41]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_40_ ( .D(id_rs_1[42]), .CLK(n4076), .Q(
        n_T_635[42]) );
  DFFX1_LVT mem_reg_rs2_reg_42_ ( .D(N503), .CLK(n4089), .Q(mem_reg_rs2[42])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_41_ ( .D(id_rs_1[43]), .CLK(n4076), .Q(
        n_T_635[43]) );
  DFFX1_LVT mem_reg_rs2_reg_43_ ( .D(N504), .CLK(n4089), .Q(mem_reg_rs2[43])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_42_ ( .D(id_rs_1[44]), .CLK(n4076), .Q(
        n_T_635[44]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_43_ ( .D(id_rs_1[45]), .CLK(n4075), .Q(
        n_T_635[45]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_44_ ( .D(id_rs_1[46]), .CLK(n4075), .Q(
        n_T_635[46]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_45_ ( .D(id_rs_1[47]), .CLK(n4075), .Q(
        n_T_635[47]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_46_ ( .D(id_rs_1[48]), .CLK(n4075), .Q(
        n_T_635[48]) );
  DFFX1_LVT mem_reg_rs2_reg_48_ ( .D(N509), .CLK(n4089), .Q(mem_reg_rs2[48])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_47_ ( .D(id_rs_1[49]), .CLK(n4075), .Q(
        n_T_635[49]) );
  DFFX1_LVT mem_reg_rs2_reg_49_ ( .D(N510), .CLK(n4089), .Q(mem_reg_rs2[49])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_2_ ( .D(id_rs_1[4]), .CLK(n4075), .Q(
        n_T_635[4]) );
  DFFX1_LVT mem_reg_rs2_reg_36_ ( .D(N497), .CLK(n4089), .Q(mem_reg_rs2[36])
         );
  DFFX1_LVT mem_reg_rs2_reg_28_ ( .D(N489), .CLK(n4089), .Q(mem_reg_rs2[28])
         );
  DFFX1_LVT mem_reg_rs2_reg_20_ ( .D(N481), .CLK(n4089), .Q(mem_reg_rs2[20])
         );
  DFFX1_LVT mem_reg_rs2_reg_44_ ( .D(N505), .CLK(n4089), .Q(mem_reg_rs2[44])
         );
  DFFX1_LVT mem_reg_rs2_reg_12_ ( .D(N473), .CLK(n4089), .Q(mem_reg_rs2[12])
         );
  DFFX1_LVT mem_reg_rs2_reg_4_ ( .D(n_T_702[4]), .CLK(n4089), .Q(
        mem_reg_rs2[4]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_48_ ( .D(id_rs_1[50]), .CLK(n4075), .Q(
        n_T_635[50]) );
  DFFX1_LVT mem_reg_rs2_reg_50_ ( .D(N511), .CLK(n4089), .Q(mem_reg_rs2[50])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_49_ ( .D(id_rs_1[51]), .CLK(n4075), .Q(
        n_T_635[51]) );
  DFFX1_LVT mem_reg_rs2_reg_51_ ( .D(N512), .CLK(n4089), .Q(mem_reg_rs2[51])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_50_ ( .D(id_rs_1[52]), .CLK(n4075), .Q(
        n_T_635[52]) );
  DFFX1_LVT mem_reg_rs2_reg_52_ ( .D(N513), .CLK(n4088), .Q(mem_reg_rs2[52])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_51_ ( .D(id_rs_1[53]), .CLK(n4075), .Q(
        n_T_635[53]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_52_ ( .D(id_rs_1[54]), .CLK(n4075), .Q(
        n_T_635[54]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_53_ ( .D(id_rs_1[55]), .CLK(n4075), .Q(
        n_T_635[55]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_54_ ( .D(id_rs_1[56]), .CLK(n4074), .Q(
        n_T_635[56]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_55_ ( .D(id_rs_1[57]), .CLK(n4074), .Q(
        n_T_635[57]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_56_ ( .D(id_rs_1[58]), .CLK(n4074), .Q(
        n_T_635[58]) );
  DFFX1_LVT mem_reg_rs2_reg_58_ ( .D(N519), .CLK(n4088), .Q(mem_reg_rs2[58])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_57_ ( .D(id_rs_1[59]), .CLK(n4074), .Q(
        n_T_635[59]) );
  DFFX1_LVT mem_reg_rs2_reg_59_ ( .D(N520), .CLK(n4088), .Q(mem_reg_rs2[59])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_3_ ( .D(id_rs_1[5]), .CLK(n4074), .Q(
        n_T_635[5]) );
  DFFX1_LVT mem_reg_rs2_reg_37_ ( .D(N498), .CLK(n4088), .Q(mem_reg_rs2[37])
         );
  DFFX1_LVT mem_reg_rs2_reg_29_ ( .D(N490), .CLK(n4088), .Q(mem_reg_rs2[29])
         );
  DFFX1_LVT mem_reg_rs2_reg_53_ ( .D(N514), .CLK(n4088), .Q(mem_reg_rs2[53])
         );
  DFFX1_LVT mem_reg_rs2_reg_21_ ( .D(N482), .CLK(n4088), .Q(mem_reg_rs2[21])
         );
  DFFX1_LVT mem_reg_rs2_reg_45_ ( .D(N506), .CLK(n4088), .Q(mem_reg_rs2[45])
         );
  DFFX1_LVT mem_reg_rs2_reg_13_ ( .D(N474), .CLK(n4088), .Q(mem_reg_rs2[13])
         );
  DFFX1_LVT mem_reg_rs2_reg_5_ ( .D(n_T_702[5]), .CLK(n4088), .Q(
        mem_reg_rs2[5]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_58_ ( .D(id_rs_1[60]), .CLK(n4074), .Q(
        n_T_635[60]) );
  DFFX1_LVT mem_reg_rs2_reg_60_ ( .D(N521), .CLK(n4088), .Q(mem_reg_rs2[60])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_59_ ( .D(id_rs_1[61]), .CLK(n4074), .Q(
        n_T_635[61]) );
  DFFX1_LVT mem_reg_rs2_reg_61_ ( .D(N522), .CLK(n4088), .Q(mem_reg_rs2[61])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_60_ ( .D(id_rs_1[62]), .CLK(n4074), .Q(
        n_T_635[62]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_4_ ( .D(id_rs_1[6]), .CLK(n4074), .Q(
        n_T_635[6]) );
  DFFX1_LVT mem_reg_rs2_reg_38_ ( .D(N499), .CLK(n4087), .Q(mem_reg_rs2[38])
         );
  DFFX1_LVT mem_reg_rs2_reg_62_ ( .D(N523), .CLK(n4087), .Q(mem_reg_rs2[62])
         );
  DFFX1_LVT mem_reg_rs2_reg_30_ ( .D(N491), .CLK(n4087), .Q(mem_reg_rs2[30])
         );
  DFFX1_LVT mem_reg_rs2_reg_54_ ( .D(N515), .CLK(n4087), .Q(mem_reg_rs2[54])
         );
  DFFX1_LVT mem_reg_rs2_reg_22_ ( .D(N483), .CLK(n4087), .Q(mem_reg_rs2[22])
         );
  DFFX1_LVT mem_reg_rs2_reg_46_ ( .D(N507), .CLK(n4087), .Q(mem_reg_rs2[46])
         );
  DFFX1_LVT mem_reg_rs2_reg_14_ ( .D(N475), .CLK(n4087), .Q(mem_reg_rs2[14])
         );
  DFFX1_LVT mem_reg_rs2_reg_6_ ( .D(n_T_702[6]), .CLK(n4087), .Q(
        mem_reg_rs2[6]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_5_ ( .D(id_rs_1[7]), .CLK(n4074), .Q(
        n_T_635[7]) );
  DFFX1_LVT mem_reg_rs2_reg_39_ ( .D(N500), .CLK(n4087), .Q(mem_reg_rs2[39])
         );
  DFFX1_LVT mem_reg_rs2_reg_63_ ( .D(N524), .CLK(n4087), .Q(mem_reg_rs2[63])
         );
  DFFX1_LVT mem_reg_rs2_reg_31_ ( .D(N492), .CLK(n4087), .Q(mem_reg_rs2[31])
         );
  DFFX1_LVT mem_reg_rs2_reg_55_ ( .D(N516), .CLK(n4087), .Q(mem_reg_rs2[55])
         );
  DFFX1_LVT mem_reg_rs2_reg_23_ ( .D(N484), .CLK(n4086), .Q(mem_reg_rs2[23])
         );
  DFFX1_LVT mem_reg_rs2_reg_47_ ( .D(N508), .CLK(n4086), .Q(mem_reg_rs2[47])
         );
  DFFX1_LVT mem_reg_rs2_reg_15_ ( .D(N476), .CLK(n4086), .Q(mem_reg_rs2[15])
         );
  DFFX1_LVT mem_reg_rs2_reg_7_ ( .D(n_T_702[7]), .CLK(n4086), .Q(
        mem_reg_rs2[7]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_6_ ( .D(id_rs_1[8]), .CLK(n4074), .Q(
        n_T_635[8]) );
  DFFX1_LVT mem_reg_rs2_reg_40_ ( .D(N501), .CLK(n4086), .Q(mem_reg_rs2[40])
         );
  DFFX1_LVT mem_reg_rs2_reg_56_ ( .D(N517), .CLK(n4086), .Q(mem_reg_rs2[56])
         );
  DFFX1_LVT mem_reg_rs2_reg_24_ ( .D(N485), .CLK(n4086), .Q(mem_reg_rs2[24])
         );
  DFFX1_LVT mem_reg_rs2_reg_8_ ( .D(N469), .CLK(n4086), .Q(mem_reg_rs2[8]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_7_ ( .D(id_rs_1[9]), .CLK(n4074), .Q(
        n_T_635[9]) );
  DFFX1_LVT mem_reg_rs2_reg_41_ ( .D(N502), .CLK(n4086), .Q(mem_reg_rs2[41])
         );
  DFFX1_LVT mem_reg_rs2_reg_57_ ( .D(N518), .CLK(n4086), .Q(mem_reg_rs2[57])
         );
  DFFX1_LVT mem_reg_rs2_reg_25_ ( .D(N486), .CLK(n4086), .Q(mem_reg_rs2[25])
         );
  DFFX1_LVT mem_reg_rs2_reg_9_ ( .D(N470), .CLK(n4086), .Q(mem_reg_rs2[9]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_60_ ( .D(N742), .CLK(n4085), .Q(n_T_628[62])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_58_ ( .D(N740), .CLK(n4084), .Q(n_T_628[60])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_57_ ( .D(N739), .CLK(n4084), .Q(n_T_628[59])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_55_ ( .D(N737), .CLK(n4084), .Q(n_T_628[57])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_54_ ( .D(N736), .CLK(n4084), .Q(n_T_628[56])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_52_ ( .D(N734), .CLK(n4084), .Q(n_T_628[54])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_51_ ( .D(N733), .CLK(n4084), .Q(n_T_628[53])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_49_ ( .D(N731), .CLK(n4084), .Q(n_T_628[51])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_48_ ( .D(N730), .CLK(n4084), .Q(n_T_628[50])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_47_ ( .D(N729), .CLK(n4083), .Q(n_T_628[49])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_46_ ( .D(N728), .CLK(n4083), .Q(n_T_628[48])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_45_ ( .D(N727), .CLK(n4083), .Q(n_T_628[47])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_44_ ( .D(N726), .CLK(n4083), .Q(n_T_628[46])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_43_ ( .D(N725), .CLK(n4083), .Q(n_T_628[45])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_42_ ( .D(N724), .CLK(n4083), .Q(n_T_628[44])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_41_ ( .D(N723), .CLK(n4083), .Q(n_T_628[43])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_40_ ( .D(N722), .CLK(n4083), .Q(n_T_628[42])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_37_ ( .D(N719), .CLK(n4083), .Q(n_T_628[39])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_36_ ( .D(N718), .CLK(n4083), .Q(n_T_628[38])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_35_ ( .D(N717), .CLK(n4082), .Q(n_T_628[37])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_34_ ( .D(N716), .CLK(n4082), .Q(n_T_628[36])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_31_ ( .D(N713), .CLK(n4082), .Q(n_T_628[33])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_30_ ( .D(N712), .CLK(n4082), .Q(n_T_628[32])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_29_ ( .D(N711), .CLK(n4082), .Q(n_T_628[31])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_28_ ( .D(N710), .CLK(n4082), .Q(n_T_628[30])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_27_ ( .D(N709), .CLK(n4082), .Q(n_T_628[29])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_26_ ( .D(N708), .CLK(n4082), .Q(n_T_628[28])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_25_ ( .D(N707), .CLK(n4082), .Q(n_T_628[27])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_24_ ( .D(N706), .CLK(n4082), .Q(n_T_628[26])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_23_ ( .D(N705), .CLK(n4081), .Q(n_T_628[25])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_22_ ( .D(N704), .CLK(n4081), .Q(n_T_628[24])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_21_ ( .D(N703), .CLK(n4081), .Q(n_T_628[23])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_20_ ( .D(N702), .CLK(n4081), .Q(n_T_628[22])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_19_ ( .D(N701), .CLK(n4081), .Q(n_T_628[21])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_18_ ( .D(N700), .CLK(n4081), .Q(n_T_628[20])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_17_ ( .D(N699), .CLK(n4081), .Q(n_T_628[19])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_16_ ( .D(N698), .CLK(n4081), .Q(n_T_628[18])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_15_ ( .D(N697), .CLK(n4081), .Q(n_T_628[17])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_14_ ( .D(N696), .CLK(n4081), .Q(n_T_628[16])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_13_ ( .D(N695), .CLK(n4081), .Q(n_T_628[15])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_12_ ( .D(N694), .CLK(n4081), .Q(n_T_628[14])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_11_ ( .D(N693), .CLK(n4080), .Q(n_T_628[13])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_10_ ( .D(N692), .CLK(n4080), .Q(n_T_628[12])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_9_ ( .D(N691), .CLK(n4080), .Q(n_T_628[11]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_8_ ( .D(N690), .CLK(n4080), .Q(n_T_628[10]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_7_ ( .D(N689), .CLK(n4080), .Q(n_T_628[9]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_6_ ( .D(N688), .CLK(n4080), .Q(n_T_628[8]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_5_ ( .D(N687), .CLK(n4080), .Q(n_T_628[7]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_4_ ( .D(N686), .CLK(n4080), .Q(n_T_628[6]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_3_ ( .D(N685), .CLK(n4080), .Q(n_T_628[5]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_2_ ( .D(N684), .CLK(n4080), .Q(n_T_628[4]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_1_ ( .D(N683), .CLK(n4080), .Q(n_T_628[3]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_0_ ( .D(N682), .CLK(n4080), .Q(n_T_628[2]) );
  DFFX1_LVT ex_reg_rs_lsb_0_reg_1_ ( .D(N673), .CLK(n4312), .Q(n_T_628[1]), 
        .QN(n3255) );
  DFFX1_LVT ex_reg_rs_lsb_0_reg_0_ ( .D(N672), .CLK(n4313), .Q(n7019), .QN(
        n569) );
  DFFX1_LVT u_T_427_reg_0__63_ ( .D(n4494), .CLK(n4284), .Q(n_T_427[1942]), 
        .QN(n3529) );
  DFFX1_LVT u_T_427_reg_0__62_ ( .D(n4491), .CLK(n4284), .Q(n_T_427[1941]), 
        .QN(n3484) );
  DFFX1_LVT u_T_427_reg_0__61_ ( .D(n4488), .CLK(n4284), .Q(n_T_427[1940]), 
        .QN(n3483) );
  DFFX1_LVT u_T_427_reg_0__60_ ( .D(n4485), .CLK(n4284), .Q(n_T_427[1939]) );
  DFFX1_LVT u_T_427_reg_0__58_ ( .D(n4479), .CLK(n4283), .Q(n_T_427[1937]), 
        .QN(n3492) );
  DFFX1_LVT u_T_427_reg_0__56_ ( .D(n4473), .CLK(n4283), .Q(n_T_427[1935]), 
        .QN(n3564) );
  DFFX1_LVT u_T_427_reg_0__54_ ( .D(n4467), .CLK(n4283), .Q(n_T_427[1933]), 
        .QN(n3562) );
  DFFX1_LVT u_T_427_reg_0__52_ ( .D(n4461), .CLK(n4283), .Q(n_T_427[1931]), 
        .QN(n3560) );
  DFFX1_LVT u_T_427_reg_0__51_ ( .D(n4458), .CLK(n4283), .Q(n_T_427[1930]), 
        .QN(n3559) );
  DFFX1_LVT u_T_427_reg_0__49_ ( .D(n4452), .CLK(n4283), .Q(n_T_427[1929]), 
        .QN(n3558) );
  DFFX1_LVT u_T_427_reg_0__46_ ( .D(n4443), .CLK(n4282), .Q(n_T_427[1926]) );
  DFFX1_LVT u_T_427_reg_0__45_ ( .D(n4440), .CLK(n4282), .Q(n_T_427[1925]), 
        .QN(n3555) );
  DFFX1_LVT u_T_427_reg_0__44_ ( .D(n4437), .CLK(n4282), .Q(n_T_427[1924]), 
        .QN(n2496) );
  DFFX1_LVT u_T_427_reg_0__43_ ( .D(n4434), .CLK(n4282), .Q(n_T_427[1923]), 
        .QN(n3554) );
  DFFX1_LVT u_T_427_reg_0__42_ ( .D(n4431), .CLK(n4282), .Q(n_T_427[1922]), 
        .QN(n3553) );
  DFFX1_LVT u_T_427_reg_0__41_ ( .D(n4428), .CLK(n4282), .Q(n_T_427[1921]), 
        .QN(n3552) );
  DFFX1_LVT u_T_427_reg_0__39_ ( .D(n4422), .CLK(n4282), .Q(n_T_427[1919]) );
  DFFX1_LVT u_T_427_reg_0__38_ ( .D(n4420), .CLK(n4282), .Q(n_T_427[1918]) );
  DFFX1_LVT u_T_427_reg_0__36_ ( .D(n4414), .CLK(n4282), .Q(n_T_427[1916]), 
        .QN(n3549) );
  DFFX1_LVT u_T_427_reg_0__35_ ( .D(n4412), .CLK(n4281), .Q(n_T_427[1915]) );
  DFFX1_LVT u_T_427_reg_0__34_ ( .D(n4409), .CLK(n4281), .Q(n_T_427[1914]) );
  DFFX1_LVT u_T_427_reg_0__33_ ( .D(n4407), .CLK(n4281), .Q(n_T_427[1913]) );
  DFFX1_LVT u_T_427_reg_0__31_ ( .D(n4402), .CLK(n4281), .Q(n_T_427[1912]) );
  DFFX1_LVT u_T_427_reg_0__30_ ( .D(n4399), .CLK(n4281), .Q(n_T_427[1911]), 
        .QN(n3547) );
  DFFX1_LVT u_T_427_reg_0__29_ ( .D(n4396), .CLK(n4281), .Q(n_T_427[1910]) );
  DFFX1_LVT u_T_427_reg_0__28_ ( .D(n4394), .CLK(n4281), .Q(n_T_427[1909]) );
  DFFX1_LVT u_T_427_reg_0__27_ ( .D(n4391), .CLK(n4281), .Q(n_T_427[1908]) );
  DFFX1_LVT u_T_427_reg_0__26_ ( .D(n4389), .CLK(n4281), .Q(n_T_427[1907]) );
  DFFX1_LVT u_T_427_reg_0__25_ ( .D(n4387), .CLK(n4281), .Q(n_T_427[1906]) );
  DFFX1_LVT u_T_427_reg_0__24_ ( .D(n4384), .CLK(n4281), .Q(n_T_427[1905]), 
        .QN(n3545) );
  DFFX1_LVT u_T_427_reg_0__23_ ( .D(n4381), .CLK(n4280), .Q(n_T_427[1904]) );
  DFFX1_LVT u_T_427_reg_0__22_ ( .D(n4379), .CLK(n4280), .Q(n_T_427[1903]), 
        .QN(n2684) );
  DFFX1_LVT u_T_427_reg_0__21_ ( .D(n4377), .CLK(n4280), .Q(n_T_427[1902]) );
  DFFX1_LVT u_T_427_reg_0__20_ ( .D(n4374), .CLK(n4280), .Q(n_T_427[1901]), 
        .QN(n3544) );
  DFFX1_LVT u_T_427_reg_0__19_ ( .D(n4371), .CLK(n4280), .Q(n_T_427[1900]), 
        .QN(n3543) );
  DFFX1_LVT u_T_427_reg_0__18_ ( .D(n4368), .CLK(n4280), .Q(n_T_427[1899]), 
        .QN(n3542) );
  DFFX1_LVT u_T_427_reg_0__14_ ( .D(n4357), .CLK(n4280), .Q(n_T_427[1895]) );
  DFFX1_LVT u_T_427_reg_0__11_ ( .D(n4351), .CLK(n4279), .Q(n_T_427[1892]) );
  DFFX1_LVT u_T_427_reg_0__5_ ( .D(n4331), .CLK(n4279), .Q(n_T_427[1886]) );
  DFFX1_LVT u_T_427_reg_0__4_ ( .D(n4328), .CLK(n4279), .Q(n_T_427[1885]) );
  DFFX1_LVT u_T_427_reg_0__2_ ( .D(n4322), .CLK(n4279), .Q(n_T_427[1884]) );
  DFFX1_LVT u_T_427_reg_0__0_ ( .D(n4316), .CLK(n4279), .Q(n_T_427[1882]), 
        .QN(n3490) );
  DFFX1_LVT u_T_427_reg_1__63_ ( .D(n4494), .CLK(n4278), .QN(n3170) );
  DFFX1_LVT u_T_427_reg_1__62_ ( .D(n4491), .CLK(n4278), .QN(n3169) );
  DFFX1_LVT u_T_427_reg_1__61_ ( .D(n4488), .CLK(n4278), .QN(n3167) );
  DFFX1_LVT u_T_427_reg_1__60_ ( .D(n4485), .CLK(n4278), .Q(n_T_427[1881]), 
        .QN(n3409) );
  DFFX1_LVT u_T_427_reg_1__59_ ( .D(n4482), .CLK(n4277), .QN(n3165) );
  DFFX1_LVT u_T_427_reg_1__58_ ( .D(n4481), .CLK(n4277), .QN(n3164) );
  DFFX1_LVT u_T_427_reg_1__57_ ( .D(n4476), .CLK(n4277), .QN(n3163) );
  DFFX1_LVT u_T_427_reg_1__56_ ( .D(n4475), .CLK(n4277), .QN(n3162) );
  DFFX1_LVT u_T_427_reg_1__55_ ( .D(n4470), .CLK(n4277), .QN(n3160) );
  DFFX1_LVT u_T_427_reg_1__54_ ( .D(n4469), .CLK(n4277), .QN(n3159) );
  DFFX1_LVT u_T_427_reg_1__53_ ( .D(n4464), .CLK(n4277), .QN(n3158) );
  DFFX1_LVT u_T_427_reg_1__52_ ( .D(n4463), .CLK(n4277), .QN(n3157) );
  DFFX1_LVT u_T_427_reg_1__51_ ( .D(n4460), .CLK(n4277), .QN(n3156) );
  DFFX1_LVT u_T_427_reg_1__50_ ( .D(n4455), .CLK(n4277), .QN(n3155) );
  DFFX1_LVT u_T_427_reg_1__49_ ( .D(n4454), .CLK(n4277), .QN(n3154) );
  DFFX1_LVT u_T_427_reg_1__48_ ( .D(n4449), .CLK(n4277), .QN(n3153) );
  DFFX1_LVT u_T_427_reg_1__47_ ( .D(n4446), .CLK(n4276), .QN(n3152) );
  DFFX1_LVT u_T_427_reg_1__45_ ( .D(n4442), .CLK(n4276), .QN(n3151) );
  DFFX1_LVT u_T_427_reg_1__43_ ( .D(n4436), .CLK(n4276), .QN(n3150) );
  DFFX1_LVT u_T_427_reg_1__42_ ( .D(n4433), .CLK(n4276), .QN(n3149) );
  DFFX1_LVT u_T_427_reg_1__41_ ( .D(n4430), .CLK(n4276), .QN(n3148) );
  DFFX1_LVT u_T_427_reg_1__40_ ( .D(n4425), .CLK(n4276), .QN(n3147) );
  DFFX1_LVT u_T_427_reg_1__37_ ( .D(n4417), .CLK(n4276), .QN(n3146) );
  DFFX1_LVT u_T_427_reg_1__36_ ( .D(n4416), .CLK(n4276), .QN(n3145) );
  DFFX1_LVT u_T_427_reg_1__32_ ( .D(n4404), .CLK(n4275), .QN(n3144) );
  DFFX1_LVT u_T_427_reg_1__30_ ( .D(n4401), .CLK(n4275), .QN(n3140) );
  DFFX1_LVT u_T_427_reg_1__29_ ( .D(n4398), .CLK(n4275), .Q(n_T_427[1872]), 
        .QN(n3375) );
  DFFX1_LVT u_T_427_reg_1__27_ ( .D(n4391), .CLK(n4275), .Q(n_T_427[1870]), 
        .QN(n3330) );
  DFFX1_LVT u_T_427_reg_1__24_ ( .D(n4386), .CLK(n4275), .QN(n3137) );
  DFFX1_LVT u_T_427_reg_1__20_ ( .D(n4376), .CLK(n4274), .Q(n_T_427[1865]), 
        .QN(n3322) );
  DFFX1_LVT u_T_427_reg_1__19_ ( .D(n4373), .CLK(n4274), .Q(n_T_427[1864]), 
        .QN(n3319) );
  DFFX1_LVT u_T_427_reg_1__18_ ( .D(n4370), .CLK(n4274), .Q(n_T_427[1863]), 
        .QN(n3316) );
  DFFX1_LVT u_T_427_reg_1__17_ ( .D(n4365), .CLK(n4274), .QN(n3139) );
  DFFX1_LVT u_T_427_reg_1__16_ ( .D(n4362), .CLK(n4274), .Q(n_T_427[1862]), 
        .QN(n3178) );
  DFFX1_LVT u_T_427_reg_1__15_ ( .D(n4360), .CLK(n4274), .Q(n_T_427[1861]) );
  DFFX1_LVT u_T_427_reg_1__14_ ( .D(n4357), .CLK(n4274), .Q(n_T_427[1860]) );
  DFFX1_LVT u_T_427_reg_1__13_ ( .D(n4355), .CLK(n4274), .Q(n_T_427[1859]) );
  DFFX1_LVT u_T_427_reg_1__12_ ( .D(n4352), .CLK(n4274), .Q(n_T_427[1858]) );
  DFFX1_LVT u_T_427_reg_1__11_ ( .D(n4351), .CLK(n4273), .Q(n_T_427[1857]) );
  DFFX1_LVT u_T_427_reg_1__10_ ( .D(n4346), .CLK(n4273), .Q(n_T_427[1856]) );
  DFFX1_LVT u_T_427_reg_1__9_ ( .D(n4343), .CLK(n4273), .Q(n_T_427[1855]) );
  DFFX1_LVT u_T_427_reg_1__8_ ( .D(n4340), .CLK(n4273), .Q(n_T_427[1854]) );
  DFFX1_LVT u_T_427_reg_1__7_ ( .D(n4337), .CLK(n4273), .Q(n_T_427[1853]) );
  DFFX1_LVT u_T_427_reg_1__6_ ( .D(n4334), .CLK(n4273), .Q(n_T_427[1852]) );
  DFFX1_LVT u_T_427_reg_1__5_ ( .D(n4331), .CLK(n4273), .Q(n_T_427[1851]) );
  DFFX1_LVT u_T_427_reg_1__4_ ( .D(n4328), .CLK(n4273), .Q(n_T_427[1850]) );
  DFFX1_LVT u_T_427_reg_1__3_ ( .D(n4325), .CLK(n4273), .Q(n_T_427[1849]) );
  DFFX1_LVT u_T_427_reg_1__2_ ( .D(n4322), .CLK(n4273), .Q(n_T_427[1848]) );
  DFFX1_LVT u_T_427_reg_1__1_ ( .D(n4321), .CLK(n4273), .QN(n3654) );
  DFFX1_LVT u_T_427_reg_1__0_ ( .D(n4318), .CLK(n4273), .QN(n3633) );
  DFFX1_LVT u_T_427_reg_2__63_ ( .D(n4494), .CLK(n4272), .QN(n3171) );
  DFFX1_LVT u_T_427_reg_2__62_ ( .D(n4491), .CLK(n4272), .Q(n_T_427[1847]), 
        .QN(n3411) );
  DFFX1_LVT u_T_427_reg_2__61_ ( .D(n4488), .CLK(n4272), .QN(n3168) );
  DFFX1_LVT u_T_427_reg_2__60_ ( .D(n4485), .CLK(n4272), .Q(n_T_427[1846]), 
        .QN(n3410) );
  DFFX1_LVT u_T_427_reg_2__59_ ( .D(n4482), .CLK(n4271), .QN(n3166) );
  DFFX1_LVT u_T_427_reg_2__58_ ( .D(n4481), .CLK(n4271), .Q(n_T_427[1845]), 
        .QN(n3474) );
  DFFX1_LVT u_T_427_reg_2__56_ ( .D(n4475), .CLK(n4271), .Q(n_T_427[1843]), 
        .QN(n3472) );
  DFFX1_LVT u_T_427_reg_2__55_ ( .D(n4470), .CLK(n4271), .QN(n3161) );
  DFFX1_LVT u_T_427_reg_2__54_ ( .D(n4469), .CLK(n4271), .Q(n_T_427[1842]), 
        .QN(n3471) );
  DFFX1_LVT u_T_427_reg_2__52_ ( .D(n4463), .CLK(n4271), .Q(n_T_427[1840]), 
        .QN(n3469) );
  DFFX1_LVT u_T_427_reg_2__51_ ( .D(n4460), .CLK(n4271), .Q(n_T_427[1839]), 
        .QN(n3412) );
  DFFX1_LVT u_T_427_reg_2__49_ ( .D(n4454), .CLK(n4271), .Q(n_T_427[1837]), 
        .QN(n3468) );
  DFFX1_LVT u_T_427_reg_2__45_ ( .D(n4442), .CLK(n4270), .Q(n_T_427[1833]), 
        .QN(n3413) );
  DFFX1_LVT u_T_427_reg_2__43_ ( .D(n4436), .CLK(n4270), .Q(n_T_427[1831]), 
        .QN(n3464) );
  DFFX1_LVT u_T_427_reg_2__42_ ( .D(n4433), .CLK(n4270), .Q(n_T_427[1830]), 
        .QN(n3462) );
  DFFX1_LVT u_T_427_reg_2__41_ ( .D(n4430), .CLK(n4270), .Q(n_T_427[1829]), 
        .QN(n3475) );
  DFFX1_LVT u_T_427_reg_2__36_ ( .D(n4416), .CLK(n4270), .Q(n_T_427[1824]), 
        .QN(n3454) );
  DFFX1_LVT u_T_427_reg_2__32_ ( .D(n4404), .CLK(n4269), .QN(n3143) );
  DFFX1_LVT u_T_427_reg_2__30_ ( .D(n4401), .CLK(n4269), .Q(n_T_427[1819]), 
        .QN(n3451) );
  DFFX1_LVT u_T_427_reg_2__29_ ( .D(n4398), .CLK(n4269), .Q(n_T_427[1818]), 
        .QN(n3396) );
  DFFX1_LVT u_T_427_reg_2__27_ ( .D(n4391), .CLK(n4269), .Q(n_T_427[1816]), 
        .QN(n3450) );
  DFFX1_LVT u_T_427_reg_2__24_ ( .D(n4386), .CLK(n4269), .Q(n_T_427[1813]), 
        .QN(n3449) );
  DFFX1_LVT u_T_427_reg_2__20_ ( .D(n4376), .CLK(n4268), .Q(n_T_427[1809]), 
        .QN(n3447) );
  DFFX1_LVT u_T_427_reg_2__19_ ( .D(n4373), .CLK(n4268), .Q(n_T_427[1808]), 
        .QN(n3446) );
  DFFX1_LVT u_T_427_reg_2__18_ ( .D(n4370), .CLK(n4268), .Q(n_T_427[1807]), 
        .QN(n3445) );
  DFFX1_LVT u_T_427_reg_2__17_ ( .D(n4365), .CLK(n4268), .QN(n3142) );
  DFFX1_LVT u_T_427_reg_2__15_ ( .D(n4360), .CLK(n4268), .Q(n_T_427[1805]) );
  DFFX1_LVT u_T_427_reg_2__14_ ( .D(n4357), .CLK(n4268), .Q(n_T_427[1804]) );
  DFFX1_LVT u_T_427_reg_2__13_ ( .D(n4355), .CLK(n4268), .Q(n_T_427[1803]) );
  DFFX1_LVT u_T_427_reg_2__12_ ( .D(n4352), .CLK(n4268), .Q(n_T_427[1802]) );
  DFFX1_LVT u_T_427_reg_2__11_ ( .D(n4351), .CLK(n4267), .Q(n_T_427[1801]) );
  DFFX1_LVT u_T_427_reg_2__10_ ( .D(n4346), .CLK(n4267), .Q(n_T_427[1800]) );
  DFFX1_LVT u_T_427_reg_2__9_ ( .D(n4343), .CLK(n4267), .Q(n_T_427[1799]) );
  DFFX1_LVT u_T_427_reg_2__8_ ( .D(n4340), .CLK(n4267), .Q(n_T_427[1798]) );
  DFFX1_LVT u_T_427_reg_2__7_ ( .D(n4337), .CLK(n4267), .Q(n_T_427[1797]) );
  DFFX1_LVT u_T_427_reg_2__6_ ( .D(n4334), .CLK(n4267), .Q(n_T_427[1796]) );
  DFFX1_LVT u_T_427_reg_2__5_ ( .D(n4331), .CLK(n4267), .Q(n_T_427[1795]) );
  DFFX1_LVT u_T_427_reg_2__4_ ( .D(n4328), .CLK(n4267), .Q(n_T_427[1794]) );
  DFFX1_LVT u_T_427_reg_2__3_ ( .D(n4325), .CLK(n4267), .Q(n_T_427[1793]) );
  DFFX1_LVT u_T_427_reg_2__2_ ( .D(n4322), .CLK(n4267), .Q(n_T_427[1792]) );
  DFFX1_LVT u_T_427_reg_2__1_ ( .D(n4321), .CLK(n4267), .QN(n3138) );
  DFFX1_LVT u_T_427_reg_2__0_ ( .D(n4318), .CLK(n4267), .Q(n_T_427[1791]), 
        .QN(n3311) );
  DFFX1_LVT u_T_427_reg_3__63_ ( .D(n4494), .CLK(n4266), .Q(n_T_427[1790]), 
        .QN(n3488) );
  DFFX1_LVT u_T_427_reg_3__62_ ( .D(n4491), .CLK(n4266), .Q(n_T_427[1789]), 
        .QN(n3487) );
  DFFX1_LVT u_T_427_reg_3__61_ ( .D(n4488), .CLK(n4266), .Q(n_T_427[1788]), 
        .QN(n3485) );
  DFFX1_LVT u_T_427_reg_3__60_ ( .D(n4485), .CLK(n4266), .Q(n_T_427[1787]) );
  DFFX1_LVT u_T_427_reg_3__58_ ( .D(n4481), .CLK(n4265), .Q(n_T_427[1785]), 
        .QN(n3516) );
  DFFX1_LVT u_T_427_reg_3__56_ ( .D(n4475), .CLK(n4265), .Q(n_T_427[1783]), 
        .QN(n3514) );
  DFFX1_LVT u_T_427_reg_3__54_ ( .D(n4469), .CLK(n4265), .Q(n_T_427[1781]), 
        .QN(n3511) );
  DFFX1_LVT u_T_427_reg_3__52_ ( .D(n4463), .CLK(n4265), .Q(n_T_427[1779]), 
        .QN(n3509) );
  DFFX1_LVT u_T_427_reg_3__51_ ( .D(n4460), .CLK(n4265), .Q(n_T_427[1778]), 
        .QN(n3508) );
  DFFX1_LVT u_T_427_reg_3__49_ ( .D(n4454), .CLK(n4265), .Q(n_T_427[1776]), 
        .QN(n3506) );
  DFFX1_LVT u_T_427_reg_3__46_ ( .D(n4443), .CLK(n4264), .Q(n_T_427[1773]) );
  DFFX1_LVT u_T_427_reg_3__45_ ( .D(n4442), .CLK(n4264), .Q(n_T_427[1772]), 
        .QN(n3503) );
  DFFX1_LVT u_T_427_reg_3__44_ ( .D(n4437), .CLK(n4264), .Q(n_T_427[1771]) );
  DFFX1_LVT u_T_427_reg_3__43_ ( .D(n4436), .CLK(n4264), .Q(n_T_427[1770]), 
        .QN(n3502) );
  DFFX1_LVT u_T_427_reg_3__42_ ( .D(n4433), .CLK(n4264), .Q(n_T_427[1769]), 
        .QN(n3501) );
  DFFX1_LVT u_T_427_reg_3__41_ ( .D(n4430), .CLK(n4264), .Q(n_T_427[1768]), 
        .QN(n3500) );
  DFFX1_LVT u_T_427_reg_3__39_ ( .D(n4422), .CLK(n4264), .Q(n_T_427[1766]) );
  DFFX1_LVT u_T_427_reg_3__38_ ( .D(n4420), .CLK(n4264), .Q(n_T_427[1765]) );
  DFFX1_LVT u_T_427_reg_3__36_ ( .D(n4416), .CLK(n4264), .Q(n_T_427[1763]), 
        .QN(n3497) );
  DFFX1_LVT u_T_427_reg_3__35_ ( .D(n4412), .CLK(n4263), .Q(n_T_427[1762]) );
  DFFX1_LVT u_T_427_reg_3__34_ ( .D(n4409), .CLK(n4263), .Q(n_T_427[1761]) );
  DFFX1_LVT u_T_427_reg_3__33_ ( .D(n4407), .CLK(n4263), .Q(n_T_427[1760]) );
  DFFX1_LVT u_T_427_reg_3__31_ ( .D(n4402), .CLK(n4263), .Q(n_T_427[1758]) );
  DFFX1_LVT u_T_427_reg_3__30_ ( .D(n4401), .CLK(n4263), .Q(n_T_427[1757]), 
        .QN(n3548) );
  DFFX1_LVT u_T_427_reg_3__29_ ( .D(n4398), .CLK(n4263), .Q(n_T_427[1756]) );
  DFFX1_LVT u_T_427_reg_3__28_ ( .D(n4394), .CLK(n4263), .Q(n_T_427[1755]) );
  DFFX1_LVT u_T_427_reg_3__27_ ( .D(n4391), .CLK(n4263), .Q(n_T_427[1754]) );
  DFFX1_LVT u_T_427_reg_3__26_ ( .D(n4389), .CLK(n4263), .Q(n_T_427[1753]) );
  DFFX1_LVT u_T_427_reg_3__25_ ( .D(n4387), .CLK(n4263), .Q(n_T_427[1752]) );
  DFFX1_LVT u_T_427_reg_3__24_ ( .D(n4386), .CLK(n4263), .Q(n_T_427[1751]), 
        .QN(n3546) );
  DFFX1_LVT u_T_427_reg_3__23_ ( .D(n4381), .CLK(n4262), .Q(n_T_427[1750]) );
  DFFX1_LVT u_T_427_reg_3__22_ ( .D(n4379), .CLK(n4262), .Q(n_T_427[1749]) );
  DFFX1_LVT u_T_427_reg_3__21_ ( .D(n4377), .CLK(n4262), .Q(n_T_427[1748]) );
  DFFX1_LVT u_T_427_reg_3__20_ ( .D(n4376), .CLK(n4262), .Q(n_T_427[1747]) );
  DFFX1_LVT u_T_427_reg_3__19_ ( .D(n4373), .CLK(n4262), .Q(n_T_427[1746]) );
  DFFX1_LVT u_T_427_reg_3__18_ ( .D(n4370), .CLK(n4262), .Q(n_T_427[1745]) );
  DFFX1_LVT u_T_427_reg_3__16_ ( .D(n4362), .CLK(n4262), .Q(n_T_427[1743]) );
  DFFX1_LVT u_T_427_reg_3__15_ ( .D(n4360), .CLK(n4262), .Q(n_T_427[1742]) );
  DFFX1_LVT u_T_427_reg_3__14_ ( .D(n4357), .CLK(n4262), .Q(n_T_427[1741]) );
  DFFX1_LVT u_T_427_reg_3__13_ ( .D(n4355), .CLK(n4262), .Q(n_T_427[1740]) );
  DFFX1_LVT u_T_427_reg_3__12_ ( .D(n4352), .CLK(n4262), .Q(n_T_427[1739]) );
  DFFX1_LVT u_T_427_reg_3__11_ ( .D(n4351), .CLK(n4261), .Q(n_T_427[1738]) );
  DFFX1_LVT u_T_427_reg_3__10_ ( .D(n4346), .CLK(n4261), .Q(n_T_427[1737]) );
  DFFX1_LVT u_T_427_reg_3__9_ ( .D(n4343), .CLK(n4261), .Q(n_T_427[1736]) );
  DFFX1_LVT u_T_427_reg_3__8_ ( .D(n4340), .CLK(n4261), .Q(n_T_427[1735]) );
  DFFX1_LVT u_T_427_reg_3__7_ ( .D(n4337), .CLK(n4261), .Q(n_T_427[1734]) );
  DFFX1_LVT u_T_427_reg_3__6_ ( .D(n4334), .CLK(n4261), .Q(n_T_427[1733]) );
  DFFX1_LVT u_T_427_reg_3__5_ ( .D(n4331), .CLK(n4261), .Q(n_T_427[1732]) );
  DFFX1_LVT u_T_427_reg_3__4_ ( .D(n4328), .CLK(n4261), .Q(n_T_427[1731]) );
  DFFX1_LVT u_T_427_reg_3__3_ ( .D(n4325), .CLK(n4261), .Q(n_T_427[1730]) );
  DFFX1_LVT u_T_427_reg_3__2_ ( .D(n4322), .CLK(n4261), .Q(n_T_427[1729]) );
  DFFX1_LVT u_T_427_reg_3__1_ ( .D(n4321), .CLK(n4261), .Q(n_T_427[1728]), 
        .QN(n3257) );
  DFFX1_LVT u_T_427_reg_3__0_ ( .D(n4318), .CLK(n4261), .Q(n_T_427[1727]), 
        .QN(n3256) );
  DFFX1_LVT u_T_427_reg_4__63_ ( .D(n4494), .CLK(n4260), .Q(n_T_427[1726]), 
        .QN(n3489) );
  DFFX1_LVT u_T_427_reg_4__62_ ( .D(n4491), .CLK(n4260), .Q(n_T_427[1725]) );
  DFFX1_LVT u_T_427_reg_4__61_ ( .D(n4488), .CLK(n4260), .Q(n_T_427[1724]), 
        .QN(n3486) );
  DFFX1_LVT u_T_427_reg_4__60_ ( .D(n4485), .CLK(n4260), .Q(n_T_427[1723]) );
  DFFX1_LVT u_T_427_reg_4__58_ ( .D(n4481), .CLK(n4259), .Q(n_T_427[1721]) );
  DFFX1_LVT u_T_427_reg_4__57_ ( .D(n4476), .CLK(n4259), .Q(n_T_427[1720]) );
  DFFX1_LVT u_T_427_reg_4__56_ ( .D(n4475), .CLK(n4259), .Q(n_T_427[1719]) );
  DFFX1_LVT u_T_427_reg_4__54_ ( .D(n4469), .CLK(n4259), .Q(n_T_427[1717]) );
  DFFX1_LVT u_T_427_reg_4__53_ ( .D(n4464), .CLK(n4259), .Q(n_T_427[1716]) );
  DFFX1_LVT u_T_427_reg_4__52_ ( .D(n4463), .CLK(n4259), .Q(n_T_427[1715]) );
  DFFX1_LVT u_T_427_reg_4__51_ ( .D(n4460), .CLK(n4259), .Q(n_T_427[1714]) );
  DFFX1_LVT u_T_427_reg_4__50_ ( .D(n4455), .CLK(n4259), .Q(n_T_427[1713]) );
  DFFX1_LVT u_T_427_reg_4__49_ ( .D(n4454), .CLK(n4259), .Q(n_T_427[1712]) );
  DFFX1_LVT u_T_427_reg_4__48_ ( .D(n4449), .CLK(n4259), .Q(n_T_427[1711]) );
  DFFX1_LVT u_T_427_reg_4__47_ ( .D(n4446), .CLK(n4258), .Q(n_T_427[1710]) );
  DFFX1_LVT u_T_427_reg_4__46_ ( .D(n4443), .CLK(n4258), .Q(n_T_427[1709]) );
  DFFX1_LVT u_T_427_reg_4__45_ ( .D(n4442), .CLK(n4258), .Q(n_T_427[1708]) );
  DFFX1_LVT u_T_427_reg_4__44_ ( .D(n4437), .CLK(n4258), .Q(n_T_427[1707]) );
  DFFX1_LVT u_T_427_reg_4__43_ ( .D(n4436), .CLK(n4258), .Q(n_T_427[1706]) );
  DFFX1_LVT u_T_427_reg_4__42_ ( .D(n4433), .CLK(n4258), .Q(n_T_427[1705]) );
  DFFX1_LVT u_T_427_reg_4__41_ ( .D(n4430), .CLK(n4258), .Q(n_T_427[1704]), 
        .QN(n2980) );
  DFFX1_LVT u_T_427_reg_4__40_ ( .D(n4425), .CLK(n4258), .Q(n_T_427[1703]) );
  DFFX1_LVT u_T_427_reg_4__39_ ( .D(n4422), .CLK(n4258), .Q(n_T_427[1702]) );
  DFFX1_LVT u_T_427_reg_4__37_ ( .D(n4417), .CLK(n4258), .Q(n_T_427[1700]) );
  DFFX1_LVT u_T_427_reg_4__36_ ( .D(n4416), .CLK(n4258), .Q(n_T_427[1699]) );
  DFFX1_LVT u_T_427_reg_4__35_ ( .D(n4412), .CLK(n4257), .Q(n_T_427[1698]) );
  DFFX1_LVT u_T_427_reg_4__34_ ( .D(n4409), .CLK(n4257), .Q(n_T_427[1697]) );
  DFFX1_LVT u_T_427_reg_4__31_ ( .D(n4402), .CLK(n4257), .Q(n_T_427[1694]) );
  DFFX1_LVT u_T_427_reg_4__30_ ( .D(n4401), .CLK(n4257), .Q(n_T_427[1693]) );
  DFFX1_LVT u_T_427_reg_4__29_ ( .D(n4398), .CLK(n4257), .Q(n_T_427[1692]) );
  DFFX1_LVT u_T_427_reg_4__28_ ( .D(n4394), .CLK(n4257), .Q(n_T_427[1691]) );
  DFFX1_LVT u_T_427_reg_4__27_ ( .D(n4391), .CLK(n4257), .Q(n_T_427[1690]) );
  DFFX1_LVT u_T_427_reg_4__26_ ( .D(n4389), .CLK(n4257), .Q(n_T_427[1689]) );
  DFFX1_LVT u_T_427_reg_4__25_ ( .D(n4387), .CLK(n4257), .Q(n_T_427[1688]) );
  DFFX1_LVT u_T_427_reg_4__24_ ( .D(n4386), .CLK(n4257), .Q(n_T_427[1687]) );
  DFFX1_LVT u_T_427_reg_4__23_ ( .D(n4381), .CLK(n4256), .Q(n_T_427[1686]) );
  DFFX1_LVT u_T_427_reg_4__22_ ( .D(n4379), .CLK(n4256), .Q(n_T_427[1685]) );
  DFFX1_LVT u_T_427_reg_4__21_ ( .D(n4377), .CLK(n4256), .Q(n_T_427[1684]) );
  DFFX1_LVT u_T_427_reg_4__20_ ( .D(n4376), .CLK(n4256), .Q(n_T_427[1683]) );
  DFFX1_LVT u_T_427_reg_4__19_ ( .D(n4373), .CLK(n4256), .Q(n_T_427[1682]) );
  DFFX1_LVT u_T_427_reg_4__18_ ( .D(n4370), .CLK(n4256), .Q(n_T_427[1681]) );
  DFFX1_LVT u_T_427_reg_4__16_ ( .D(n4362), .CLK(n4256), .Q(n_T_427[1679]) );
  DFFX1_LVT u_T_427_reg_4__11_ ( .D(n4351), .CLK(n4255), .Q(n_T_427[1674]), 
        .QN(n3435) );
  DFFX1_LVT u_T_427_reg_4__1_ ( .D(n4321), .CLK(n4255), .Q(n_T_427[1664]) );
  DFFX1_LVT u_T_427_reg_4__0_ ( .D(n4318), .CLK(n4255), .Q(n_T_427[1663]) );
  DFFX1_LVT u_T_427_reg_5__63_ ( .D(n4494), .CLK(n4254), .Q(n_T_427[1662]) );
  DFFX1_LVT u_T_427_reg_5__62_ ( .D(n4491), .CLK(n4254), .Q(n_T_427[1661]) );
  DFFX1_LVT u_T_427_reg_5__61_ ( .D(n4488), .CLK(n4254), .Q(n_T_427[1660]) );
  DFFX1_LVT u_T_427_reg_5__60_ ( .D(n4485), .CLK(n4254), .Q(n_T_427[1659]) );
  DFFX1_LVT u_T_427_reg_5__59_ ( .D(n4482), .CLK(n4253), .Q(n_T_427[1658]) );
  DFFX1_LVT u_T_427_reg_5__58_ ( .D(n4481), .CLK(n4253), .Q(n_T_427[1657]) );
  DFFX1_LVT u_T_427_reg_5__57_ ( .D(n4476), .CLK(n4253), .Q(n_T_427[1656]) );
  DFFX1_LVT u_T_427_reg_5__56_ ( .D(n4475), .CLK(n4253), .Q(n_T_427[1655]) );
  DFFX1_LVT u_T_427_reg_5__55_ ( .D(n4470), .CLK(n4253), .Q(n_T_427[1654]) );
  DFFX1_LVT u_T_427_reg_5__54_ ( .D(n4469), .CLK(n4253), .Q(n_T_427[1653]) );
  DFFX1_LVT u_T_427_reg_5__53_ ( .D(n4464), .CLK(n4253), .Q(n_T_427[1652]) );
  DFFX1_LVT u_T_427_reg_5__52_ ( .D(n4463), .CLK(n4253), .Q(n_T_427[1651]) );
  DFFX1_LVT u_T_427_reg_5__51_ ( .D(n4460), .CLK(n4253), .Q(n_T_427[1650]) );
  DFFX1_LVT u_T_427_reg_5__50_ ( .D(n4455), .CLK(n4253), .Q(n_T_427[1649]) );
  DFFX1_LVT u_T_427_reg_5__49_ ( .D(n4454), .CLK(n4253), .Q(n_T_427[1648]) );
  DFFX1_LVT u_T_427_reg_5__48_ ( .D(n4449), .CLK(n4253), .Q(n_T_427[1647]) );
  DFFX1_LVT u_T_427_reg_5__47_ ( .D(n4446), .CLK(n4252), .Q(n_T_427[1646]) );
  DFFX1_LVT u_T_427_reg_5__46_ ( .D(n4443), .CLK(n4252), .Q(n_T_427[1645]) );
  DFFX1_LVT u_T_427_reg_5__45_ ( .D(n4442), .CLK(n4252), .Q(n_T_427[1644]) );
  DFFX1_LVT u_T_427_reg_5__44_ ( .D(n4437), .CLK(n4252), .Q(n_T_427[1643]) );
  DFFX1_LVT u_T_427_reg_5__43_ ( .D(n4436), .CLK(n4252), .Q(n_T_427[1642]) );
  DFFX1_LVT u_T_427_reg_5__42_ ( .D(n4433), .CLK(n4252), .Q(n_T_427[1641]) );
  DFFX1_LVT u_T_427_reg_5__41_ ( .D(n4430), .CLK(n4252), .Q(n_T_427[1640]) );
  DFFX1_LVT u_T_427_reg_5__40_ ( .D(n4425), .CLK(n4252), .Q(n_T_427[1639]) );
  DFFX1_LVT u_T_427_reg_5__39_ ( .D(n4422), .CLK(n4252), .Q(n_T_427[1638]) );
  DFFX1_LVT u_T_427_reg_5__38_ ( .D(n4420), .CLK(n4252), .Q(n_T_427[1637]) );
  DFFX1_LVT u_T_427_reg_5__37_ ( .D(n4417), .CLK(n4252), .Q(n_T_427[1636]) );
  DFFX1_LVT u_T_427_reg_5__36_ ( .D(n4416), .CLK(n4252), .Q(n_T_427[1635]) );
  DFFX1_LVT u_T_427_reg_5__35_ ( .D(n4412), .CLK(n4251), .Q(n_T_427[1634]) );
  DFFX1_LVT u_T_427_reg_5__34_ ( .D(n4409), .CLK(n4251), .Q(n_T_427[1633]) );
  DFFX1_LVT u_T_427_reg_5__33_ ( .D(n4407), .CLK(n4251), .Q(n_T_427[1632]) );
  DFFX1_LVT u_T_427_reg_5__32_ ( .D(n4404), .CLK(n4251), .Q(n_T_427[1631]) );
  DFFX1_LVT u_T_427_reg_5__31_ ( .D(n4402), .CLK(n4251), .Q(n_T_427[1630]) );
  DFFX1_LVT u_T_427_reg_5__30_ ( .D(n4401), .CLK(n4251), .Q(n_T_427[1629]) );
  DFFX1_LVT u_T_427_reg_5__29_ ( .D(n4398), .CLK(n4251), .Q(n_T_427[1628]) );
  DFFX1_LVT u_T_427_reg_5__28_ ( .D(n4394), .CLK(n4251), .Q(n_T_427[1627]) );
  DFFX1_LVT u_T_427_reg_5__27_ ( .D(n4391), .CLK(n4251), .Q(n_T_427[1626]) );
  DFFX1_LVT u_T_427_reg_5__26_ ( .D(n4389), .CLK(n4251), .Q(n_T_427[1625]) );
  DFFX1_LVT u_T_427_reg_5__25_ ( .D(n4387), .CLK(n4251), .Q(n_T_427[1624]) );
  DFFX1_LVT u_T_427_reg_5__24_ ( .D(n4386), .CLK(n4251), .Q(n_T_427[1623]) );
  DFFX1_LVT u_T_427_reg_5__23_ ( .D(n4381), .CLK(n4250), .Q(n_T_427[1622]) );
  DFFX1_LVT u_T_427_reg_5__22_ ( .D(n4379), .CLK(n4250), .Q(n_T_427[1621]) );
  DFFX1_LVT u_T_427_reg_5__21_ ( .D(n4377), .CLK(n4250), .Q(n_T_427[1620]) );
  DFFX1_LVT u_T_427_reg_5__20_ ( .D(n4376), .CLK(n4250), .Q(n_T_427[1619]) );
  DFFX1_LVT u_T_427_reg_5__19_ ( .D(n4373), .CLK(n4250), .Q(n_T_427[1618]) );
  DFFX1_LVT u_T_427_reg_5__18_ ( .D(n4370), .CLK(n4250), .Q(n_T_427[1617]) );
  DFFX1_LVT u_T_427_reg_5__17_ ( .D(n4365), .CLK(n4250), .Q(n_T_427[1616]) );
  DFFX1_LVT u_T_427_reg_5__16_ ( .D(n4362), .CLK(n4250), .Q(n_T_427[1615]) );
  DFFX1_LVT u_T_427_reg_5__15_ ( .D(n4360), .CLK(n4250), .Q(n_T_427[1614]) );
  DFFX1_LVT u_T_427_reg_5__14_ ( .D(n4357), .CLK(n4250), .Q(n_T_427[1613]) );
  DFFX1_LVT u_T_427_reg_5__13_ ( .D(n4355), .CLK(n4250), .Q(n_T_427[1612]) );
  DFFX1_LVT u_T_427_reg_5__12_ ( .D(n4352), .CLK(n4250), .Q(n_T_427[1611]) );
  DFFX1_LVT u_T_427_reg_5__11_ ( .D(n4351), .CLK(n4249), .Q(n_T_427[1610]) );
  DFFX1_LVT u_T_427_reg_5__10_ ( .D(n4346), .CLK(n4249), .Q(n_T_427[1609]) );
  DFFX1_LVT u_T_427_reg_5__9_ ( .D(n4343), .CLK(n4249), .Q(n_T_427[1608]) );
  DFFX1_LVT u_T_427_reg_5__8_ ( .D(n4340), .CLK(n4249), .Q(n_T_427[1607]) );
  DFFX1_LVT u_T_427_reg_5__7_ ( .D(n4337), .CLK(n4249), .Q(n_T_427[1606]) );
  DFFX1_LVT u_T_427_reg_5__6_ ( .D(n4334), .CLK(n4249), .Q(n_T_427[1605]) );
  DFFX1_LVT u_T_427_reg_5__5_ ( .D(n4331), .CLK(n4249), .Q(n_T_427[1604]) );
  DFFX1_LVT u_T_427_reg_5__4_ ( .D(n4328), .CLK(n4249), .Q(n_T_427[1603]) );
  DFFX1_LVT u_T_427_reg_5__3_ ( .D(n4325), .CLK(n4249), .Q(n_T_427[1602]) );
  DFFX1_LVT u_T_427_reg_5__2_ ( .D(n4322), .CLK(n4249), .Q(n_T_427[1601]) );
  DFFX1_LVT u_T_427_reg_5__1_ ( .D(n4321), .CLK(n4249), .Q(n_T_427[1600]) );
  DFFX1_LVT u_T_427_reg_5__0_ ( .D(n4318), .CLK(n4249), .Q(n_T_427[1599]) );
  DFFX1_LVT u_T_427_reg_6__63_ ( .D(n4494), .CLK(n4248), .Q(n_T_427[1598]) );
  DFFX1_LVT u_T_427_reg_6__62_ ( .D(n4491), .CLK(n4248), .Q(n_T_427[1597]) );
  DFFX1_LVT u_T_427_reg_6__61_ ( .D(n4488), .CLK(n4248), .Q(n_T_427[1596]) );
  DFFX1_LVT u_T_427_reg_6__60_ ( .D(n4485), .CLK(n4248), .Q(n_T_427[1595]) );
  DFFX1_LVT u_T_427_reg_6__59_ ( .D(n4482), .CLK(n4247), .Q(n_T_427[1594]) );
  DFFX1_LVT u_T_427_reg_6__58_ ( .D(n4481), .CLK(n4247), .Q(n_T_427[1593]) );
  DFFX1_LVT u_T_427_reg_6__57_ ( .D(n4476), .CLK(n4247), .Q(n_T_427[1592]) );
  DFFX1_LVT u_T_427_reg_6__56_ ( .D(n4475), .CLK(n4247), .Q(n_T_427[1591]) );
  DFFX1_LVT u_T_427_reg_6__55_ ( .D(n4470), .CLK(n4247), .Q(n_T_427[1590]) );
  DFFX1_LVT u_T_427_reg_6__54_ ( .D(n4469), .CLK(n4247), .Q(n_T_427[1589]) );
  DFFX1_LVT u_T_427_reg_6__53_ ( .D(n4464), .CLK(n4247), .Q(n_T_427[1588]) );
  DFFX1_LVT u_T_427_reg_6__52_ ( .D(n4463), .CLK(n4247), .Q(n_T_427[1587]) );
  DFFX1_LVT u_T_427_reg_6__51_ ( .D(n4460), .CLK(n4247), .Q(n_T_427[1586]) );
  DFFX1_LVT u_T_427_reg_6__50_ ( .D(n4455), .CLK(n4247), .Q(n_T_427[1585]) );
  DFFX1_LVT u_T_427_reg_6__49_ ( .D(n4454), .CLK(n4247), .Q(n_T_427[1584]) );
  DFFX1_LVT u_T_427_reg_6__48_ ( .D(n4449), .CLK(n4247), .Q(n_T_427[1583]) );
  DFFX1_LVT u_T_427_reg_6__47_ ( .D(n4446), .CLK(n4246), .Q(n_T_427[1582]) );
  DFFX1_LVT u_T_427_reg_6__46_ ( .D(n4443), .CLK(n4246), .Q(n_T_427[1581]) );
  DFFX1_LVT u_T_427_reg_6__45_ ( .D(n4442), .CLK(n4246), .Q(n_T_427[1580]) );
  DFFX1_LVT u_T_427_reg_6__44_ ( .D(n4437), .CLK(n4246), .Q(n_T_427[1579]) );
  DFFX1_LVT u_T_427_reg_6__43_ ( .D(n4436), .CLK(n4246), .Q(n_T_427[1578]) );
  DFFX1_LVT u_T_427_reg_6__42_ ( .D(n4433), .CLK(n4246), .Q(n_T_427[1577]) );
  DFFX1_LVT u_T_427_reg_6__41_ ( .D(n4430), .CLK(n4246), .Q(n_T_427[1576]) );
  DFFX1_LVT u_T_427_reg_6__40_ ( .D(n4425), .CLK(n4246), .Q(n_T_427[1575]) );
  DFFX1_LVT u_T_427_reg_6__39_ ( .D(n4422), .CLK(n4246), .Q(n_T_427[1574]) );
  DFFX1_LVT u_T_427_reg_6__38_ ( .D(n4420), .CLK(n4246), .Q(n_T_427[1573]) );
  DFFX1_LVT u_T_427_reg_6__37_ ( .D(n4417), .CLK(n4246), .Q(n_T_427[1572]) );
  DFFX1_LVT u_T_427_reg_6__36_ ( .D(n4416), .CLK(n4246), .Q(n_T_427[1571]) );
  DFFX1_LVT u_T_427_reg_6__35_ ( .D(n4412), .CLK(n4245), .Q(n_T_427[1570]) );
  DFFX1_LVT u_T_427_reg_6__34_ ( .D(n4409), .CLK(n4245), .Q(n_T_427[1569]) );
  DFFX1_LVT u_T_427_reg_6__33_ ( .D(n4407), .CLK(n4245), .Q(n_T_427[1568]) );
  DFFX1_LVT u_T_427_reg_6__32_ ( .D(n4404), .CLK(n4245), .Q(n_T_427[1567]) );
  DFFX1_LVT u_T_427_reg_6__31_ ( .D(n4402), .CLK(n4245), .Q(n_T_427[1566]) );
  DFFX1_LVT u_T_427_reg_6__30_ ( .D(n4401), .CLK(n4245), .Q(n_T_427[1565]) );
  DFFX1_LVT u_T_427_reg_6__29_ ( .D(n4398), .CLK(n4245), .Q(n_T_427[1564]) );
  DFFX1_LVT u_T_427_reg_6__28_ ( .D(n4394), .CLK(n4245), .Q(n_T_427[1563]) );
  DFFX1_LVT u_T_427_reg_6__27_ ( .D(n4391), .CLK(n4245), .Q(n_T_427[1562]) );
  DFFX1_LVT u_T_427_reg_6__26_ ( .D(n4389), .CLK(n4245), .Q(n_T_427[1561]) );
  DFFX1_LVT u_T_427_reg_6__25_ ( .D(n4387), .CLK(n4245), .Q(n_T_427[1560]) );
  DFFX1_LVT u_T_427_reg_6__24_ ( .D(n4386), .CLK(n4245), .Q(n_T_427[1559]) );
  DFFX1_LVT u_T_427_reg_6__23_ ( .D(n4381), .CLK(n4244), .Q(n_T_427[1558]) );
  DFFX1_LVT u_T_427_reg_6__22_ ( .D(n4379), .CLK(n4244), .Q(n_T_427[1557]) );
  DFFX1_LVT u_T_427_reg_6__21_ ( .D(n4377), .CLK(n4244), .Q(n_T_427[1556]) );
  DFFX1_LVT u_T_427_reg_6__20_ ( .D(n4376), .CLK(n4244), .Q(n_T_427[1555]) );
  DFFX1_LVT u_T_427_reg_6__19_ ( .D(n4373), .CLK(n4244), .Q(n_T_427[1554]) );
  DFFX1_LVT u_T_427_reg_6__18_ ( .D(n4370), .CLK(n4244), .Q(n_T_427[1553]) );
  DFFX1_LVT u_T_427_reg_6__17_ ( .D(n4365), .CLK(n4244), .Q(n_T_427[1552]) );
  DFFX1_LVT u_T_427_reg_6__16_ ( .D(n4362), .CLK(n4244), .Q(n_T_427[1551]) );
  DFFX1_LVT u_T_427_reg_6__15_ ( .D(n4360), .CLK(n4244), .Q(n_T_427[1550]) );
  DFFX1_LVT u_T_427_reg_6__14_ ( .D(n4357), .CLK(n4244), .Q(n_T_427[1549]) );
  DFFX1_LVT u_T_427_reg_6__13_ ( .D(n4355), .CLK(n4244), .Q(n_T_427[1548]) );
  DFFX1_LVT u_T_427_reg_6__12_ ( .D(n4352), .CLK(n4244), .Q(n_T_427[1547]) );
  DFFX1_LVT u_T_427_reg_6__11_ ( .D(n4351), .CLK(n4243), .Q(n_T_427[1546]) );
  DFFX1_LVT u_T_427_reg_6__10_ ( .D(n4346), .CLK(n4243), .Q(n_T_427[1545]) );
  DFFX1_LVT u_T_427_reg_6__9_ ( .D(n4343), .CLK(n4243), .Q(n_T_427[1544]) );
  DFFX1_LVT u_T_427_reg_6__8_ ( .D(n4340), .CLK(n4243), .Q(n_T_427[1543]) );
  DFFX1_LVT u_T_427_reg_6__7_ ( .D(n4337), .CLK(n4243), .Q(n_T_427[1542]) );
  DFFX1_LVT u_T_427_reg_6__6_ ( .D(n4334), .CLK(n4243), .Q(n_T_427[1541]) );
  DFFX1_LVT u_T_427_reg_6__5_ ( .D(n4331), .CLK(n4243), .Q(n_T_427[1540]) );
  DFFX1_LVT u_T_427_reg_6__4_ ( .D(n4328), .CLK(n4243), .Q(n_T_427[1539]) );
  DFFX1_LVT u_T_427_reg_6__3_ ( .D(n4325), .CLK(n4243), .Q(n_T_427[1538]) );
  DFFX1_LVT u_T_427_reg_6__2_ ( .D(n4322), .CLK(n4243), .Q(n_T_427[1537]) );
  DFFX1_LVT u_T_427_reg_6__1_ ( .D(n4321), .CLK(n4243), .Q(n_T_427[1536]) );
  DFFX1_LVT u_T_427_reg_6__0_ ( .D(n4318), .CLK(n4243), .Q(n_T_427[1535]) );
  DFFX1_LVT u_T_427_reg_7__63_ ( .D(n4494), .CLK(n4242), .Q(n_T_427[1534]) );
  DFFX1_LVT u_T_427_reg_7__62_ ( .D(n4491), .CLK(n4242), .Q(n_T_427[1533]) );
  DFFX1_LVT u_T_427_reg_7__61_ ( .D(n4488), .CLK(n4242), .Q(n_T_427[1532]) );
  DFFX1_LVT u_T_427_reg_7__60_ ( .D(n4485), .CLK(n4242), .Q(n_T_427[1531]) );
  DFFX1_LVT u_T_427_reg_7__59_ ( .D(n4482), .CLK(n4241), .Q(n_T_427[1530]) );
  DFFX1_LVT u_T_427_reg_7__58_ ( .D(n4481), .CLK(n4241), .Q(n_T_427[1529]) );
  DFFX1_LVT u_T_427_reg_7__57_ ( .D(n4476), .CLK(n4241), .Q(n_T_427[1528]) );
  DFFX1_LVT u_T_427_reg_7__56_ ( .D(n4475), .CLK(n4241), .Q(n_T_427[1527]) );
  DFFX1_LVT u_T_427_reg_7__55_ ( .D(n4470), .CLK(n4241), .Q(n_T_427[1526]) );
  DFFX1_LVT u_T_427_reg_7__54_ ( .D(n4469), .CLK(n4241), .Q(n_T_427[1525]) );
  DFFX1_LVT u_T_427_reg_7__53_ ( .D(n4464), .CLK(n4241), .Q(n_T_427[1524]) );
  DFFX1_LVT u_T_427_reg_7__52_ ( .D(n4463), .CLK(n4241), .Q(n_T_427[1523]) );
  DFFX1_LVT u_T_427_reg_7__51_ ( .D(n4460), .CLK(n4241), .Q(n_T_427[1522]) );
  DFFX1_LVT u_T_427_reg_7__50_ ( .D(n4455), .CLK(n4241), .Q(n_T_427[1521]) );
  DFFX1_LVT u_T_427_reg_7__49_ ( .D(n4454), .CLK(n4241), .Q(n_T_427[1520]) );
  DFFX1_LVT u_T_427_reg_7__48_ ( .D(n4449), .CLK(n4241), .Q(n_T_427[1519]), 
        .QN(n3774) );
  DFFX1_LVT u_T_427_reg_7__47_ ( .D(n4446), .CLK(n4240), .Q(n_T_427[1518]) );
  DFFX1_LVT u_T_427_reg_7__46_ ( .D(n4443), .CLK(n4240), .Q(n_T_427[1517]) );
  DFFX1_LVT u_T_427_reg_7__45_ ( .D(n4442), .CLK(n4240), .Q(n_T_427[1516]) );
  DFFX1_LVT u_T_427_reg_7__44_ ( .D(n4437), .CLK(n4240), .Q(n_T_427[1515]) );
  DFFX1_LVT u_T_427_reg_7__43_ ( .D(n4436), .CLK(n4240), .Q(n_T_427[1514]) );
  DFFX1_LVT u_T_427_reg_7__42_ ( .D(n4433), .CLK(n4240), .Q(n_T_427[1513]), 
        .QN(n3463) );
  DFFX1_LVT u_T_427_reg_7__41_ ( .D(n4430), .CLK(n4240), .Q(n_T_427[1512]) );
  DFFX1_LVT u_T_427_reg_7__40_ ( .D(n4425), .CLK(n4240), .Q(n_T_427[1511]) );
  DFFX1_LVT u_T_427_reg_7__37_ ( .D(n4417), .CLK(n4240), .Q(n_T_427[1508]) );
  DFFX1_LVT u_T_427_reg_7__36_ ( .D(n4416), .CLK(n4240), .Q(n_T_427[1507]), 
        .QN(n3455) );
  DFFX1_LVT u_T_427_reg_7__35_ ( .D(n4412), .CLK(n4239), .Q(n_T_427[1506]) );
  DFFX1_LVT u_T_427_reg_7__34_ ( .D(n4409), .CLK(n4239), .Q(n_T_427[1505]) );
  DFFX1_LVT u_T_427_reg_7__33_ ( .D(n4407), .CLK(n4239), .Q(n_T_427[1504]) );
  DFFX1_LVT u_T_427_reg_7__32_ ( .D(n4404), .CLK(n4239), .Q(n_T_427[1503]) );
  DFFX1_LVT u_T_427_reg_7__31_ ( .D(n4402), .CLK(n4239), .Q(n_T_427[1502]) );
  DFFX1_LVT u_T_427_reg_7__30_ ( .D(n4401), .CLK(n4239), .Q(n_T_427[1501]) );
  DFFX1_LVT u_T_427_reg_7__29_ ( .D(n4398), .CLK(n4239), .Q(n_T_427[1500]) );
  DFFX1_LVT u_T_427_reg_7__28_ ( .D(n4394), .CLK(n4239), .Q(n_T_427[1499]) );
  DFFX1_LVT u_T_427_reg_7__27_ ( .D(n4391), .CLK(n4239), .Q(n_T_427[1498]) );
  DFFX1_LVT u_T_427_reg_7__26_ ( .D(n4389), .CLK(n4239), .Q(n_T_427[1497]) );
  DFFX1_LVT u_T_427_reg_7__25_ ( .D(n4387), .CLK(n4239), .Q(n_T_427[1496]) );
  DFFX1_LVT u_T_427_reg_7__24_ ( .D(n4386), .CLK(n4239), .Q(n_T_427[1495]) );
  DFFX1_LVT u_T_427_reg_7__23_ ( .D(n4381), .CLK(n4238), .Q(n_T_427[1494]) );
  DFFX1_LVT u_T_427_reg_7__22_ ( .D(n4379), .CLK(n4238), .Q(n_T_427[1493]) );
  DFFX1_LVT u_T_427_reg_7__21_ ( .D(n4377), .CLK(n4238), .Q(n_T_427[1492]) );
  DFFX1_LVT u_T_427_reg_7__20_ ( .D(n4376), .CLK(n4238), .Q(n_T_427[1491]) );
  DFFX1_LVT u_T_427_reg_7__19_ ( .D(n4373), .CLK(n4238), .Q(n_T_427[1490]) );
  DFFX1_LVT u_T_427_reg_7__18_ ( .D(n4370), .CLK(n4238), .Q(n_T_427[1489]) );
  DFFX1_LVT u_T_427_reg_7__17_ ( .D(n4365), .CLK(n4238), .Q(n_T_427[1488]) );
  DFFX1_LVT u_T_427_reg_7__16_ ( .D(n4362), .CLK(n4238), .Q(n_T_427[1487]) );
  DFFX1_LVT u_T_427_reg_7__1_ ( .D(n4321), .CLK(n4237), .Q(n_T_427[1472]), 
        .QN(n3416) );
  DFFX1_LVT u_T_427_reg_7__0_ ( .D(n4318), .CLK(n4237), .Q(n_T_427[1471]), 
        .QN(n3417) );
  DFFX1_LVT u_T_427_reg_8__63_ ( .D(n4494), .CLK(n4236), .Q(n_T_427[1470]) );
  DFFX1_LVT u_T_427_reg_8__62_ ( .D(n4491), .CLK(n4236), .Q(n_T_427[1469]) );
  DFFX1_LVT u_T_427_reg_8__61_ ( .D(n4488), .CLK(n4236), .Q(n_T_427[1468]) );
  DFFX1_LVT u_T_427_reg_8__60_ ( .D(n4485), .CLK(n4236), .Q(n_T_427[1467]) );
  DFFX1_LVT u_T_427_reg_8__59_ ( .D(n4482), .CLK(n4235), .Q(n_T_427[1466]) );
  DFFX1_LVT u_T_427_reg_8__58_ ( .D(n4480), .CLK(n4235), .Q(n_T_427[1465]) );
  DFFX1_LVT u_T_427_reg_8__57_ ( .D(n4476), .CLK(n4235), .Q(n_T_427[1464]) );
  DFFX1_LVT u_T_427_reg_8__56_ ( .D(n4474), .CLK(n4235), .Q(n_T_427[1463]) );
  DFFX1_LVT u_T_427_reg_8__55_ ( .D(n4470), .CLK(n4235), .Q(n_T_427[1462]) );
  DFFX1_LVT u_T_427_reg_8__54_ ( .D(n4468), .CLK(n4235), .Q(n_T_427[1461]) );
  DFFX1_LVT u_T_427_reg_8__53_ ( .D(n4464), .CLK(n4235), .Q(n_T_427[1460]) );
  DFFX1_LVT u_T_427_reg_8__52_ ( .D(n4462), .CLK(n4235), .Q(n_T_427[1459]) );
  DFFX1_LVT u_T_427_reg_8__51_ ( .D(n4459), .CLK(n4235), .Q(n_T_427[1458]) );
  DFFX1_LVT u_T_427_reg_8__50_ ( .D(n4455), .CLK(n4235), .Q(n_T_427[1457]) );
  DFFX1_LVT u_T_427_reg_8__49_ ( .D(n4453), .CLK(n4235), .Q(n_T_427[1456]) );
  DFFX1_LVT u_T_427_reg_8__48_ ( .D(n4449), .CLK(n4235), .Q(n_T_427[1455]) );
  DFFX1_LVT u_T_427_reg_8__47_ ( .D(n4446), .CLK(n4234), .Q(n_T_427[1454]) );
  DFFX1_LVT u_T_427_reg_8__46_ ( .D(n4443), .CLK(n4234), .Q(n_T_427[1453]) );
  DFFX1_LVT u_T_427_reg_8__45_ ( .D(n4441), .CLK(n4234), .Q(n_T_427[1452]) );
  DFFX1_LVT u_T_427_reg_8__44_ ( .D(n4437), .CLK(n4234), .Q(n_T_427[1451]) );
  DFFX1_LVT u_T_427_reg_8__43_ ( .D(n4435), .CLK(n4234), .Q(n_T_427[1450]) );
  DFFX1_LVT u_T_427_reg_8__42_ ( .D(n4432), .CLK(n4234), .Q(n_T_427[1449]) );
  DFFX1_LVT u_T_427_reg_8__41_ ( .D(n4429), .CLK(n4234), .Q(n_T_427[1448]) );
  DFFX1_LVT u_T_427_reg_8__40_ ( .D(n4425), .CLK(n4234), .Q(n_T_427[1447]) );
  DFFX1_LVT u_T_427_reg_8__39_ ( .D(n4422), .CLK(n4234), .Q(n_T_427[1446]) );
  DFFX1_LVT u_T_427_reg_8__38_ ( .D(n4420), .CLK(n4234), .Q(n_T_427[1445]) );
  DFFX1_LVT u_T_427_reg_8__37_ ( .D(n4417), .CLK(n4234), .Q(n_T_427[1444]) );
  DFFX1_LVT u_T_427_reg_8__36_ ( .D(n4415), .CLK(n4234), .Q(n_T_427[1443]) );
  DFFX1_LVT u_T_427_reg_8__35_ ( .D(n4412), .CLK(n4233), .Q(n_T_427[1442]) );
  DFFX1_LVT u_T_427_reg_8__34_ ( .D(n4409), .CLK(n4233), .Q(n_T_427[1441]) );
  DFFX1_LVT u_T_427_reg_8__33_ ( .D(n4407), .CLK(n4233), .Q(n_T_427[1440]) );
  DFFX1_LVT u_T_427_reg_8__32_ ( .D(n4404), .CLK(n4233), .Q(n_T_427[1439]) );
  DFFX1_LVT u_T_427_reg_8__31_ ( .D(n4402), .CLK(n4233), .Q(n_T_427[1438]) );
  DFFX1_LVT u_T_427_reg_8__30_ ( .D(n4400), .CLK(n4233), .Q(n_T_427[1437]) );
  DFFX1_LVT u_T_427_reg_8__29_ ( .D(n4397), .CLK(n4233), .Q(n_T_427[1436]) );
  DFFX1_LVT u_T_427_reg_8__28_ ( .D(n4394), .CLK(n4233), .Q(n_T_427[1435]) );
  DFFX1_LVT u_T_427_reg_8__27_ ( .D(n4391), .CLK(n4233), .Q(n_T_427[1434]) );
  DFFX1_LVT u_T_427_reg_8__26_ ( .D(n4389), .CLK(n4233), .Q(n_T_427[1433]) );
  DFFX1_LVT u_T_427_reg_8__25_ ( .D(n4387), .CLK(n4233), .Q(n_T_427[1432]) );
  DFFX1_LVT u_T_427_reg_8__24_ ( .D(n4385), .CLK(n4233), .Q(n_T_427[1431]) );
  DFFX1_LVT u_T_427_reg_8__23_ ( .D(n4381), .CLK(n4232), .Q(n_T_427[1430]) );
  DFFX1_LVT u_T_427_reg_8__22_ ( .D(n4379), .CLK(n4232), .Q(n_T_427[1429]) );
  DFFX1_LVT u_T_427_reg_8__21_ ( .D(n4377), .CLK(n4232), .Q(n_T_427[1428]) );
  DFFX1_LVT u_T_427_reg_8__20_ ( .D(n4375), .CLK(n4232), .Q(n_T_427[1427]) );
  DFFX1_LVT u_T_427_reg_8__19_ ( .D(n4372), .CLK(n4232), .Q(n_T_427[1426]) );
  DFFX1_LVT u_T_427_reg_8__18_ ( .D(n4369), .CLK(n4232), .Q(n_T_427[1425]) );
  DFFX1_LVT u_T_427_reg_8__17_ ( .D(n4365), .CLK(n4232), .Q(n_T_427[1424]) );
  DFFX1_LVT u_T_427_reg_8__16_ ( .D(n4362), .CLK(n4232), .Q(n_T_427[1423]) );
  DFFX1_LVT u_T_427_reg_8__15_ ( .D(n4360), .CLK(n4232), .Q(n_T_427[1422]) );
  DFFX1_LVT u_T_427_reg_8__14_ ( .D(n4357), .CLK(n4232), .Q(n_T_427[1421]) );
  DFFX1_LVT u_T_427_reg_8__13_ ( .D(n4355), .CLK(n4232), .Q(n_T_427[1420]) );
  DFFX1_LVT u_T_427_reg_8__12_ ( .D(n4352), .CLK(n4232), .Q(n_T_427[1419]) );
  DFFX1_LVT u_T_427_reg_8__11_ ( .D(n4350), .CLK(n4231), .Q(n_T_427[1418]) );
  DFFX1_LVT u_T_427_reg_8__10_ ( .D(n4346), .CLK(n4231), .Q(n_T_427[1417]) );
  DFFX1_LVT u_T_427_reg_8__9_ ( .D(n4343), .CLK(n4231), .Q(n_T_427[1416]) );
  DFFX1_LVT u_T_427_reg_8__8_ ( .D(n4340), .CLK(n4231), .Q(n_T_427[1415]) );
  DFFX1_LVT u_T_427_reg_8__7_ ( .D(n4337), .CLK(n4231), .Q(n_T_427[1414]) );
  DFFX1_LVT u_T_427_reg_8__6_ ( .D(n4334), .CLK(n4231), .Q(n_T_427[1413]) );
  DFFX1_LVT u_T_427_reg_8__5_ ( .D(n4331), .CLK(n4231), .Q(n_T_427[1412]) );
  DFFX1_LVT u_T_427_reg_8__4_ ( .D(n4328), .CLK(n4231), .Q(n_T_427[1411]) );
  DFFX1_LVT u_T_427_reg_8__3_ ( .D(n4325), .CLK(n4231), .Q(n_T_427[1410]) );
  DFFX1_LVT u_T_427_reg_8__2_ ( .D(n4322), .CLK(n4231), .Q(n_T_427[1409]) );
  DFFX1_LVT u_T_427_reg_8__1_ ( .D(n4320), .CLK(n4231), .Q(n_T_427[1408]) );
  DFFX1_LVT u_T_427_reg_8__0_ ( .D(n4317), .CLK(n4231), .Q(n_T_427[1407]) );
  DFFX1_LVT u_T_427_reg_9__63_ ( .D(n4494), .CLK(n4230), .Q(n_T_427[1406]) );
  DFFX1_LVT u_T_427_reg_9__62_ ( .D(n4491), .CLK(n4230), .Q(n_T_427[1405]) );
  DFFX1_LVT u_T_427_reg_9__61_ ( .D(n4488), .CLK(n4230), .Q(n_T_427[1404]) );
  DFFX1_LVT u_T_427_reg_9__60_ ( .D(n4485), .CLK(n4230), .Q(n_T_427[1403]) );
  DFFX1_LVT u_T_427_reg_9__59_ ( .D(n4482), .CLK(n4229), .Q(n_T_427[1402]) );
  DFFX1_LVT u_T_427_reg_9__58_ ( .D(n4480), .CLK(n4229), .Q(n_T_427[1401]) );
  DFFX1_LVT u_T_427_reg_9__57_ ( .D(n4476), .CLK(n4229), .Q(n_T_427[1400]) );
  DFFX1_LVT u_T_427_reg_9__56_ ( .D(n4474), .CLK(n4229), .Q(n_T_427[1399]) );
  DFFX1_LVT u_T_427_reg_9__55_ ( .D(n4470), .CLK(n4229), .Q(n_T_427[1398]) );
  DFFX1_LVT u_T_427_reg_9__54_ ( .D(n4468), .CLK(n4229), .Q(n_T_427[1397]) );
  DFFX1_LVT u_T_427_reg_9__53_ ( .D(n4464), .CLK(n4229), .Q(n_T_427[1396]) );
  DFFX1_LVT u_T_427_reg_9__52_ ( .D(n4462), .CLK(n4229), .Q(n_T_427[1395]) );
  DFFX1_LVT u_T_427_reg_9__51_ ( .D(n4459), .CLK(n4229), .Q(n_T_427[1394]) );
  DFFX1_LVT u_T_427_reg_9__50_ ( .D(n4455), .CLK(n4229), .Q(n_T_427[1393]) );
  DFFX1_LVT u_T_427_reg_9__49_ ( .D(n4453), .CLK(n4229), .Q(n_T_427[1392]) );
  DFFX1_LVT u_T_427_reg_9__48_ ( .D(n4449), .CLK(n4229), .Q(n_T_427[1391]) );
  DFFX1_LVT u_T_427_reg_9__47_ ( .D(n4446), .CLK(n4228), .Q(n_T_427[1390]) );
  DFFX1_LVT u_T_427_reg_9__46_ ( .D(n4443), .CLK(n4228), .Q(n_T_427[1389]) );
  DFFX1_LVT u_T_427_reg_9__45_ ( .D(n4441), .CLK(n4228), .Q(n_T_427[1388]) );
  DFFX1_LVT u_T_427_reg_9__44_ ( .D(n4437), .CLK(n4228), .Q(n_T_427[1387]) );
  DFFX1_LVT u_T_427_reg_9__43_ ( .D(n4435), .CLK(n4228), .Q(n_T_427[1386]) );
  DFFX1_LVT u_T_427_reg_9__42_ ( .D(n4432), .CLK(n4228), .Q(n_T_427[1385]) );
  DFFX1_LVT u_T_427_reg_9__41_ ( .D(n4429), .CLK(n4228), .Q(n_T_427[1384]) );
  DFFX1_LVT u_T_427_reg_9__40_ ( .D(n4425), .CLK(n4228), .Q(n_T_427[1383]) );
  DFFX1_LVT u_T_427_reg_9__39_ ( .D(n4422), .CLK(n4228), .Q(n_T_427[1382]) );
  DFFX1_LVT u_T_427_reg_9__38_ ( .D(n4420), .CLK(n4228), .Q(n_T_427[1381]) );
  DFFX1_LVT u_T_427_reg_9__37_ ( .D(n4417), .CLK(n4228), .Q(n_T_427[1380]) );
  DFFX1_LVT u_T_427_reg_9__36_ ( .D(n4415), .CLK(n4228), .Q(n_T_427[1379]) );
  DFFX1_LVT u_T_427_reg_9__35_ ( .D(n4412), .CLK(n4227), .Q(n_T_427[1378]) );
  DFFX1_LVT u_T_427_reg_9__34_ ( .D(n4409), .CLK(n4227), .Q(n_T_427[1377]) );
  DFFX1_LVT u_T_427_reg_9__33_ ( .D(n4407), .CLK(n4227), .Q(n_T_427[1376]) );
  DFFX1_LVT u_T_427_reg_9__32_ ( .D(n4404), .CLK(n4227), .Q(n_T_427[1375]) );
  DFFX1_LVT u_T_427_reg_9__31_ ( .D(n4402), .CLK(n4227), .Q(n_T_427[1374]) );
  DFFX1_LVT u_T_427_reg_9__30_ ( .D(n4400), .CLK(n4227), .Q(n_T_427[1373]) );
  DFFX1_LVT u_T_427_reg_9__29_ ( .D(n4397), .CLK(n4227), .Q(n_T_427[1372]) );
  DFFX1_LVT u_T_427_reg_9__28_ ( .D(n4394), .CLK(n4227), .Q(n_T_427[1371]) );
  DFFX1_LVT u_T_427_reg_9__27_ ( .D(n4391), .CLK(n4227), .Q(n_T_427[1370]) );
  DFFX1_LVT u_T_427_reg_9__26_ ( .D(n4389), .CLK(n4227), .Q(n_T_427[1369]) );
  DFFX1_LVT u_T_427_reg_9__25_ ( .D(n4387), .CLK(n4227), .Q(n_T_427[1368]) );
  DFFX1_LVT u_T_427_reg_9__24_ ( .D(n4385), .CLK(n4227), .Q(n_T_427[1367]) );
  DFFX1_LVT u_T_427_reg_9__23_ ( .D(n4381), .CLK(n4226), .Q(n_T_427[1366]) );
  DFFX1_LVT u_T_427_reg_9__22_ ( .D(n4379), .CLK(n4226), .Q(n_T_427[1365]) );
  DFFX1_LVT u_T_427_reg_9__21_ ( .D(n4377), .CLK(n4226), .Q(n_T_427[1364]) );
  DFFX1_LVT u_T_427_reg_9__20_ ( .D(n4375), .CLK(n4226), .Q(n_T_427[1363]) );
  DFFX1_LVT u_T_427_reg_9__19_ ( .D(n4372), .CLK(n4226), .Q(n_T_427[1362]) );
  DFFX1_LVT u_T_427_reg_9__18_ ( .D(n4369), .CLK(n4226), .Q(n_T_427[1361]) );
  DFFX1_LVT u_T_427_reg_9__17_ ( .D(n4365), .CLK(n4226), .Q(n_T_427[1360]) );
  DFFX1_LVT u_T_427_reg_9__16_ ( .D(n4362), .CLK(n4226), .Q(n_T_427[1359]) );
  DFFX1_LVT u_T_427_reg_9__15_ ( .D(n4360), .CLK(n4226), .Q(n_T_427[1358]) );
  DFFX1_LVT u_T_427_reg_9__14_ ( .D(n4357), .CLK(n4226), .Q(n_T_427[1357]) );
  DFFX1_LVT u_T_427_reg_9__13_ ( .D(n4355), .CLK(n4226), .Q(n_T_427[1356]) );
  DFFX1_LVT u_T_427_reg_9__12_ ( .D(n4352), .CLK(n4226), .Q(n_T_427[1355]) );
  DFFX1_LVT u_T_427_reg_9__11_ ( .D(n4350), .CLK(n4225), .Q(n_T_427[1354]) );
  DFFX1_LVT u_T_427_reg_9__10_ ( .D(n4346), .CLK(n4225), .Q(n_T_427[1353]) );
  DFFX1_LVT u_T_427_reg_9__9_ ( .D(n4343), .CLK(n4225), .Q(n_T_427[1352]) );
  DFFX1_LVT u_T_427_reg_9__8_ ( .D(n4340), .CLK(n4225), .Q(n_T_427[1351]) );
  DFFX1_LVT u_T_427_reg_9__7_ ( .D(n4337), .CLK(n4225), .Q(n_T_427[1350]) );
  DFFX1_LVT u_T_427_reg_9__6_ ( .D(n4334), .CLK(n4225), .Q(n_T_427[1349]) );
  DFFX1_LVT u_T_427_reg_9__5_ ( .D(n4331), .CLK(n4225), .Q(n_T_427[1348]) );
  DFFX1_LVT u_T_427_reg_9__4_ ( .D(n4328), .CLK(n4225), .Q(n_T_427[1347]) );
  DFFX1_LVT u_T_427_reg_9__3_ ( .D(n4325), .CLK(n4225), .Q(n_T_427[1346]) );
  DFFX1_LVT u_T_427_reg_9__2_ ( .D(n4322), .CLK(n4225), .Q(n_T_427[1345]) );
  DFFX1_LVT u_T_427_reg_9__1_ ( .D(n4320), .CLK(n4225), .Q(n_T_427[1344]) );
  DFFX1_LVT u_T_427_reg_9__0_ ( .D(n4317), .CLK(n4225), .Q(n_T_427[1343]) );
  DFFX1_LVT u_T_427_reg_10__63_ ( .D(n4494), .CLK(n4224), .Q(n_T_427[1342]) );
  DFFX1_LVT u_T_427_reg_10__62_ ( .D(n4491), .CLK(n4224), .Q(n_T_427[1341]) );
  DFFX1_LVT u_T_427_reg_10__61_ ( .D(n4488), .CLK(n4224), .Q(n_T_427[1340]) );
  DFFX1_LVT u_T_427_reg_10__60_ ( .D(n4485), .CLK(n4224), .Q(n_T_427[1339]) );
  DFFX1_LVT u_T_427_reg_10__59_ ( .D(n4482), .CLK(n4223), .Q(n_T_427[1338]) );
  DFFX1_LVT u_T_427_reg_10__58_ ( .D(n4480), .CLK(n4223), .Q(n_T_427[1337]) );
  DFFX1_LVT u_T_427_reg_10__57_ ( .D(n4476), .CLK(n4223), .Q(n_T_427[1336]) );
  DFFX1_LVT u_T_427_reg_10__56_ ( .D(n4474), .CLK(n4223), .Q(n_T_427[1335]) );
  DFFX1_LVT u_T_427_reg_10__55_ ( .D(n4470), .CLK(n4223), .Q(n_T_427[1334]) );
  DFFX1_LVT u_T_427_reg_10__54_ ( .D(n4468), .CLK(n4223), .Q(n_T_427[1333]) );
  DFFX1_LVT u_T_427_reg_10__53_ ( .D(n4464), .CLK(n4223), .Q(n_T_427[1332]) );
  DFFX1_LVT u_T_427_reg_10__52_ ( .D(n4462), .CLK(n4223), .Q(n_T_427[1331]) );
  DFFX1_LVT u_T_427_reg_10__51_ ( .D(n4459), .CLK(n4223), .Q(n_T_427[1330]) );
  DFFX1_LVT u_T_427_reg_10__50_ ( .D(n4455), .CLK(n4223), .Q(n_T_427[1329]) );
  DFFX1_LVT u_T_427_reg_10__49_ ( .D(n4453), .CLK(n4223), .Q(n_T_427[1328]) );
  DFFX1_LVT u_T_427_reg_10__48_ ( .D(n4449), .CLK(n4223), .Q(n_T_427[1327]) );
  DFFX1_LVT u_T_427_reg_10__47_ ( .D(n4446), .CLK(n4222), .Q(n_T_427[1326]) );
  DFFX1_LVT u_T_427_reg_10__46_ ( .D(n4443), .CLK(n4222), .Q(n_T_427[1325]) );
  DFFX1_LVT u_T_427_reg_10__45_ ( .D(n4441), .CLK(n4222), .Q(n_T_427[1324]) );
  DFFX1_LVT u_T_427_reg_10__44_ ( .D(n4437), .CLK(n4222), .Q(n_T_427[1323]) );
  DFFX1_LVT u_T_427_reg_10__43_ ( .D(n4435), .CLK(n4222), .Q(n_T_427[1322]) );
  DFFX1_LVT u_T_427_reg_10__42_ ( .D(n4432), .CLK(n4222), .Q(n_T_427[1321]) );
  DFFX1_LVT u_T_427_reg_10__41_ ( .D(n4429), .CLK(n4222), .Q(n_T_427[1320]) );
  DFFX1_LVT u_T_427_reg_10__40_ ( .D(n4425), .CLK(n4222), .Q(n_T_427[1319]) );
  DFFX1_LVT u_T_427_reg_10__39_ ( .D(n4422), .CLK(n4222), .Q(n_T_427[1318]) );
  DFFX1_LVT u_T_427_reg_10__38_ ( .D(n4420), .CLK(n4222), .Q(n_T_427[1317]) );
  DFFX1_LVT u_T_427_reg_10__37_ ( .D(n4417), .CLK(n4222), .Q(n_T_427[1316]) );
  DFFX1_LVT u_T_427_reg_10__36_ ( .D(n4415), .CLK(n4222), .Q(n_T_427[1315]) );
  DFFX1_LVT u_T_427_reg_10__35_ ( .D(n4412), .CLK(n4221), .Q(n_T_427[1314]) );
  DFFX1_LVT u_T_427_reg_10__34_ ( .D(n4409), .CLK(n4221), .Q(n_T_427[1313]) );
  DFFX1_LVT u_T_427_reg_10__33_ ( .D(n4407), .CLK(n4221), .Q(n_T_427[1312]) );
  DFFX1_LVT u_T_427_reg_10__32_ ( .D(n4404), .CLK(n4221), .Q(n_T_427[1311]) );
  DFFX1_LVT u_T_427_reg_10__31_ ( .D(n4402), .CLK(n4221), .Q(n_T_427[1310]) );
  DFFX1_LVT u_T_427_reg_10__30_ ( .D(n4400), .CLK(n4221), .Q(n_T_427[1309]) );
  DFFX1_LVT u_T_427_reg_10__29_ ( .D(n4397), .CLK(n4221), .Q(n_T_427[1308]) );
  DFFX1_LVT u_T_427_reg_10__28_ ( .D(n4394), .CLK(n4221), .Q(n_T_427[1307]) );
  DFFX1_LVT u_T_427_reg_10__27_ ( .D(n4391), .CLK(n4221), .Q(n_T_427[1306]) );
  DFFX1_LVT u_T_427_reg_10__26_ ( .D(n4389), .CLK(n4221), .Q(n_T_427[1305]) );
  DFFX1_LVT u_T_427_reg_10__25_ ( .D(n4387), .CLK(n4221), .Q(n_T_427[1304]) );
  DFFX1_LVT u_T_427_reg_10__24_ ( .D(n4385), .CLK(n4221), .Q(n_T_427[1303]) );
  DFFX1_LVT u_T_427_reg_10__23_ ( .D(n4381), .CLK(n4220), .Q(n_T_427[1302]) );
  DFFX1_LVT u_T_427_reg_10__22_ ( .D(n4379), .CLK(n4220), .Q(n_T_427[1301]) );
  DFFX1_LVT u_T_427_reg_10__21_ ( .D(n4377), .CLK(n4220), .Q(n_T_427[1300]) );
  DFFX1_LVT u_T_427_reg_10__20_ ( .D(n4375), .CLK(n4220), .Q(n_T_427[1299]) );
  DFFX1_LVT u_T_427_reg_10__19_ ( .D(n4372), .CLK(n4220), .Q(n_T_427[1298]) );
  DFFX1_LVT u_T_427_reg_10__18_ ( .D(n4369), .CLK(n4220), .Q(n_T_427[1297]) );
  DFFX1_LVT u_T_427_reg_10__17_ ( .D(n4365), .CLK(n4220), .Q(n_T_427[1296]) );
  DFFX1_LVT u_T_427_reg_10__16_ ( .D(n4362), .CLK(n4220), .Q(n_T_427[1295]) );
  DFFX1_LVT u_T_427_reg_10__15_ ( .D(n4360), .CLK(n4220), .Q(n_T_427[1294]) );
  DFFX1_LVT u_T_427_reg_10__14_ ( .D(n4357), .CLK(n4220), .Q(n_T_427[1293]) );
  DFFX1_LVT u_T_427_reg_10__13_ ( .D(n4355), .CLK(n4220), .Q(n_T_427[1292]) );
  DFFX1_LVT u_T_427_reg_10__12_ ( .D(n4352), .CLK(n4220), .Q(n_T_427[1291]) );
  DFFX1_LVT u_T_427_reg_10__11_ ( .D(n4350), .CLK(n4219), .Q(n_T_427[1290]) );
  DFFX1_LVT u_T_427_reg_10__10_ ( .D(n4346), .CLK(n4219), .Q(n_T_427[1289]) );
  DFFX1_LVT u_T_427_reg_10__9_ ( .D(n4343), .CLK(n4219), .Q(n_T_427[1288]) );
  DFFX1_LVT u_T_427_reg_10__8_ ( .D(n4340), .CLK(n4219), .Q(n_T_427[1287]) );
  DFFX1_LVT u_T_427_reg_10__7_ ( .D(n4337), .CLK(n4219), .Q(n_T_427[1286]) );
  DFFX1_LVT u_T_427_reg_10__6_ ( .D(n4334), .CLK(n4219), .Q(n_T_427[1285]) );
  DFFX1_LVT u_T_427_reg_10__5_ ( .D(n4331), .CLK(n4219), .Q(n_T_427[1284]) );
  DFFX1_LVT u_T_427_reg_10__4_ ( .D(n4328), .CLK(n4219), .Q(n_T_427[1283]) );
  DFFX1_LVT u_T_427_reg_10__3_ ( .D(n4325), .CLK(n4219), .Q(n_T_427[1282]) );
  DFFX1_LVT u_T_427_reg_10__2_ ( .D(n4322), .CLK(n4219), .Q(n_T_427[1281]) );
  DFFX1_LVT u_T_427_reg_10__1_ ( .D(n4320), .CLK(n4219), .Q(n_T_427[1280]) );
  DFFX1_LVT u_T_427_reg_10__0_ ( .D(n4317), .CLK(n4219), .Q(n_T_427[1279]) );
  DFFX1_LVT u_T_427_reg_11__63_ ( .D(n4494), .CLK(n4218), .Q(n_T_427[1278]) );
  DFFX1_LVT u_T_427_reg_11__62_ ( .D(n4491), .CLK(n4218), .Q(n_T_427[1277]) );
  DFFX1_LVT u_T_427_reg_11__61_ ( .D(n4488), .CLK(n4218), .Q(n_T_427[1276]) );
  DFFX1_LVT u_T_427_reg_11__60_ ( .D(n4485), .CLK(n4218), .Q(n_T_427[1275]) );
  DFFX1_LVT u_T_427_reg_11__59_ ( .D(n4482), .CLK(n4217), .Q(n_T_427[1274]) );
  DFFX1_LVT u_T_427_reg_11__58_ ( .D(n4480), .CLK(n4217), .Q(n_T_427[1273]) );
  DFFX1_LVT u_T_427_reg_11__57_ ( .D(n4476), .CLK(n4217), .Q(n_T_427[1272]) );
  DFFX1_LVT u_T_427_reg_11__56_ ( .D(n4474), .CLK(n4217), .Q(n_T_427[1271]) );
  DFFX1_LVT u_T_427_reg_11__55_ ( .D(n4470), .CLK(n4217), .Q(n_T_427[1270]) );
  DFFX1_LVT u_T_427_reg_11__54_ ( .D(n4468), .CLK(n4217), .Q(n_T_427[1269]) );
  DFFX1_LVT u_T_427_reg_11__53_ ( .D(n4464), .CLK(n4217), .Q(n_T_427[1268]) );
  DFFX1_LVT u_T_427_reg_11__52_ ( .D(n4462), .CLK(n4217), .Q(n_T_427[1267]) );
  DFFX1_LVT u_T_427_reg_11__51_ ( .D(n4459), .CLK(n4217), .Q(n_T_427[1266]) );
  DFFX1_LVT u_T_427_reg_11__50_ ( .D(n4455), .CLK(n4217), .Q(n_T_427[1265]) );
  DFFX1_LVT u_T_427_reg_11__49_ ( .D(n4453), .CLK(n4217), .Q(n_T_427[1264]) );
  DFFX1_LVT u_T_427_reg_11__48_ ( .D(n4449), .CLK(n4217), .Q(n_T_427[1263]) );
  DFFX1_LVT u_T_427_reg_11__47_ ( .D(n4446), .CLK(n4216), .Q(n_T_427[1262]) );
  DFFX1_LVT u_T_427_reg_11__46_ ( .D(n4443), .CLK(n4216), .Q(n_T_427[1261]) );
  DFFX1_LVT u_T_427_reg_11__45_ ( .D(n4441), .CLK(n4216), .Q(n_T_427[1260]) );
  DFFX1_LVT u_T_427_reg_11__44_ ( .D(n4437), .CLK(n4216), .Q(n_T_427[1259]) );
  DFFX1_LVT u_T_427_reg_11__43_ ( .D(n4435), .CLK(n4216), .Q(n_T_427[1258]) );
  DFFX1_LVT u_T_427_reg_11__42_ ( .D(n4432), .CLK(n4216), .Q(n_T_427[1257]) );
  DFFX1_LVT u_T_427_reg_11__41_ ( .D(n4429), .CLK(n4216), .Q(n_T_427[1256]) );
  DFFX1_LVT u_T_427_reg_11__40_ ( .D(n4425), .CLK(n4216), .Q(n_T_427[1255]) );
  DFFX1_LVT u_T_427_reg_11__39_ ( .D(n4422), .CLK(n4216), .Q(n_T_427[1254]) );
  DFFX1_LVT u_T_427_reg_11__38_ ( .D(n4420), .CLK(n4216), .Q(n_T_427[1253]) );
  DFFX1_LVT u_T_427_reg_11__37_ ( .D(n4417), .CLK(n4216), .Q(n_T_427[1252]) );
  DFFX1_LVT u_T_427_reg_11__36_ ( .D(n4415), .CLK(n4216), .Q(n_T_427[1251]) );
  DFFX1_LVT u_T_427_reg_11__35_ ( .D(n4412), .CLK(n4215), .Q(n_T_427[1250]) );
  DFFX1_LVT u_T_427_reg_11__34_ ( .D(n4409), .CLK(n4215), .Q(n_T_427[1249]) );
  DFFX1_LVT u_T_427_reg_11__33_ ( .D(n4407), .CLK(n4215), .Q(n_T_427[1248]) );
  DFFX1_LVT u_T_427_reg_11__32_ ( .D(n4404), .CLK(n4215), .Q(n_T_427[1247]) );
  DFFX1_LVT u_T_427_reg_11__31_ ( .D(n4402), .CLK(n4215), .Q(n_T_427[1246]) );
  DFFX1_LVT u_T_427_reg_11__30_ ( .D(n4400), .CLK(n4215), .Q(n_T_427[1245]) );
  DFFX1_LVT u_T_427_reg_11__29_ ( .D(n4397), .CLK(n4215), .Q(n_T_427[1244]) );
  DFFX1_LVT u_T_427_reg_11__28_ ( .D(n4394), .CLK(n4215), .Q(n_T_427[1243]) );
  DFFX1_LVT u_T_427_reg_11__27_ ( .D(n4391), .CLK(n4215), .Q(n_T_427[1242]) );
  DFFX1_LVT u_T_427_reg_11__26_ ( .D(n4389), .CLK(n4215), .Q(n_T_427[1241]) );
  DFFX1_LVT u_T_427_reg_11__25_ ( .D(n4387), .CLK(n4215), .Q(n_T_427[1240]) );
  DFFX1_LVT u_T_427_reg_11__24_ ( .D(n4385), .CLK(n4215), .Q(n_T_427[1239]) );
  DFFX1_LVT u_T_427_reg_11__23_ ( .D(n4381), .CLK(n4214), .Q(n_T_427[1238]) );
  DFFX1_LVT u_T_427_reg_11__22_ ( .D(n4379), .CLK(n4214), .Q(n_T_427[1237]) );
  DFFX1_LVT u_T_427_reg_11__21_ ( .D(n4377), .CLK(n4214), .Q(n_T_427[1236]) );
  DFFX1_LVT u_T_427_reg_11__20_ ( .D(n4375), .CLK(n4214), .Q(n_T_427[1235]) );
  DFFX1_LVT u_T_427_reg_11__19_ ( .D(n4372), .CLK(n4214), .Q(n_T_427[1234]) );
  DFFX1_LVT u_T_427_reg_11__18_ ( .D(n4369), .CLK(n4214), .Q(n_T_427[1233]) );
  DFFX1_LVT u_T_427_reg_11__17_ ( .D(n4365), .CLK(n4214), .Q(n_T_427[1232]) );
  DFFX1_LVT u_T_427_reg_11__16_ ( .D(n4362), .CLK(n4214), .Q(n_T_427[1231]) );
  DFFX1_LVT u_T_427_reg_11__15_ ( .D(n4360), .CLK(n4214), .Q(n_T_427[1230]) );
  DFFX1_LVT u_T_427_reg_11__14_ ( .D(n4357), .CLK(n4214), .Q(n_T_427[1229]) );
  DFFX1_LVT u_T_427_reg_11__13_ ( .D(n4355), .CLK(n4214), .Q(n_T_427[1228]) );
  DFFX1_LVT u_T_427_reg_11__12_ ( .D(n4352), .CLK(n4214), .Q(n_T_427[1227]) );
  DFFX1_LVT u_T_427_reg_11__11_ ( .D(n4350), .CLK(n4213), .Q(n_T_427[1226]) );
  DFFX1_LVT u_T_427_reg_11__10_ ( .D(n4346), .CLK(n4213), .Q(n_T_427[1225]) );
  DFFX1_LVT u_T_427_reg_11__9_ ( .D(n4343), .CLK(n4213), .Q(n_T_427[1224]) );
  DFFX1_LVT u_T_427_reg_11__8_ ( .D(n4340), .CLK(n4213), .Q(n_T_427[1223]) );
  DFFX1_LVT u_T_427_reg_11__7_ ( .D(n4337), .CLK(n4213), .Q(n_T_427[1222]) );
  DFFX1_LVT u_T_427_reg_11__6_ ( .D(n4334), .CLK(n4213), .Q(n_T_427[1221]) );
  DFFX1_LVT u_T_427_reg_11__5_ ( .D(n4331), .CLK(n4213), .Q(n_T_427[1220]) );
  DFFX1_LVT u_T_427_reg_11__4_ ( .D(n4328), .CLK(n4213), .Q(n_T_427[1219]) );
  DFFX1_LVT u_T_427_reg_11__3_ ( .D(n4325), .CLK(n4213), .Q(n_T_427[1218]) );
  DFFX1_LVT u_T_427_reg_11__2_ ( .D(n4322), .CLK(n4213), .Q(n_T_427[1217]) );
  DFFX1_LVT u_T_427_reg_11__1_ ( .D(n4320), .CLK(n4213), .Q(n_T_427[1216]) );
  DFFX1_LVT u_T_427_reg_11__0_ ( .D(n4317), .CLK(n4213), .Q(n_T_427[1215]) );
  DFFX1_LVT u_T_427_reg_12__63_ ( .D(n4495), .CLK(n4212), .Q(n_T_427[1214]), 
        .QN(n3308) );
  DFFX1_LVT u_T_427_reg_12__62_ ( .D(n4492), .CLK(n4212), .Q(n_T_427[1213]), 
        .QN(n3306) );
  DFFX1_LVT u_T_427_reg_12__61_ ( .D(n4489), .CLK(n4212), .Q(n_T_427[1212]), 
        .QN(n3305) );
  DFFX1_LVT u_T_427_reg_12__60_ ( .D(n4486), .CLK(n4212), .Q(n_T_427[1211]), 
        .QN(n3304) );
  DFFX1_LVT u_T_427_reg_12__58_ ( .D(n4480), .CLK(n4211), .Q(n_T_427[1209]), 
        .QN(n3365) );
  DFFX1_LVT u_T_427_reg_12__56_ ( .D(n4474), .CLK(n4211), .Q(n_T_427[1207]), 
        .QN(n3362) );
  DFFX1_LVT u_T_427_reg_12__54_ ( .D(n4468), .CLK(n4211), .Q(n_T_427[1205]), 
        .QN(n3360) );
  DFFX1_LVT u_T_427_reg_12__52_ ( .D(n4462), .CLK(n4211), .Q(n_T_427[1203]), 
        .QN(n3355) );
  DFFX1_LVT u_T_427_reg_12__51_ ( .D(n4459), .CLK(n4211), .Q(n_T_427[1202]), 
        .QN(n3354) );
  DFFX1_LVT u_T_427_reg_12__49_ ( .D(n4453), .CLK(n4211), .Q(n_T_427[1200]), 
        .QN(n3349) );
  DFFX1_LVT u_T_427_reg_12__45_ ( .D(n4441), .CLK(n4210), .Q(n_T_427[1196]), 
        .QN(n3343) );
  DFFX1_LVT u_T_427_reg_12__43_ ( .D(n4435), .CLK(n4210), .Q(n_T_427[1194]), 
        .QN(n3340) );
  DFFX1_LVT u_T_427_reg_12__42_ ( .D(n4432), .CLK(n4210), .Q(n_T_427[1193]) );
  DFFX1_LVT u_T_427_reg_12__41_ ( .D(n4429), .CLK(n4210), .Q(n_T_427[1192]), 
        .QN(n3339) );
  DFFX1_LVT u_T_427_reg_12__39_ ( .D(n4423), .CLK(n4210), .Q(n_T_427[1190]) );
  DFFX1_LVT u_T_427_reg_12__38_ ( .D(n4420), .CLK(n4210), .Q(n_T_427[1189]) );
  DFFX1_LVT u_T_427_reg_12__36_ ( .D(n4415), .CLK(n4210), .Q(n_T_427[1187]) );
  DFFX1_LVT u_T_427_reg_12__30_ ( .D(n4400), .CLK(n4209), .Q(n_T_427[1181]), 
        .QN(n3331) );
  DFFX1_LVT u_T_427_reg_12__29_ ( .D(n4397), .CLK(n4209), .Q(n_T_427[1180]), 
        .QN(n3294) );
  DFFX1_LVT u_T_427_reg_12__27_ ( .D(n4392), .CLK(n4209), .Q(n_T_427[1178]), 
        .QN(n3328) );
  DFFX1_LVT u_T_427_reg_12__24_ ( .D(n4385), .CLK(n4209), .Q(n_T_427[1175]), 
        .QN(n3326) );
  DFFX1_LVT u_T_427_reg_12__20_ ( .D(n4375), .CLK(n4208), .Q(n_T_427[1171]), 
        .QN(n3320) );
  DFFX1_LVT u_T_427_reg_12__19_ ( .D(n4372), .CLK(n4208), .Q(n_T_427[1170]), 
        .QN(n3317) );
  DFFX1_LVT u_T_427_reg_12__18_ ( .D(n4369), .CLK(n4208), .Q(n_T_427[1169]), 
        .QN(n3314) );
  DFFX1_LVT u_T_427_reg_12__1_ ( .D(n4320), .CLK(n4207), .Q(n_T_427[1152]) );
  DFFX1_LVT u_T_427_reg_12__0_ ( .D(n4317), .CLK(n4207), .Q(n_T_427[1151]) );
  DFFX1_LVT u_T_427_reg_13__63_ ( .D(n4495), .CLK(n4206), .Q(n_T_427[1150]) );
  DFFX1_LVT u_T_427_reg_13__62_ ( .D(n4492), .CLK(n4206), .Q(n_T_427[1149]) );
  DFFX1_LVT u_T_427_reg_13__61_ ( .D(n4489), .CLK(n4206), .Q(n_T_427[1148]) );
  DFFX1_LVT u_T_427_reg_13__60_ ( .D(n4486), .CLK(n4206), .Q(n_T_427[1147]) );
  DFFX1_LVT u_T_427_reg_13__59_ ( .D(n4483), .CLK(n4205), .Q(n_T_427[1146]) );
  DFFX1_LVT u_T_427_reg_13__58_ ( .D(n4480), .CLK(n4205), .Q(n_T_427[1145]) );
  DFFX1_LVT u_T_427_reg_13__57_ ( .D(n4477), .CLK(n4205), .Q(n_T_427[1144]) );
  DFFX1_LVT u_T_427_reg_13__56_ ( .D(n4474), .CLK(n4205), .Q(n_T_427[1143]) );
  DFFX1_LVT u_T_427_reg_13__55_ ( .D(n4471), .CLK(n4205), .Q(n_T_427[1142]) );
  DFFX1_LVT u_T_427_reg_13__54_ ( .D(n4468), .CLK(n4205), .Q(n_T_427[1141]) );
  DFFX1_LVT u_T_427_reg_13__53_ ( .D(n4465), .CLK(n4205), .Q(n_T_427[1140]) );
  DFFX1_LVT u_T_427_reg_13__52_ ( .D(n4462), .CLK(n4205), .Q(n_T_427[1139]) );
  DFFX1_LVT u_T_427_reg_13__51_ ( .D(n4459), .CLK(n4205), .Q(n_T_427[1138]) );
  DFFX1_LVT u_T_427_reg_13__50_ ( .D(n4456), .CLK(n4205), .Q(n_T_427[1137]) );
  DFFX1_LVT u_T_427_reg_13__49_ ( .D(n4453), .CLK(n4205), .Q(n_T_427[1136]) );
  DFFX1_LVT u_T_427_reg_13__48_ ( .D(n4450), .CLK(n4205), .Q(n_T_427[1135]) );
  DFFX1_LVT u_T_427_reg_13__47_ ( .D(n4447), .CLK(n4204), .Q(n_T_427[1134]) );
  DFFX1_LVT u_T_427_reg_13__46_ ( .D(n4444), .CLK(n4204), .Q(n_T_427[1133]) );
  DFFX1_LVT u_T_427_reg_13__45_ ( .D(n4441), .CLK(n4204), .Q(n_T_427[1132]) );
  DFFX1_LVT u_T_427_reg_13__44_ ( .D(n4438), .CLK(n4204), .Q(n_T_427[1131]) );
  DFFX1_LVT u_T_427_reg_13__43_ ( .D(n4435), .CLK(n4204), .Q(n_T_427[1130]) );
  DFFX1_LVT u_T_427_reg_13__42_ ( .D(n4432), .CLK(n4204), .Q(n_T_427[1129]) );
  DFFX1_LVT u_T_427_reg_13__41_ ( .D(n4429), .CLK(n4204), .Q(n_T_427[1128]) );
  DFFX1_LVT u_T_427_reg_13__40_ ( .D(n4426), .CLK(n4204), .Q(n_T_427[1127]) );
  DFFX1_LVT u_T_427_reg_13__39_ ( .D(n4423), .CLK(n4204), .Q(n_T_427[1126]) );
  DFFX1_LVT u_T_427_reg_13__38_ ( .D(n4420), .CLK(n4204), .Q(n_T_427[1125]) );
  DFFX1_LVT u_T_427_reg_13__37_ ( .D(n4418), .CLK(n4204), .Q(n_T_427[1124]) );
  DFFX1_LVT u_T_427_reg_13__36_ ( .D(n4415), .CLK(n4204), .Q(n_T_427[1123]) );
  DFFX1_LVT u_T_427_reg_13__35_ ( .D(n4412), .CLK(n4203), .Q(n_T_427[1122]) );
  DFFX1_LVT u_T_427_reg_13__34_ ( .D(n4410), .CLK(n4203), .Q(n_T_427[1121]) );
  DFFX1_LVT u_T_427_reg_13__33_ ( .D(n4407), .CLK(n4203), .Q(n_T_427[1120]) );
  DFFX1_LVT u_T_427_reg_13__32_ ( .D(n4405), .CLK(n4203), .Q(n_T_427[1119]) );
  DFFX1_LVT u_T_427_reg_13__31_ ( .D(n4402), .CLK(n4203), .Q(n_T_427[1118]) );
  DFFX1_LVT u_T_427_reg_13__30_ ( .D(n4400), .CLK(n4203), .Q(n_T_427[1117]) );
  DFFX1_LVT u_T_427_reg_13__29_ ( .D(n4397), .CLK(n4203), .Q(n_T_427[1116]) );
  DFFX1_LVT u_T_427_reg_13__28_ ( .D(n4394), .CLK(n4203), .Q(n_T_427[1115]) );
  DFFX1_LVT u_T_427_reg_13__27_ ( .D(n4392), .CLK(n4203), .Q(n_T_427[1114]) );
  DFFX1_LVT u_T_427_reg_13__26_ ( .D(n4389), .CLK(n4203), .Q(n_T_427[1113]) );
  DFFX1_LVT u_T_427_reg_13__25_ ( .D(n4387), .CLK(n4203), .Q(n_T_427[1112]) );
  DFFX1_LVT u_T_427_reg_13__24_ ( .D(n4385), .CLK(n4203), .Q(n_T_427[1111]) );
  DFFX1_LVT u_T_427_reg_13__23_ ( .D(n4382), .CLK(n4202), .Q(n_T_427[1110]) );
  DFFX1_LVT u_T_427_reg_13__22_ ( .D(n4379), .CLK(n4202), .Q(n_T_427[1109]) );
  DFFX1_LVT u_T_427_reg_13__21_ ( .D(n4377), .CLK(n4202), .Q(n_T_427[1108]) );
  DFFX1_LVT u_T_427_reg_13__20_ ( .D(n4375), .CLK(n4202), .Q(n_T_427[1107]) );
  DFFX1_LVT u_T_427_reg_13__19_ ( .D(n4372), .CLK(n4202), .Q(n_T_427[1106]) );
  DFFX1_LVT u_T_427_reg_13__18_ ( .D(n4369), .CLK(n4202), .Q(n_T_427[1105]) );
  DFFX1_LVT u_T_427_reg_13__17_ ( .D(n4366), .CLK(n4202), .Q(n_T_427[1104]) );
  DFFX1_LVT u_T_427_reg_13__16_ ( .D(n4363), .CLK(n4202), .Q(n_T_427[1103]) );
  DFFX1_LVT u_T_427_reg_13__15_ ( .D(n4360), .CLK(n4202), .Q(n_T_427[1102]) );
  DFFX1_LVT u_T_427_reg_13__14_ ( .D(n4358), .CLK(n4202), .Q(n_T_427[1101]) );
  DFFX1_LVT u_T_427_reg_13__13_ ( .D(n4355), .CLK(n4202), .Q(n_T_427[1100]) );
  DFFX1_LVT u_T_427_reg_13__12_ ( .D(n4353), .CLK(n4202), .Q(n_T_427[1099]) );
  DFFX1_LVT u_T_427_reg_13__11_ ( .D(n4350), .CLK(n4201), .Q(n_T_427[1098]) );
  DFFX1_LVT u_T_427_reg_13__10_ ( .D(n4347), .CLK(n4201), .Q(n_T_427[1097]) );
  DFFX1_LVT u_T_427_reg_13__9_ ( .D(n4344), .CLK(n4201), .Q(n_T_427[1096]) );
  DFFX1_LVT u_T_427_reg_13__8_ ( .D(n4341), .CLK(n4201), .Q(n_T_427[1095]) );
  DFFX1_LVT u_T_427_reg_13__7_ ( .D(n4338), .CLK(n4201), .Q(n_T_427[1094]) );
  DFFX1_LVT u_T_427_reg_13__6_ ( .D(n4335), .CLK(n4201), .Q(n_T_427[1093]) );
  DFFX1_LVT u_T_427_reg_13__5_ ( .D(n4332), .CLK(n4201), .Q(n_T_427[1092]) );
  DFFX1_LVT u_T_427_reg_13__4_ ( .D(n4329), .CLK(n4201), .Q(n_T_427[1091]) );
  DFFX1_LVT u_T_427_reg_13__3_ ( .D(n4326), .CLK(n4201), .Q(n_T_427[1090]) );
  DFFX1_LVT u_T_427_reg_13__2_ ( .D(n4323), .CLK(n4201), .Q(n_T_427[1089]) );
  DFFX1_LVT u_T_427_reg_13__1_ ( .D(n4320), .CLK(n4201), .Q(n_T_427[1088]) );
  DFFX1_LVT u_T_427_reg_13__0_ ( .D(n4317), .CLK(n4201), .Q(n_T_427[1087]) );
  DFFX1_LVT u_T_427_reg_14__63_ ( .D(n4495), .CLK(n4200), .Q(n_T_427[1086]), 
        .QN(n3309) );
  DFFX1_LVT u_T_427_reg_14__62_ ( .D(n4492), .CLK(n4200), .Q(n_T_427[1085]), 
        .QN(n3307) );
  DFFX1_LVT u_T_427_reg_14__61_ ( .D(n4489), .CLK(n4200), .Q(n_T_427[1084]), 
        .QN(n3281) );
  DFFX1_LVT u_T_427_reg_14__60_ ( .D(n4486), .CLK(n4200), .Q(n_T_427[1083]), 
        .QN(n3303) );
  DFFX1_LVT u_T_427_reg_14__58_ ( .D(n4480), .CLK(n4199), .Q(n_T_427[1081]), 
        .QN(n3366) );
  DFFX1_LVT u_T_427_reg_14__56_ ( .D(n4474), .CLK(n4199), .Q(n_T_427[1079]) );
  DFFX1_LVT u_T_427_reg_14__55_ ( .D(n4471), .CLK(n4199), .Q(n_T_427[1078]) );
  DFFX1_LVT u_T_427_reg_14__54_ ( .D(n4468), .CLK(n4199), .Q(n_T_427[1077]), 
        .QN(n3359) );
  DFFX1_LVT u_T_427_reg_14__52_ ( .D(n4462), .CLK(n4199), .Q(n_T_427[1075]), 
        .QN(n3356) );
  DFFX1_LVT u_T_427_reg_14__51_ ( .D(n4459), .CLK(n4199), .Q(n_T_427[1074]), 
        .QN(n3353) );
  DFFX1_LVT u_T_427_reg_14__49_ ( .D(n4453), .CLK(n4199), .Q(n_T_427[1072]), 
        .QN(n3350) );
  DFFX1_LVT u_T_427_reg_14__48_ ( .D(n4450), .CLK(n4199), .Q(n_T_427[1071]) );
  DFFX1_LVT u_T_427_reg_14__45_ ( .D(n4441), .CLK(n4198), .Q(n_T_427[1068]), 
        .QN(n3344) );
  DFFX1_LVT u_T_427_reg_14__44_ ( .D(n4438), .CLK(n4198), .Q(n_T_427[1067]) );
  DFFX1_LVT u_T_427_reg_14__43_ ( .D(n4435), .CLK(n4198), .Q(n_T_427[1066]), 
        .QN(n3341) );
  DFFX1_LVT u_T_427_reg_14__42_ ( .D(n4432), .CLK(n4198), .Q(n_T_427[1065]) );
  DFFX1_LVT u_T_427_reg_14__41_ ( .D(n4429), .CLK(n4198), .Q(n_T_427[1064]) );
  DFFX1_LVT u_T_427_reg_14__39_ ( .D(n4423), .CLK(n4198), .Q(n_T_427[1062]) );
  DFFX1_LVT u_T_427_reg_14__38_ ( .D(n4420), .CLK(n4198), .Q(n_T_427[1061]) );
  DFFX1_LVT u_T_427_reg_14__37_ ( .D(n4418), .CLK(n4198), .Q(n_T_427[1060]) );
  DFFX1_LVT u_T_427_reg_14__36_ ( .D(n4415), .CLK(n4198), .Q(n_T_427[1059]) );
  DFFX1_LVT u_T_427_reg_14__35_ ( .D(n4412), .CLK(n4197), .Q(n_T_427[1058]) );
  DFFX1_LVT u_T_427_reg_14__34_ ( .D(n4410), .CLK(n4197), .Q(n_T_427[1057]) );
  DFFX1_LVT u_T_427_reg_14__33_ ( .D(n4407), .CLK(n4197), .Q(n_T_427[1056]) );
  DFFX1_LVT u_T_427_reg_14__30_ ( .D(n4400), .CLK(n4197), .Q(n_T_427[1053]), 
        .QN(n3332) );
  DFFX1_LVT u_T_427_reg_14__29_ ( .D(n4397), .CLK(n4197), .Q(n_T_427[1052]), 
        .QN(n3295) );
  DFFX1_LVT u_T_427_reg_14__27_ ( .D(n4392), .CLK(n4197), .Q(n_T_427[1050]), 
        .QN(n3329) );
  DFFX1_LVT u_T_427_reg_14__24_ ( .D(n4385), .CLK(n4197), .Q(n_T_427[1047]), 
        .QN(n3327) );
  DFFX1_LVT u_T_427_reg_14__20_ ( .D(n4375), .CLK(n4196), .Q(n_T_427[1043]), 
        .QN(n3321) );
  DFFX1_LVT u_T_427_reg_14__19_ ( .D(n4372), .CLK(n4196), .Q(n_T_427[1042]), 
        .QN(n3318) );
  DFFX1_LVT u_T_427_reg_14__18_ ( .D(n4369), .CLK(n4196), .Q(n_T_427[1041]), 
        .QN(n3315) );
  DFFX1_LVT u_T_427_reg_14__15_ ( .D(n4360), .CLK(n4196), .Q(n_T_427[1038]) );
  DFFX1_LVT u_T_427_reg_14__14_ ( .D(n4358), .CLK(n4196), .Q(n_T_427[1037]) );
  DFFX1_LVT u_T_427_reg_14__13_ ( .D(n4355), .CLK(n4196), .Q(n_T_427[1036]) );
  DFFX1_LVT u_T_427_reg_14__12_ ( .D(n4353), .CLK(n4196), .Q(n_T_427[1035]) );
  DFFX1_LVT u_T_427_reg_14__11_ ( .D(n4350), .CLK(n4195), .Q(n_T_427[1034]) );
  DFFX1_LVT u_T_427_reg_14__10_ ( .D(n4347), .CLK(n4195), .Q(n_T_427[1033]) );
  DFFX1_LVT u_T_427_reg_14__9_ ( .D(n4344), .CLK(n4195), .Q(n_T_427[1032]) );
  DFFX1_LVT u_T_427_reg_14__8_ ( .D(n4341), .CLK(n4195), .Q(n_T_427[1031]) );
  DFFX1_LVT u_T_427_reg_14__7_ ( .D(n4338), .CLK(n4195), .Q(n_T_427[1030]) );
  DFFX1_LVT u_T_427_reg_14__6_ ( .D(n4335), .CLK(n4195), .Q(n_T_427[1029]) );
  DFFX1_LVT u_T_427_reg_14__5_ ( .D(n4332), .CLK(n4195), .Q(n_T_427[1028]) );
  DFFX1_LVT u_T_427_reg_14__4_ ( .D(n4329), .CLK(n4195), .Q(n_T_427[1027]) );
  DFFX1_LVT u_T_427_reg_14__3_ ( .D(n4326), .CLK(n4195), .Q(n_T_427[1026]) );
  DFFX1_LVT u_T_427_reg_14__2_ ( .D(n4323), .CLK(n4195), .Q(n_T_427[1025]) );
  DFFX1_LVT u_T_427_reg_14__1_ ( .D(n4320), .CLK(n4195), .Q(n_T_427[1024]) );
  DFFX1_LVT u_T_427_reg_14__0_ ( .D(n4317), .CLK(n4195), .Q(n_T_427[1023]) );
  DFFX1_LVT u_T_427_reg_15__63_ ( .D(n4495), .CLK(n4194), .Q(n_T_427[1022]) );
  DFFX1_LVT u_T_427_reg_15__62_ ( .D(n4492), .CLK(n4194), .Q(n_T_427[1021]) );
  DFFX1_LVT u_T_427_reg_15__61_ ( .D(n4489), .CLK(n4194), .Q(n_T_427[1020]) );
  DFFX1_LVT u_T_427_reg_15__60_ ( .D(n4486), .CLK(n4194), .Q(n_T_427[1019]) );
  DFFX1_LVT u_T_427_reg_15__59_ ( .D(n4483), .CLK(n4193), .Q(n_T_427[1018]) );
  DFFX1_LVT u_T_427_reg_15__58_ ( .D(n4480), .CLK(n4193), .Q(n_T_427[1017]) );
  DFFX1_LVT u_T_427_reg_15__57_ ( .D(n4477), .CLK(n4193), .Q(n_T_427[1016]) );
  DFFX1_LVT u_T_427_reg_15__56_ ( .D(n4474), .CLK(n4193), .Q(n_T_427[1015]) );
  DFFX1_LVT u_T_427_reg_15__55_ ( .D(n4471), .CLK(n4193), .Q(n_T_427[1014]) );
  DFFX1_LVT u_T_427_reg_15__54_ ( .D(n4468), .CLK(n4193), .Q(n_T_427[1013]) );
  DFFX1_LVT u_T_427_reg_15__53_ ( .D(n4465), .CLK(n4193), .Q(n_T_427[1012]) );
  DFFX1_LVT u_T_427_reg_15__52_ ( .D(n4462), .CLK(n4193), .Q(n_T_427[1011]) );
  DFFX1_LVT u_T_427_reg_15__51_ ( .D(n4459), .CLK(n4193), .Q(n_T_427[1010]) );
  DFFX1_LVT u_T_427_reg_15__50_ ( .D(n4456), .CLK(n4193), .Q(n_T_427[1009]) );
  DFFX1_LVT u_T_427_reg_15__49_ ( .D(n4453), .CLK(n4193), .Q(n_T_427[1008]) );
  DFFX1_LVT u_T_427_reg_15__48_ ( .D(n4450), .CLK(n4193), .Q(n_T_427[1007]) );
  DFFX1_LVT u_T_427_reg_15__47_ ( .D(n4447), .CLK(n4192), .Q(n_T_427[1006]) );
  DFFX1_LVT u_T_427_reg_15__46_ ( .D(n4444), .CLK(n4192), .Q(n_T_427[1005]) );
  DFFX1_LVT u_T_427_reg_15__45_ ( .D(n4441), .CLK(n4192), .Q(n_T_427[1004]) );
  DFFX1_LVT u_T_427_reg_15__44_ ( .D(n4438), .CLK(n4192), .Q(n_T_427[1003]) );
  DFFX1_LVT u_T_427_reg_15__43_ ( .D(n4435), .CLK(n4192), .Q(n_T_427[1002]) );
  DFFX1_LVT u_T_427_reg_15__42_ ( .D(n4432), .CLK(n4192), .Q(n_T_427[1001]) );
  DFFX1_LVT u_T_427_reg_15__41_ ( .D(n4429), .CLK(n4192), .Q(n_T_427[1000]) );
  DFFX1_LVT u_T_427_reg_15__40_ ( .D(n4426), .CLK(n4192), .Q(n_T_427[999]) );
  DFFX1_LVT u_T_427_reg_15__39_ ( .D(n4423), .CLK(n4192), .Q(n_T_427[998]) );
  DFFX1_LVT u_T_427_reg_15__38_ ( .D(n4420), .CLK(n4192), .Q(n_T_427[997]) );
  DFFX1_LVT u_T_427_reg_15__37_ ( .D(n4418), .CLK(n4192), .Q(n_T_427[996]) );
  DFFX1_LVT u_T_427_reg_15__36_ ( .D(n4415), .CLK(n4192), .Q(n_T_427[995]) );
  DFFX1_LVT u_T_427_reg_15__35_ ( .D(n4412), .CLK(n4191), .Q(n_T_427[994]) );
  DFFX1_LVT u_T_427_reg_15__34_ ( .D(n4410), .CLK(n4191), .Q(n_T_427[993]) );
  DFFX1_LVT u_T_427_reg_15__33_ ( .D(n4407), .CLK(n4191), .Q(n_T_427[992]) );
  DFFX1_LVT u_T_427_reg_15__32_ ( .D(n4405), .CLK(n4191), .Q(n_T_427[991]) );
  DFFX1_LVT u_T_427_reg_15__31_ ( .D(n4402), .CLK(n4191), .Q(n_T_427[990]) );
  DFFX1_LVT u_T_427_reg_15__30_ ( .D(n4400), .CLK(n4191), .Q(n_T_427[989]) );
  DFFX1_LVT u_T_427_reg_15__29_ ( .D(n4397), .CLK(n4191), .Q(n_T_427[988]) );
  DFFX1_LVT u_T_427_reg_15__28_ ( .D(n4394), .CLK(n4191), .Q(n_T_427[987]) );
  DFFX1_LVT u_T_427_reg_15__27_ ( .D(n4392), .CLK(n4191), .Q(n_T_427[986]) );
  DFFX1_LVT u_T_427_reg_15__26_ ( .D(n4389), .CLK(n4191), .Q(n_T_427[985]) );
  DFFX1_LVT u_T_427_reg_15__25_ ( .D(n4387), .CLK(n4191), .Q(n_T_427[984]) );
  DFFX1_LVT u_T_427_reg_15__24_ ( .D(n4385), .CLK(n4191), .Q(n_T_427[983]) );
  DFFX1_LVT u_T_427_reg_15__23_ ( .D(n4382), .CLK(n4190), .Q(n_T_427[982]) );
  DFFX1_LVT u_T_427_reg_15__22_ ( .D(n4379), .CLK(n4190), .Q(n_T_427[981]) );
  DFFX1_LVT u_T_427_reg_15__21_ ( .D(n4377), .CLK(n4190), .Q(n_T_427[980]) );
  DFFX1_LVT u_T_427_reg_15__20_ ( .D(n4375), .CLK(n4190), .Q(n_T_427[979]) );
  DFFX1_LVT u_T_427_reg_15__19_ ( .D(n4372), .CLK(n4190), .Q(n_T_427[978]) );
  DFFX1_LVT u_T_427_reg_15__18_ ( .D(n4369), .CLK(n4190), .Q(n_T_427[977]) );
  DFFX1_LVT u_T_427_reg_15__17_ ( .D(n4366), .CLK(n4190), .Q(n_T_427[976]) );
  DFFX1_LVT u_T_427_reg_15__16_ ( .D(n4363), .CLK(n4190), .Q(n_T_427[975]) );
  DFFX1_LVT u_T_427_reg_15__15_ ( .D(n4360), .CLK(n4190), .Q(n_T_427[974]) );
  DFFX1_LVT u_T_427_reg_15__14_ ( .D(n4358), .CLK(n4190), .Q(n_T_427[973]) );
  DFFX1_LVT u_T_427_reg_15__13_ ( .D(n4355), .CLK(n4190), .Q(n_T_427[972]) );
  DFFX1_LVT u_T_427_reg_15__12_ ( .D(n4353), .CLK(n4190), .Q(n_T_427[971]) );
  DFFX1_LVT u_T_427_reg_15__11_ ( .D(n4350), .CLK(n4189), .Q(n_T_427[970]) );
  DFFX1_LVT u_T_427_reg_15__10_ ( .D(n4347), .CLK(n4189), .Q(n_T_427[969]) );
  DFFX1_LVT u_T_427_reg_15__9_ ( .D(n4344), .CLK(n4189), .Q(n_T_427[968]) );
  DFFX1_LVT u_T_427_reg_15__8_ ( .D(n4341), .CLK(n4189), .Q(n_T_427[967]) );
  DFFX1_LVT u_T_427_reg_15__7_ ( .D(n4338), .CLK(n4189), .Q(n_T_427[966]) );
  DFFX1_LVT u_T_427_reg_15__6_ ( .D(n4335), .CLK(n4189), .Q(n_T_427[965]) );
  DFFX1_LVT u_T_427_reg_15__5_ ( .D(n4332), .CLK(n4189), .Q(n_T_427[964]) );
  DFFX1_LVT u_T_427_reg_15__4_ ( .D(n4329), .CLK(n4189), .Q(n_T_427[963]) );
  DFFX1_LVT u_T_427_reg_15__3_ ( .D(n4326), .CLK(n4189), .Q(n_T_427[962]) );
  DFFX1_LVT u_T_427_reg_15__2_ ( .D(n4323), .CLK(n4189), .Q(n_T_427[961]) );
  DFFX1_LVT u_T_427_reg_15__1_ ( .D(n4320), .CLK(n4189), .Q(n_T_427[960]) );
  DFFX1_LVT u_T_427_reg_15__0_ ( .D(n4317), .CLK(n4189), .Q(n_T_427[959]) );
  DFFX1_LVT u_T_427_reg_16__63_ ( .D(n4495), .CLK(n4188), .Q(n_T_427[958]) );
  DFFX1_LVT u_T_427_reg_16__62_ ( .D(n4492), .CLK(n4188), .Q(n_T_427[957]) );
  DFFX1_LVT u_T_427_reg_16__61_ ( .D(n4489), .CLK(n4188), .Q(n_T_427[956]) );
  DFFX1_LVT u_T_427_reg_16__60_ ( .D(n4486), .CLK(n4188), .Q(n_T_427[955]) );
  DFFX1_LVT u_T_427_reg_16__59_ ( .D(n4483), .CLK(n4187), .Q(n_T_427[954]) );
  DFFX1_LVT u_T_427_reg_16__58_ ( .D(n4480), .CLK(n4187), .Q(n_T_427[953]) );
  DFFX1_LVT u_T_427_reg_16__57_ ( .D(n4477), .CLK(n4187), .Q(n_T_427[952]) );
  DFFX1_LVT u_T_427_reg_16__56_ ( .D(n4474), .CLK(n4187), .Q(n_T_427[951]) );
  DFFX1_LVT u_T_427_reg_16__55_ ( .D(n4471), .CLK(n4187), .Q(n_T_427[950]) );
  DFFX1_LVT u_T_427_reg_16__54_ ( .D(n4468), .CLK(n4187), .Q(n_T_427[949]) );
  DFFX1_LVT u_T_427_reg_16__53_ ( .D(n4465), .CLK(n4187), .Q(n_T_427[948]) );
  DFFX1_LVT u_T_427_reg_16__52_ ( .D(n4462), .CLK(n4187), .Q(n_T_427[947]) );
  DFFX1_LVT u_T_427_reg_16__51_ ( .D(n4459), .CLK(n4187), .Q(n_T_427[946]) );
  DFFX1_LVT u_T_427_reg_16__50_ ( .D(n4456), .CLK(n4187), .Q(n_T_427[945]) );
  DFFX1_LVT u_T_427_reg_16__49_ ( .D(n4453), .CLK(n4187), .Q(n_T_427[944]) );
  DFFX1_LVT u_T_427_reg_16__48_ ( .D(n4450), .CLK(n4187), .Q(n_T_427[943]) );
  DFFX1_LVT u_T_427_reg_16__47_ ( .D(n4447), .CLK(n4186), .Q(n_T_427[942]) );
  DFFX1_LVT u_T_427_reg_16__46_ ( .D(n4444), .CLK(n4186), .Q(n_T_427[941]) );
  DFFX1_LVT u_T_427_reg_16__45_ ( .D(n4441), .CLK(n4186), .Q(n_T_427[940]) );
  DFFX1_LVT u_T_427_reg_16__44_ ( .D(n4438), .CLK(n4186), .Q(n_T_427[939]) );
  DFFX1_LVT u_T_427_reg_16__43_ ( .D(n4435), .CLK(n4186), .Q(n_T_427[938]) );
  DFFX1_LVT u_T_427_reg_16__42_ ( .D(n4432), .CLK(n4186), .Q(n_T_427[937]) );
  DFFX1_LVT u_T_427_reg_16__41_ ( .D(n4429), .CLK(n4186), .Q(n_T_427[936]) );
  DFFX1_LVT u_T_427_reg_16__40_ ( .D(n4426), .CLK(n4186), .Q(n_T_427[935]) );
  DFFX1_LVT u_T_427_reg_16__39_ ( .D(n4423), .CLK(n4186), .Q(n_T_427[934]) );
  DFFX1_LVT u_T_427_reg_16__38_ ( .D(n4420), .CLK(n4186), .Q(n_T_427[933]) );
  DFFX1_LVT u_T_427_reg_16__37_ ( .D(n4418), .CLK(n4186), .Q(n_T_427[932]) );
  DFFX1_LVT u_T_427_reg_16__36_ ( .D(n4415), .CLK(n4186), .Q(n_T_427[931]) );
  DFFX1_LVT u_T_427_reg_16__35_ ( .D(n4412), .CLK(n4185), .Q(n_T_427[930]) );
  DFFX1_LVT u_T_427_reg_16__34_ ( .D(n4410), .CLK(n4185), .Q(n_T_427[929]) );
  DFFX1_LVT u_T_427_reg_16__33_ ( .D(n4407), .CLK(n4185), .Q(n_T_427[928]) );
  DFFX1_LVT u_T_427_reg_16__32_ ( .D(n4405), .CLK(n4185), .Q(n_T_427[927]) );
  DFFX1_LVT u_T_427_reg_16__31_ ( .D(n4402), .CLK(n4185), .Q(n_T_427[926]) );
  DFFX1_LVT u_T_427_reg_16__30_ ( .D(n4400), .CLK(n4185), .Q(n_T_427[925]) );
  DFFX1_LVT u_T_427_reg_16__29_ ( .D(n4397), .CLK(n4185), .Q(n_T_427[924]) );
  DFFX1_LVT u_T_427_reg_16__28_ ( .D(n4394), .CLK(n4185), .Q(n_T_427[923]) );
  DFFX1_LVT u_T_427_reg_16__27_ ( .D(n4392), .CLK(n4185), .Q(n_T_427[922]) );
  DFFX1_LVT u_T_427_reg_16__26_ ( .D(n4389), .CLK(n4185), .Q(n_T_427[921]) );
  DFFX1_LVT u_T_427_reg_16__25_ ( .D(n4387), .CLK(n4185), .Q(n_T_427[920]) );
  DFFX1_LVT u_T_427_reg_16__24_ ( .D(n4385), .CLK(n4185), .Q(n_T_427[919]) );
  DFFX1_LVT u_T_427_reg_16__23_ ( .D(n4382), .CLK(n4184), .Q(n_T_427[918]) );
  DFFX1_LVT u_T_427_reg_16__22_ ( .D(n4379), .CLK(n4184), .Q(n_T_427[917]) );
  DFFX1_LVT u_T_427_reg_16__21_ ( .D(n4377), .CLK(n4184), .Q(n_T_427[916]) );
  DFFX1_LVT u_T_427_reg_16__20_ ( .D(n4375), .CLK(n4184), .Q(n_T_427[915]) );
  DFFX1_LVT u_T_427_reg_16__19_ ( .D(n4372), .CLK(n4184), .Q(n_T_427[914]) );
  DFFX1_LVT u_T_427_reg_16__18_ ( .D(n4369), .CLK(n4184), .Q(n_T_427[913]) );
  DFFX1_LVT u_T_427_reg_16__17_ ( .D(n4366), .CLK(n4184), .Q(n_T_427[912]) );
  DFFX1_LVT u_T_427_reg_16__16_ ( .D(n4363), .CLK(n4184), .Q(n_T_427[911]) );
  DFFX1_LVT u_T_427_reg_16__15_ ( .D(n4360), .CLK(n4184), .Q(n_T_427[910]) );
  DFFX1_LVT u_T_427_reg_16__14_ ( .D(n4358), .CLK(n4184), .Q(n_T_427[909]) );
  DFFX1_LVT u_T_427_reg_16__13_ ( .D(n4355), .CLK(n4184), .Q(n_T_427[908]) );
  DFFX1_LVT u_T_427_reg_16__12_ ( .D(n4353), .CLK(n4184), .Q(n_T_427[907]) );
  DFFX1_LVT u_T_427_reg_16__11_ ( .D(n4350), .CLK(n4183), .Q(n_T_427[906]) );
  DFFX1_LVT u_T_427_reg_16__10_ ( .D(n4347), .CLK(n4183), .Q(n_T_427[905]) );
  DFFX1_LVT u_T_427_reg_16__9_ ( .D(n4344), .CLK(n4183), .Q(n_T_427[904]) );
  DFFX1_LVT u_T_427_reg_16__8_ ( .D(n4341), .CLK(n4183), .Q(n_T_427[903]) );
  DFFX1_LVT u_T_427_reg_16__7_ ( .D(n4338), .CLK(n4183), .Q(n_T_427[902]) );
  DFFX1_LVT u_T_427_reg_16__6_ ( .D(n4335), .CLK(n4183), .Q(n_T_427[901]) );
  DFFX1_LVT u_T_427_reg_16__5_ ( .D(n4332), .CLK(n4183), .Q(n_T_427[900]) );
  DFFX1_LVT u_T_427_reg_16__4_ ( .D(n4329), .CLK(n4183), .Q(n_T_427[899]) );
  DFFX1_LVT u_T_427_reg_16__3_ ( .D(n4326), .CLK(n4183), .Q(n_T_427[898]) );
  DFFX1_LVT u_T_427_reg_16__2_ ( .D(n4323), .CLK(n4183), .Q(n_T_427[897]) );
  DFFX1_LVT u_T_427_reg_16__1_ ( .D(n4320), .CLK(n4183), .Q(n_T_427[896]) );
  DFFX1_LVT u_T_427_reg_16__0_ ( .D(n4317), .CLK(n4183), .Q(n_T_427[895]) );
  DFFX1_LVT u_T_427_reg_17__63_ ( .D(n4495), .CLK(n4182), .Q(n_T_427[894]) );
  DFFX1_LVT u_T_427_reg_17__62_ ( .D(n4492), .CLK(n4182), .Q(n_T_427[893]) );
  DFFX1_LVT u_T_427_reg_17__61_ ( .D(n4489), .CLK(n4182), .Q(n_T_427[892]) );
  DFFX1_LVT u_T_427_reg_17__60_ ( .D(n4486), .CLK(n4182), .Q(n_T_427[891]) );
  DFFX1_LVT u_T_427_reg_17__59_ ( .D(n4483), .CLK(n4181), .Q(n_T_427[890]) );
  DFFX1_LVT u_T_427_reg_17__58_ ( .D(n4480), .CLK(n4181), .Q(n_T_427[889]) );
  DFFX1_LVT u_T_427_reg_17__57_ ( .D(n4477), .CLK(n4181), .Q(n_T_427[888]) );
  DFFX1_LVT u_T_427_reg_17__56_ ( .D(n4474), .CLK(n4181), .Q(n_T_427[887]) );
  DFFX1_LVT u_T_427_reg_17__55_ ( .D(n4471), .CLK(n4181), .Q(n_T_427[886]) );
  DFFX1_LVT u_T_427_reg_17__54_ ( .D(n4468), .CLK(n4181), .Q(n_T_427[885]) );
  DFFX1_LVT u_T_427_reg_17__53_ ( .D(n4465), .CLK(n4181), .Q(n_T_427[884]) );
  DFFX1_LVT u_T_427_reg_17__52_ ( .D(n4462), .CLK(n4181), .Q(n_T_427[883]) );
  DFFX1_LVT u_T_427_reg_17__51_ ( .D(n4459), .CLK(n4181), .Q(n_T_427[882]) );
  DFFX1_LVT u_T_427_reg_17__50_ ( .D(n4456), .CLK(n4181), .Q(n_T_427[881]) );
  DFFX1_LVT u_T_427_reg_17__49_ ( .D(n4453), .CLK(n4181), .Q(n_T_427[880]) );
  DFFX1_LVT u_T_427_reg_17__48_ ( .D(n4450), .CLK(n4181), .Q(n_T_427[879]) );
  DFFX1_LVT u_T_427_reg_17__47_ ( .D(n4447), .CLK(n4180), .Q(n_T_427[878]) );
  DFFX1_LVT u_T_427_reg_17__46_ ( .D(n4444), .CLK(n4180), .Q(n_T_427[877]) );
  DFFX1_LVT u_T_427_reg_17__45_ ( .D(n4441), .CLK(n4180), .Q(n_T_427[876]) );
  DFFX1_LVT u_T_427_reg_17__44_ ( .D(n4438), .CLK(n4180), .Q(n_T_427[875]) );
  DFFX1_LVT u_T_427_reg_17__43_ ( .D(n4435), .CLK(n4180), .Q(n_T_427[874]) );
  DFFX1_LVT u_T_427_reg_17__42_ ( .D(n4432), .CLK(n4180), .Q(n_T_427[873]) );
  DFFX1_LVT u_T_427_reg_17__41_ ( .D(n4429), .CLK(n4180), .Q(n_T_427[872]) );
  DFFX1_LVT u_T_427_reg_17__40_ ( .D(n4426), .CLK(n4180), .Q(n_T_427[871]) );
  DFFX1_LVT u_T_427_reg_17__39_ ( .D(n4423), .CLK(n4180), .Q(n_T_427[870]) );
  DFFX1_LVT u_T_427_reg_17__38_ ( .D(n4420), .CLK(n4180), .Q(n_T_427[869]) );
  DFFX1_LVT u_T_427_reg_17__37_ ( .D(n4418), .CLK(n4180), .Q(n_T_427[868]) );
  DFFX1_LVT u_T_427_reg_17__36_ ( .D(n4415), .CLK(n4180), .Q(n_T_427[867]) );
  DFFX1_LVT u_T_427_reg_17__35_ ( .D(n4412), .CLK(n4179), .Q(n_T_427[866]) );
  DFFX1_LVT u_T_427_reg_17__34_ ( .D(n4410), .CLK(n4179), .Q(n_T_427[865]) );
  DFFX1_LVT u_T_427_reg_17__33_ ( .D(n4407), .CLK(n4179), .Q(n_T_427[864]) );
  DFFX1_LVT u_T_427_reg_17__32_ ( .D(n4405), .CLK(n4179), .Q(n_T_427[863]) );
  DFFX1_LVT u_T_427_reg_17__31_ ( .D(n4402), .CLK(n4179), .Q(n_T_427[862]) );
  DFFX1_LVT u_T_427_reg_17__30_ ( .D(n4400), .CLK(n4179), .Q(n_T_427[861]) );
  DFFX1_LVT u_T_427_reg_17__29_ ( .D(n4397), .CLK(n4179), .Q(n_T_427[860]) );
  DFFX1_LVT u_T_427_reg_17__28_ ( .D(n4394), .CLK(n4179), .Q(n_T_427[859]) );
  DFFX1_LVT u_T_427_reg_17__27_ ( .D(n4392), .CLK(n4179), .Q(n_T_427[858]) );
  DFFX1_LVT u_T_427_reg_17__26_ ( .D(n4389), .CLK(n4179), .Q(n_T_427[857]) );
  DFFX1_LVT u_T_427_reg_17__25_ ( .D(n4387), .CLK(n4179), .Q(n_T_427[856]) );
  DFFX1_LVT u_T_427_reg_17__24_ ( .D(n4385), .CLK(n4179), .Q(n_T_427[855]) );
  DFFX1_LVT u_T_427_reg_17__23_ ( .D(n4382), .CLK(n4178), .Q(n_T_427[854]) );
  DFFX1_LVT u_T_427_reg_17__22_ ( .D(n4379), .CLK(n4178), .Q(n_T_427[853]) );
  DFFX1_LVT u_T_427_reg_17__21_ ( .D(n4377), .CLK(n4178), .Q(n_T_427[852]) );
  DFFX1_LVT u_T_427_reg_17__20_ ( .D(n4375), .CLK(n4178), .Q(n_T_427[851]) );
  DFFX1_LVT u_T_427_reg_17__19_ ( .D(n4372), .CLK(n4178), .Q(n_T_427[850]) );
  DFFX1_LVT u_T_427_reg_17__18_ ( .D(n4369), .CLK(n4178), .Q(n_T_427[849]) );
  DFFX1_LVT u_T_427_reg_17__17_ ( .D(n4366), .CLK(n4178), .Q(n_T_427[848]) );
  DFFX1_LVT u_T_427_reg_17__16_ ( .D(n4363), .CLK(n4178), .Q(n_T_427[847]) );
  DFFX1_LVT u_T_427_reg_17__15_ ( .D(n4360), .CLK(n4178), .Q(n_T_427[846]) );
  DFFX1_LVT u_T_427_reg_17__14_ ( .D(n4358), .CLK(n4178), .Q(n_T_427[845]) );
  DFFX1_LVT u_T_427_reg_17__13_ ( .D(n4355), .CLK(n4178), .Q(n_T_427[844]) );
  DFFX1_LVT u_T_427_reg_17__12_ ( .D(n4353), .CLK(n4178), .Q(n_T_427[843]) );
  DFFX1_LVT u_T_427_reg_17__11_ ( .D(n4350), .CLK(n4177), .Q(n_T_427[842]) );
  DFFX1_LVT u_T_427_reg_17__10_ ( .D(n4347), .CLK(n4177), .Q(n_T_427[841]) );
  DFFX1_LVT u_T_427_reg_17__9_ ( .D(n4344), .CLK(n4177), .Q(n_T_427[840]) );
  DFFX1_LVT u_T_427_reg_17__8_ ( .D(n4341), .CLK(n4177), .Q(n_T_427[839]) );
  DFFX1_LVT u_T_427_reg_17__7_ ( .D(n4338), .CLK(n4177), .Q(n_T_427[838]) );
  DFFX1_LVT u_T_427_reg_17__6_ ( .D(n4335), .CLK(n4177), .Q(n_T_427[837]) );
  DFFX1_LVT u_T_427_reg_17__5_ ( .D(n4332), .CLK(n4177), .Q(n_T_427[836]) );
  DFFX1_LVT u_T_427_reg_17__4_ ( .D(n4329), .CLK(n4177), .Q(n_T_427[835]) );
  DFFX1_LVT u_T_427_reg_17__3_ ( .D(n4326), .CLK(n4177), .Q(n_T_427[834]) );
  DFFX1_LVT u_T_427_reg_17__2_ ( .D(n4323), .CLK(n4177), .Q(n_T_427[833]) );
  DFFX1_LVT u_T_427_reg_17__1_ ( .D(n4320), .CLK(n4177), .Q(n_T_427[832]) );
  DFFX1_LVT u_T_427_reg_17__0_ ( .D(n4317), .CLK(n4177), .Q(n_T_427[831]) );
  DFFX1_LVT u_T_427_reg_18__63_ ( .D(n4495), .CLK(n4176), .Q(n_T_427[830]) );
  DFFX1_LVT u_T_427_reg_18__62_ ( .D(n4492), .CLK(n4176), .Q(n_T_427[829]) );
  DFFX1_LVT u_T_427_reg_18__61_ ( .D(n4489), .CLK(n4176), .Q(n_T_427[828]) );
  DFFX1_LVT u_T_427_reg_18__60_ ( .D(n4486), .CLK(n4176), .Q(n_T_427[827]) );
  DFFX1_LVT u_T_427_reg_18__59_ ( .D(n4483), .CLK(n4175), .Q(n_T_427[826]) );
  DFFX1_LVT u_T_427_reg_18__58_ ( .D(n4480), .CLK(n4175), .Q(n_T_427[825]) );
  DFFX1_LVT u_T_427_reg_18__57_ ( .D(n4477), .CLK(n4175), .Q(n_T_427[824]) );
  DFFX1_LVT u_T_427_reg_18__56_ ( .D(n4474), .CLK(n4175), .Q(n_T_427[823]) );
  DFFX1_LVT u_T_427_reg_18__55_ ( .D(n4471), .CLK(n4175), .Q(n_T_427[822]) );
  DFFX1_LVT u_T_427_reg_18__54_ ( .D(n4468), .CLK(n4175), .Q(n_T_427[821]) );
  DFFX1_LVT u_T_427_reg_18__53_ ( .D(n4465), .CLK(n4175), .Q(n_T_427[820]) );
  DFFX1_LVT u_T_427_reg_18__52_ ( .D(n4462), .CLK(n4175), .Q(n_T_427[819]) );
  DFFX1_LVT u_T_427_reg_18__51_ ( .D(n4459), .CLK(n4175), .Q(n_T_427[818]) );
  DFFX1_LVT u_T_427_reg_18__50_ ( .D(n4456), .CLK(n4175), .Q(n_T_427[817]) );
  DFFX1_LVT u_T_427_reg_18__49_ ( .D(n4453), .CLK(n4175), .Q(n_T_427[816]) );
  DFFX1_LVT u_T_427_reg_18__48_ ( .D(n4450), .CLK(n4175), .Q(n_T_427[815]) );
  DFFX1_LVT u_T_427_reg_18__47_ ( .D(n4447), .CLK(n4174), .Q(n_T_427[814]) );
  DFFX1_LVT u_T_427_reg_18__46_ ( .D(n4444), .CLK(n4174), .Q(n_T_427[813]) );
  DFFX1_LVT u_T_427_reg_18__45_ ( .D(n4441), .CLK(n4174), .Q(n_T_427[812]) );
  DFFX1_LVT u_T_427_reg_18__44_ ( .D(n4438), .CLK(n4174), .Q(n_T_427[811]) );
  DFFX1_LVT u_T_427_reg_18__43_ ( .D(n4435), .CLK(n4174), .Q(n_T_427[810]) );
  DFFX1_LVT u_T_427_reg_18__42_ ( .D(n4432), .CLK(n4174), .Q(n_T_427[809]) );
  DFFX1_LVT u_T_427_reg_18__41_ ( .D(n4429), .CLK(n4174), .Q(n_T_427[808]) );
  DFFX1_LVT u_T_427_reg_18__40_ ( .D(n4426), .CLK(n4174), .Q(n_T_427[807]) );
  DFFX1_LVT u_T_427_reg_18__39_ ( .D(n4423), .CLK(n4174), .Q(n_T_427[806]) );
  DFFX1_LVT u_T_427_reg_18__38_ ( .D(n4420), .CLK(n4174), .Q(n_T_427[805]) );
  DFFX1_LVT u_T_427_reg_18__37_ ( .D(n4418), .CLK(n4174), .Q(n_T_427[804]) );
  DFFX1_LVT u_T_427_reg_18__36_ ( .D(n4415), .CLK(n4174), .Q(n_T_427[803]) );
  DFFX1_LVT u_T_427_reg_18__35_ ( .D(n4412), .CLK(n4173), .Q(n_T_427[802]) );
  DFFX1_LVT u_T_427_reg_18__34_ ( .D(n4410), .CLK(n4173), .Q(n_T_427[801]) );
  DFFX1_LVT u_T_427_reg_18__33_ ( .D(n4407), .CLK(n4173), .Q(n_T_427[800]) );
  DFFX1_LVT u_T_427_reg_18__32_ ( .D(n4405), .CLK(n4173), .Q(n_T_427[799]) );
  DFFX1_LVT u_T_427_reg_18__31_ ( .D(n4402), .CLK(n4173), .Q(n_T_427[798]) );
  DFFX1_LVT u_T_427_reg_18__30_ ( .D(n4400), .CLK(n4173), .Q(n_T_427[797]) );
  DFFX1_LVT u_T_427_reg_18__29_ ( .D(n4397), .CLK(n4173), .Q(n_T_427[796]) );
  DFFX1_LVT u_T_427_reg_18__28_ ( .D(n4394), .CLK(n4173), .Q(n_T_427[795]) );
  DFFX1_LVT u_T_427_reg_18__27_ ( .D(n4392), .CLK(n4173), .Q(n_T_427[794]) );
  DFFX1_LVT u_T_427_reg_18__26_ ( .D(n4389), .CLK(n4173), .Q(n_T_427[793]) );
  DFFX1_LVT u_T_427_reg_18__25_ ( .D(n4387), .CLK(n4173), .Q(n_T_427[792]) );
  DFFX1_LVT u_T_427_reg_18__24_ ( .D(n4385), .CLK(n4173), .Q(n_T_427[791]) );
  DFFX1_LVT u_T_427_reg_18__23_ ( .D(n4382), .CLK(n4172), .Q(n_T_427[790]) );
  DFFX1_LVT u_T_427_reg_18__22_ ( .D(n4379), .CLK(n4172), .Q(n_T_427[789]) );
  DFFX1_LVT u_T_427_reg_18__21_ ( .D(n4377), .CLK(n4172), .Q(n_T_427[788]) );
  DFFX1_LVT u_T_427_reg_18__20_ ( .D(n4375), .CLK(n4172), .Q(n_T_427[787]) );
  DFFX1_LVT u_T_427_reg_18__19_ ( .D(n4372), .CLK(n4172), .Q(n_T_427[786]) );
  DFFX1_LVT u_T_427_reg_18__18_ ( .D(n4369), .CLK(n4172), .Q(n_T_427[785]) );
  DFFX1_LVT u_T_427_reg_18__17_ ( .D(n4366), .CLK(n4172), .Q(n_T_427[784]) );
  DFFX1_LVT u_T_427_reg_18__16_ ( .D(n4363), .CLK(n4172), .Q(n_T_427[783]) );
  DFFX1_LVT u_T_427_reg_18__15_ ( .D(n4360), .CLK(n4172), .Q(n_T_427[782]) );
  DFFX1_LVT u_T_427_reg_18__14_ ( .D(n4358), .CLK(n4172), .Q(n_T_427[781]) );
  DFFX1_LVT u_T_427_reg_18__13_ ( .D(n4355), .CLK(n4172), .Q(n_T_427[780]) );
  DFFX1_LVT u_T_427_reg_18__12_ ( .D(n4353), .CLK(n4172), .Q(n_T_427[779]) );
  DFFX1_LVT u_T_427_reg_18__11_ ( .D(n4350), .CLK(n4171), .Q(n_T_427[778]) );
  DFFX1_LVT u_T_427_reg_18__10_ ( .D(n4347), .CLK(n4171), .Q(n_T_427[777]) );
  DFFX1_LVT u_T_427_reg_18__9_ ( .D(n4344), .CLK(n4171), .Q(n_T_427[776]) );
  DFFX1_LVT u_T_427_reg_18__8_ ( .D(n4341), .CLK(n4171), .Q(n_T_427[775]) );
  DFFX1_LVT u_T_427_reg_18__7_ ( .D(n4338), .CLK(n4171), .Q(n_T_427[774]) );
  DFFX1_LVT u_T_427_reg_18__6_ ( .D(n4335), .CLK(n4171), .Q(n_T_427[773]) );
  DFFX1_LVT u_T_427_reg_18__5_ ( .D(n4332), .CLK(n4171), .Q(n_T_427[772]) );
  DFFX1_LVT u_T_427_reg_18__4_ ( .D(n4329), .CLK(n4171), .Q(n_T_427[771]) );
  DFFX1_LVT u_T_427_reg_18__3_ ( .D(n4326), .CLK(n4171), .Q(n_T_427[770]) );
  DFFX1_LVT u_T_427_reg_18__2_ ( .D(n4323), .CLK(n4171), .Q(n_T_427[769]) );
  DFFX1_LVT u_T_427_reg_18__1_ ( .D(n4320), .CLK(n4171), .Q(n_T_427[768]) );
  DFFX1_LVT u_T_427_reg_18__0_ ( .D(n4317), .CLK(n4171), .Q(n_T_427[767]) );
  DFFX1_LVT u_T_427_reg_19__63_ ( .D(n4495), .CLK(n4170), .Q(n_T_427[766]) );
  DFFX1_LVT u_T_427_reg_19__62_ ( .D(n4492), .CLK(n4170), .Q(n_T_427[765]) );
  DFFX1_LVT u_T_427_reg_19__61_ ( .D(n4489), .CLK(n4170), .Q(n_T_427[764]), 
        .QN(n3280) );
  DFFX1_LVT u_T_427_reg_19__60_ ( .D(n4486), .CLK(n4170), .Q(n_T_427[763]) );
  DFFX1_LVT u_T_427_reg_19__59_ ( .D(n4483), .CLK(n4169), .Q(n_T_427[762]) );
  DFFX1_LVT u_T_427_reg_19__58_ ( .D(n4479), .CLK(n4169), .Q(n_T_427[761]) );
  DFFX1_LVT u_T_427_reg_19__56_ ( .D(n4473), .CLK(n4169), .Q(n_T_427[759]) );
  DFFX1_LVT u_T_427_reg_19__54_ ( .D(n4467), .CLK(n4169), .Q(n_T_427[757]) );
  DFFX1_LVT u_T_427_reg_19__53_ ( .D(n4465), .CLK(n4169), .Q(n_T_427[756]) );
  DFFX1_LVT u_T_427_reg_19__52_ ( .D(n4461), .CLK(n4169), .Q(n_T_427[755]), 
        .QN(n3408) );
  DFFX1_LVT u_T_427_reg_19__51_ ( .D(n4458), .CLK(n4169), .Q(n_T_427[754]) );
  DFFX1_LVT u_T_427_reg_19__49_ ( .D(n4452), .CLK(n4169), .Q(n_T_427[752]) );
  DFFX1_LVT u_T_427_reg_19__48_ ( .D(n4450), .CLK(n4169), .Q(n_T_427[751]) );
  DFFX1_LVT u_T_427_reg_19__47_ ( .D(n4447), .CLK(n4168), .Q(n_T_427[750]) );
  DFFX1_LVT u_T_427_reg_19__45_ ( .D(n4440), .CLK(n4168), .Q(n_T_427[748]) );
  DFFX1_LVT u_T_427_reg_19__44_ ( .D(n4438), .CLK(n4168), .Q(n_T_427[747]) );
  DFFX1_LVT u_T_427_reg_19__43_ ( .D(n4434), .CLK(n4168), .Q(n_T_427[746]), 
        .QN(n3405) );
  DFFX1_LVT u_T_427_reg_19__42_ ( .D(n4431), .CLK(n4168), .Q(n_T_427[745]) );
  DFFX1_LVT u_T_427_reg_19__41_ ( .D(n4428), .CLK(n4168), .Q(n_T_427[744]) );
  DFFX1_LVT u_T_427_reg_19__39_ ( .D(n4423), .CLK(n4168), .Q(n_T_427[742]) );
  DFFX1_LVT u_T_427_reg_19__38_ ( .D(n4420), .CLK(n4168), .Q(n_T_427[741]) );
  DFFX1_LVT u_T_427_reg_19__37_ ( .D(n4418), .CLK(n4168), .Q(n_T_427[740]) );
  DFFX1_LVT u_T_427_reg_19__36_ ( .D(n4414), .CLK(n4168), .Q(n_T_427[739]) );
  DFFX1_LVT u_T_427_reg_19__33_ ( .D(n4407), .CLK(n4167), .Q(n_T_427[737]) );
  DFFX1_LVT u_T_427_reg_19__31_ ( .D(n4402), .CLK(n4167), .Q(n_T_427[735]) );
  DFFX1_LVT u_T_427_reg_19__30_ ( .D(n4399), .CLK(n4167), .Q(n_T_427[734]) );
  DFFX1_LVT u_T_427_reg_19__29_ ( .D(n4396), .CLK(n4167), .Q(n_T_427[733]) );
  DFFX1_LVT u_T_427_reg_19__28_ ( .D(n4394), .CLK(n4167), .Q(n_T_427[732]) );
  DFFX1_LVT u_T_427_reg_19__27_ ( .D(n4392), .CLK(n4167), .Q(n_T_427[731]) );
  DFFX1_LVT u_T_427_reg_19__26_ ( .D(n4389), .CLK(n4167), .Q(n_T_427[730]) );
  DFFX1_LVT u_T_427_reg_19__25_ ( .D(n4387), .CLK(n4167), .Q(n_T_427[729]) );
  DFFX1_LVT u_T_427_reg_19__24_ ( .D(n4384), .CLK(n4167), .Q(n_T_427[728]) );
  DFFX1_LVT u_T_427_reg_19__23_ ( .D(n4382), .CLK(n4166), .Q(n_T_427[727]) );
  DFFX1_LVT u_T_427_reg_19__22_ ( .D(n4379), .CLK(n4166), .Q(n_T_427[726]) );
  DFFX1_LVT u_T_427_reg_19__21_ ( .D(n4377), .CLK(n4166), .Q(n_T_427[725]) );
  DFFX1_LVT u_T_427_reg_19__20_ ( .D(n4374), .CLK(n4166), .Q(n_T_427[724]) );
  DFFX1_LVT u_T_427_reg_19__19_ ( .D(n4371), .CLK(n4166), .Q(n_T_427[723]) );
  DFFX1_LVT u_T_427_reg_19__18_ ( .D(n4368), .CLK(n4166), .Q(n_T_427[722]) );
  DFFX1_LVT u_T_427_reg_19__17_ ( .D(n4366), .CLK(n4166), .Q(n_T_427[721]) );
  DFFX1_LVT u_T_427_reg_19__16_ ( .D(n4363), .CLK(n4166), .Q(n_T_427[720]) );
  DFFX1_LVT u_T_427_reg_19__15_ ( .D(n4360), .CLK(n4166), .Q(n_T_427[719]) );
  DFFX1_LVT u_T_427_reg_19__14_ ( .D(n4358), .CLK(n4166), .Q(n_T_427[718]) );
  DFFX1_LVT u_T_427_reg_19__13_ ( .D(n4355), .CLK(n4166), .Q(n_T_427[717]) );
  DFFX1_LVT u_T_427_reg_19__12_ ( .D(n4353), .CLK(n4166), .Q(n_T_427[716]) );
  DFFX1_LVT u_T_427_reg_19__11_ ( .D(n4349), .CLK(n4165), .Q(n_T_427[715]) );
  DFFX1_LVT u_T_427_reg_19__10_ ( .D(n4347), .CLK(n4165), .Q(n_T_427[714]) );
  DFFX1_LVT u_T_427_reg_19__9_ ( .D(n4344), .CLK(n4165), .Q(n_T_427[713]) );
  DFFX1_LVT u_T_427_reg_19__8_ ( .D(n4341), .CLK(n4165), .Q(n_T_427[712]) );
  DFFX1_LVT u_T_427_reg_19__7_ ( .D(n4338), .CLK(n4165), .Q(n_T_427[711]) );
  DFFX1_LVT u_T_427_reg_19__6_ ( .D(n4335), .CLK(n4165), .Q(n_T_427[710]) );
  DFFX1_LVT u_T_427_reg_19__5_ ( .D(n4332), .CLK(n4165), .Q(n_T_427[709]) );
  DFFX1_LVT u_T_427_reg_19__4_ ( .D(n4329), .CLK(n4165), .Q(n_T_427[708]) );
  DFFX1_LVT u_T_427_reg_19__3_ ( .D(n4326), .CLK(n4165), .Q(n_T_427[707]) );
  DFFX1_LVT u_T_427_reg_19__2_ ( .D(n4323), .CLK(n4165), .Q(n_T_427[706]) );
  DFFX1_LVT u_T_427_reg_19__1_ ( .D(n4319), .CLK(n4165), .Q(n_T_427[705]) );
  DFFX1_LVT u_T_427_reg_19__0_ ( .D(n4316), .CLK(n4165), .Q(n_T_427[704]) );
  DFFX1_LVT u_T_427_reg_20__63_ ( .D(n4495), .CLK(n4164), .Q(n_T_427[703]) );
  DFFX1_LVT u_T_427_reg_20__62_ ( .D(n4492), .CLK(n4164), .Q(n_T_427[702]), 
        .QN(n3478) );
  DFFX1_LVT u_T_427_reg_20__61_ ( .D(n4489), .CLK(n4164), .Q(n_T_427[701]) );
  DFFX1_LVT u_T_427_reg_20__60_ ( .D(n4486), .CLK(n4164), .Q(n_T_427[700]) );
  DFFX1_LVT u_T_427_reg_20__59_ ( .D(n4483), .CLK(n4163), .Q(n_T_427[699]) );
  DFFX1_LVT u_T_427_reg_20__58_ ( .D(n4479), .CLK(n4163), .Q(n_T_427[698]) );
  DFFX1_LVT u_T_427_reg_20__57_ ( .D(n4477), .CLK(n4163), .Q(n_T_427[697]) );
  DFFX1_LVT u_T_427_reg_20__56_ ( .D(n4473), .CLK(n4163), .Q(n_T_427[696]) );
  DFFX1_LVT u_T_427_reg_20__55_ ( .D(n4471), .CLK(n4163), .Q(n_T_427[695]) );
  DFFX1_LVT u_T_427_reg_20__54_ ( .D(n4467), .CLK(n4163), .Q(n_T_427[694]) );
  DFFX1_LVT u_T_427_reg_20__53_ ( .D(n4465), .CLK(n4163), .Q(n_T_427[693]) );
  DFFX1_LVT u_T_427_reg_20__52_ ( .D(n4461), .CLK(n4163), .Q(n_T_427[692]) );
  DFFX1_LVT u_T_427_reg_20__51_ ( .D(n4458), .CLK(n4163), .Q(n_T_427[691]) );
  DFFX1_LVT u_T_427_reg_20__50_ ( .D(n4456), .CLK(n4163), .Q(n_T_427[690]) );
  DFFX1_LVT u_T_427_reg_20__49_ ( .D(n4452), .CLK(n4163), .Q(n_T_427[689]) );
  DFFX1_LVT u_T_427_reg_20__48_ ( .D(n4450), .CLK(n4163), .Q(n_T_427[688]) );
  DFFX1_LVT u_T_427_reg_20__46_ ( .D(n4444), .CLK(n4162), .Q(n_T_427[686]) );
  DFFX1_LVT u_T_427_reg_20__45_ ( .D(n4440), .CLK(n4162), .Q(n_T_427[685]) );
  DFFX1_LVT u_T_427_reg_20__44_ ( .D(n4438), .CLK(n4162), .Q(n_T_427[684]) );
  DFFX1_LVT u_T_427_reg_20__43_ ( .D(n4434), .CLK(n4162), .Q(n_T_427[683]) );
  DFFX1_LVT u_T_427_reg_20__42_ ( .D(n4431), .CLK(n4162), .Q(n_T_427[682]) );
  DFFX1_LVT u_T_427_reg_20__41_ ( .D(n4428), .CLK(n4162), .Q(n_T_427[681]), 
        .QN(n3404) );
  DFFX1_LVT u_T_427_reg_20__40_ ( .D(n4426), .CLK(n4162), .Q(n_T_427[680]) );
  DFFX1_LVT u_T_427_reg_20__38_ ( .D(n4420), .CLK(n4162), .Q(n_T_427[678]) );
  DFFX1_LVT u_T_427_reg_20__37_ ( .D(n4418), .CLK(n4162), .Q(n_T_427[677]) );
  DFFX1_LVT u_T_427_reg_20__36_ ( .D(n4414), .CLK(n4162), .Q(n_T_427[676]) );
  DFFX1_LVT u_T_427_reg_20__34_ ( .D(n4410), .CLK(n4161), .Q(n_T_427[674]) );
  DFFX1_LVT u_T_427_reg_20__33_ ( .D(n4407), .CLK(n4161), .Q(n_T_427[673]) );
  DFFX1_LVT u_T_427_reg_20__32_ ( .D(n4405), .CLK(n4161), .Q(n_T_427[672]) );
  DFFX1_LVT u_T_427_reg_20__31_ ( .D(n4402), .CLK(n4161), .Q(n_T_427[671]) );
  DFFX1_LVT u_T_427_reg_20__30_ ( .D(n4399), .CLK(n4161), .Q(n_T_427[670]) );
  DFFX1_LVT u_T_427_reg_20__29_ ( .D(n4396), .CLK(n4161), .Q(n_T_427[669]) );
  DFFX1_LVT u_T_427_reg_20__28_ ( .D(n4394), .CLK(n4161), .Q(n_T_427[668]) );
  DFFX1_LVT u_T_427_reg_20__27_ ( .D(n4392), .CLK(n4161), .Q(n_T_427[667]) );
  DFFX1_LVT u_T_427_reg_20__26_ ( .D(n4389), .CLK(n4161), .Q(n_T_427[666]) );
  DFFX1_LVT u_T_427_reg_20__25_ ( .D(n4387), .CLK(n4161), .Q(n_T_427[665]) );
  DFFX1_LVT u_T_427_reg_20__24_ ( .D(n4384), .CLK(n4161), .Q(n_T_427[664]) );
  DFFX1_LVT u_T_427_reg_20__23_ ( .D(n4382), .CLK(n4160), .Q(n_T_427[663]) );
  DFFX1_LVT u_T_427_reg_20__22_ ( .D(n4379), .CLK(n4160), .Q(n_T_427[662]) );
  DFFX1_LVT u_T_427_reg_20__21_ ( .D(n4377), .CLK(n4160), .Q(n_T_427[661]) );
  DFFX1_LVT u_T_427_reg_20__20_ ( .D(n4374), .CLK(n4160), .Q(n_T_427[660]) );
  DFFX1_LVT u_T_427_reg_20__19_ ( .D(n4371), .CLK(n4160), .Q(n_T_427[659]) );
  DFFX1_LVT u_T_427_reg_20__18_ ( .D(n4368), .CLK(n4160), .Q(n_T_427[658]) );
  DFFX1_LVT u_T_427_reg_20__17_ ( .D(n4366), .CLK(n4160), .Q(n_T_427[657]) );
  DFFX1_LVT u_T_427_reg_20__16_ ( .D(n4363), .CLK(n4160), .Q(n_T_427[656]) );
  DFFX1_LVT u_T_427_reg_20__15_ ( .D(n4360), .CLK(n4160), .Q(n_T_427[655]) );
  DFFX1_LVT u_T_427_reg_20__14_ ( .D(n4358), .CLK(n4160), .Q(n_T_427[654]) );
  DFFX1_LVT u_T_427_reg_20__13_ ( .D(n4355), .CLK(n4160), .Q(n_T_427[653]) );
  DFFX1_LVT u_T_427_reg_20__12_ ( .D(n4353), .CLK(n4160), .Q(n_T_427[652]) );
  DFFX1_LVT u_T_427_reg_20__11_ ( .D(n4349), .CLK(n4159), .Q(n_T_427[651]) );
  DFFX1_LVT u_T_427_reg_20__10_ ( .D(n4347), .CLK(n4159), .Q(n_T_427[650]) );
  DFFX1_LVT u_T_427_reg_20__9_ ( .D(n4344), .CLK(n4159), .Q(n_T_427[649]) );
  DFFX1_LVT u_T_427_reg_20__8_ ( .D(n4341), .CLK(n4159), .Q(n_T_427[648]) );
  DFFX1_LVT u_T_427_reg_20__7_ ( .D(n4338), .CLK(n4159), .Q(n_T_427[647]) );
  DFFX1_LVT u_T_427_reg_20__6_ ( .D(n4335), .CLK(n4159), .Q(n_T_427[646]) );
  DFFX1_LVT u_T_427_reg_20__5_ ( .D(n4332), .CLK(n4159), .Q(n_T_427[645]) );
  DFFX1_LVT u_T_427_reg_20__3_ ( .D(n4326), .CLK(n4159), .Q(n_T_427[643]) );
  DFFX1_LVT u_T_427_reg_20__1_ ( .D(n4319), .CLK(n4159), .Q(n_T_427[641]) );
  DFFX1_LVT u_T_427_reg_20__0_ ( .D(n4316), .CLK(n4159), .Q(n_T_427[640]) );
  DFFX1_LVT u_T_427_reg_21__63_ ( .D(n4495), .CLK(n4158), .Q(n_T_427[639]) );
  DFFX1_LVT u_T_427_reg_21__62_ ( .D(n4492), .CLK(n4158), .Q(n_T_427[638]) );
  DFFX1_LVT u_T_427_reg_21__61_ ( .D(n4489), .CLK(n4158), .Q(n_T_427[637]) );
  DFFX1_LVT u_T_427_reg_21__60_ ( .D(n4486), .CLK(n4158), .Q(n_T_427[636]) );
  DFFX1_LVT u_T_427_reg_21__59_ ( .D(n4483), .CLK(n4157), .Q(n_T_427[635]) );
  DFFX1_LVT u_T_427_reg_21__58_ ( .D(n4479), .CLK(n4157), .Q(n_T_427[634]) );
  DFFX1_LVT u_T_427_reg_21__57_ ( .D(n4477), .CLK(n4157), .Q(n_T_427[633]) );
  DFFX1_LVT u_T_427_reg_21__56_ ( .D(n4473), .CLK(n4157), .Q(n_T_427[632]) );
  DFFX1_LVT u_T_427_reg_21__55_ ( .D(n4471), .CLK(n4157), .Q(n_T_427[631]) );
  DFFX1_LVT u_T_427_reg_21__54_ ( .D(n4467), .CLK(n4157), .Q(n_T_427[630]) );
  DFFX1_LVT u_T_427_reg_21__53_ ( .D(n4465), .CLK(n4157), .Q(n_T_427[629]) );
  DFFX1_LVT u_T_427_reg_21__52_ ( .D(n4461), .CLK(n4157), .Q(n_T_427[628]) );
  DFFX1_LVT u_T_427_reg_21__51_ ( .D(n4458), .CLK(n4157), .Q(n_T_427[627]) );
  DFFX1_LVT u_T_427_reg_21__50_ ( .D(n4456), .CLK(n4157), .Q(n_T_427[626]) );
  DFFX1_LVT u_T_427_reg_21__49_ ( .D(n4452), .CLK(n4157), .Q(n_T_427[625]) );
  DFFX1_LVT u_T_427_reg_21__48_ ( .D(n4450), .CLK(n4157), .Q(n_T_427[624]) );
  DFFX1_LVT u_T_427_reg_21__47_ ( .D(n4447), .CLK(n4156), .Q(n_T_427[623]) );
  DFFX1_LVT u_T_427_reg_21__46_ ( .D(n4444), .CLK(n4156), .Q(n_T_427[622]) );
  DFFX1_LVT u_T_427_reg_21__45_ ( .D(n4440), .CLK(n4156), .Q(n_T_427[621]) );
  DFFX1_LVT u_T_427_reg_21__44_ ( .D(n4438), .CLK(n4156), .Q(n_T_427[620]) );
  DFFX1_LVT u_T_427_reg_21__43_ ( .D(n4434), .CLK(n4156), .Q(n_T_427[619]) );
  DFFX1_LVT u_T_427_reg_21__42_ ( .D(n4431), .CLK(n4156), .Q(n_T_427[618]) );
  DFFX1_LVT u_T_427_reg_21__41_ ( .D(n4428), .CLK(n4156), .Q(n_T_427[617]) );
  DFFX1_LVT u_T_427_reg_21__40_ ( .D(n4426), .CLK(n4156), .Q(n_T_427[616]) );
  DFFX1_LVT u_T_427_reg_21__39_ ( .D(n4423), .CLK(n4156), .Q(n_T_427[615]) );
  DFFX1_LVT u_T_427_reg_21__38_ ( .D(n4420), .CLK(n4156), .Q(n_T_427[614]) );
  DFFX1_LVT u_T_427_reg_21__37_ ( .D(n4418), .CLK(n4156), .Q(n_T_427[613]) );
  DFFX1_LVT u_T_427_reg_21__36_ ( .D(n4414), .CLK(n4156), .Q(n_T_427[612]) );
  DFFX1_LVT u_T_427_reg_21__35_ ( .D(n4412), .CLK(n4155), .Q(n_T_427[611]) );
  DFFX1_LVT u_T_427_reg_21__34_ ( .D(n4410), .CLK(n4155), .Q(n_T_427[610]) );
  DFFX1_LVT u_T_427_reg_21__33_ ( .D(n4407), .CLK(n4155), .Q(n_T_427[609]) );
  DFFX1_LVT u_T_427_reg_21__32_ ( .D(n4405), .CLK(n4155), .Q(n_T_427[608]) );
  DFFX1_LVT u_T_427_reg_21__31_ ( .D(n4402), .CLK(n4155), .Q(n_T_427[607]) );
  DFFX1_LVT u_T_427_reg_21__30_ ( .D(n4399), .CLK(n4155), .Q(n_T_427[606]) );
  DFFX1_LVT u_T_427_reg_21__29_ ( .D(n4396), .CLK(n4155), .Q(n_T_427[605]) );
  DFFX1_LVT u_T_427_reg_21__28_ ( .D(n4394), .CLK(n4155), .Q(n_T_427[604]) );
  DFFX1_LVT u_T_427_reg_21__27_ ( .D(n4392), .CLK(n4155), .Q(n_T_427[603]) );
  DFFX1_LVT u_T_427_reg_21__26_ ( .D(n4389), .CLK(n4155), .Q(n_T_427[602]) );
  DFFX1_LVT u_T_427_reg_21__25_ ( .D(n4387), .CLK(n4155), .Q(n_T_427[601]) );
  DFFX1_LVT u_T_427_reg_21__24_ ( .D(n4384), .CLK(n4155), .Q(n_T_427[600]) );
  DFFX1_LVT u_T_427_reg_21__23_ ( .D(n4382), .CLK(n4154), .Q(n_T_427[599]) );
  DFFX1_LVT u_T_427_reg_21__22_ ( .D(n4379), .CLK(n4154), .Q(n_T_427[598]) );
  DFFX1_LVT u_T_427_reg_21__21_ ( .D(n4377), .CLK(n4154), .Q(n_T_427[597]) );
  DFFX1_LVT u_T_427_reg_21__20_ ( .D(n4374), .CLK(n4154), .Q(n_T_427[596]) );
  DFFX1_LVT u_T_427_reg_21__19_ ( .D(n4371), .CLK(n4154), .Q(n_T_427[595]) );
  DFFX1_LVT u_T_427_reg_21__18_ ( .D(n4368), .CLK(n4154), .Q(n_T_427[594]) );
  DFFX1_LVT u_T_427_reg_21__17_ ( .D(n4366), .CLK(n4154), .Q(n_T_427[593]) );
  DFFX1_LVT u_T_427_reg_21__16_ ( .D(n4363), .CLK(n4154), .Q(n_T_427[592]) );
  DFFX1_LVT u_T_427_reg_21__15_ ( .D(n4360), .CLK(n4154), .Q(n_T_427[591]) );
  DFFX1_LVT u_T_427_reg_21__14_ ( .D(n4358), .CLK(n4154), .Q(n_T_427[590]) );
  DFFX1_LVT u_T_427_reg_21__13_ ( .D(n4355), .CLK(n4154), .Q(n_T_427[589]) );
  DFFX1_LVT u_T_427_reg_21__12_ ( .D(n4353), .CLK(n4154), .Q(n_T_427[588]) );
  DFFX1_LVT u_T_427_reg_21__11_ ( .D(n4349), .CLK(n4153), .Q(n_T_427[587]) );
  DFFX1_LVT u_T_427_reg_21__10_ ( .D(n4347), .CLK(n4153), .Q(n_T_427[586]) );
  DFFX1_LVT u_T_427_reg_21__9_ ( .D(n4344), .CLK(n4153), .Q(n_T_427[585]) );
  DFFX1_LVT u_T_427_reg_21__8_ ( .D(n4341), .CLK(n4153), .Q(n_T_427[584]) );
  DFFX1_LVT u_T_427_reg_21__7_ ( .D(n4338), .CLK(n4153), .Q(n_T_427[583]) );
  DFFX1_LVT u_T_427_reg_21__6_ ( .D(n4335), .CLK(n4153), .Q(n_T_427[582]) );
  DFFX1_LVT u_T_427_reg_21__5_ ( .D(n4332), .CLK(n4153), .Q(n_T_427[581]) );
  DFFX1_LVT u_T_427_reg_21__4_ ( .D(n4329), .CLK(n4153), .Q(n_T_427[580]) );
  DFFX1_LVT u_T_427_reg_21__3_ ( .D(n4326), .CLK(n4153), .Q(n_T_427[579]) );
  DFFX1_LVT u_T_427_reg_21__2_ ( .D(n4323), .CLK(n4153), .Q(n_T_427[578]) );
  DFFX1_LVT u_T_427_reg_21__1_ ( .D(n4319), .CLK(n4153), .Q(n_T_427[577]) );
  DFFX1_LVT u_T_427_reg_21__0_ ( .D(n4316), .CLK(n4153), .Q(n_T_427[576]) );
  DFFX1_LVT u_T_427_reg_22__63_ ( .D(n4495), .CLK(n4152), .Q(n_T_427[575]) );
  DFFX1_LVT u_T_427_reg_22__62_ ( .D(n4492), .CLK(n4152), .Q(n_T_427[574]) );
  DFFX1_LVT u_T_427_reg_22__61_ ( .D(n4489), .CLK(n4152), .Q(n_T_427[573]) );
  DFFX1_LVT u_T_427_reg_22__60_ ( .D(n4486), .CLK(n4152), .Q(n_T_427[572]) );
  DFFX1_LVT u_T_427_reg_22__59_ ( .D(n4483), .CLK(n4151), .Q(n_T_427[571]) );
  DFFX1_LVT u_T_427_reg_22__58_ ( .D(n4479), .CLK(n4151), .Q(n_T_427[570]) );
  DFFX1_LVT u_T_427_reg_22__57_ ( .D(n4477), .CLK(n4151), .Q(n_T_427[569]) );
  DFFX1_LVT u_T_427_reg_22__56_ ( .D(n4473), .CLK(n4151), .Q(n_T_427[568]) );
  DFFX1_LVT u_T_427_reg_22__55_ ( .D(n4471), .CLK(n4151), .Q(n_T_427[567]) );
  DFFX1_LVT u_T_427_reg_22__54_ ( .D(n4467), .CLK(n4151), .Q(n_T_427[566]) );
  DFFX1_LVT u_T_427_reg_22__53_ ( .D(n4465), .CLK(n4151), .Q(n_T_427[565]) );
  DFFX1_LVT u_T_427_reg_22__52_ ( .D(n4461), .CLK(n4151), .Q(n_T_427[564]) );
  DFFX1_LVT u_T_427_reg_22__51_ ( .D(n4458), .CLK(n4151), .Q(n_T_427[563]) );
  DFFX1_LVT u_T_427_reg_22__50_ ( .D(n4456), .CLK(n4151), .Q(n_T_427[562]) );
  DFFX1_LVT u_T_427_reg_22__49_ ( .D(n4452), .CLK(n4151), .Q(n_T_427[561]) );
  DFFX1_LVT u_T_427_reg_22__48_ ( .D(n4450), .CLK(n4151), .Q(n_T_427[560]) );
  DFFX1_LVT u_T_427_reg_22__47_ ( .D(n4447), .CLK(n4150), .Q(n_T_427[559]) );
  DFFX1_LVT u_T_427_reg_22__46_ ( .D(n4444), .CLK(n4150), .Q(n_T_427[558]) );
  DFFX1_LVT u_T_427_reg_22__45_ ( .D(n4440), .CLK(n4150), .Q(n_T_427[557]) );
  DFFX1_LVT u_T_427_reg_22__44_ ( .D(n4438), .CLK(n4150), .Q(n_T_427[556]) );
  DFFX1_LVT u_T_427_reg_22__43_ ( .D(n4434), .CLK(n4150), .Q(n_T_427[555]) );
  DFFX1_LVT u_T_427_reg_22__42_ ( .D(n4431), .CLK(n4150), .Q(n_T_427[554]) );
  DFFX1_LVT u_T_427_reg_22__41_ ( .D(n4428), .CLK(n4150), .Q(n_T_427[553]) );
  DFFX1_LVT u_T_427_reg_22__40_ ( .D(n4426), .CLK(n4150), .Q(n_T_427[552]) );
  DFFX1_LVT u_T_427_reg_22__39_ ( .D(n4423), .CLK(n4150), .Q(n_T_427[551]) );
  DFFX1_LVT u_T_427_reg_22__38_ ( .D(n4420), .CLK(n4150), .Q(n_T_427[550]) );
  DFFX1_LVT u_T_427_reg_22__37_ ( .D(n4418), .CLK(n4150), .Q(n_T_427[549]) );
  DFFX1_LVT u_T_427_reg_22__36_ ( .D(n4414), .CLK(n4150), .Q(n_T_427[548]) );
  DFFX1_LVT u_T_427_reg_22__35_ ( .D(n4412), .CLK(n4149), .Q(n_T_427[547]) );
  DFFX1_LVT u_T_427_reg_22__34_ ( .D(n4410), .CLK(n4149), .Q(n_T_427[546]) );
  DFFX1_LVT u_T_427_reg_22__33_ ( .D(n4407), .CLK(n4149), .Q(n_T_427[545]) );
  DFFX1_LVT u_T_427_reg_22__32_ ( .D(n4405), .CLK(n4149), .Q(n_T_427[544]) );
  DFFX1_LVT u_T_427_reg_22__31_ ( .D(n4402), .CLK(n4149), .Q(n_T_427[543]) );
  DFFX1_LVT u_T_427_reg_22__30_ ( .D(n4399), .CLK(n4149), .Q(n_T_427[542]) );
  DFFX1_LVT u_T_427_reg_22__29_ ( .D(n4396), .CLK(n4149), .Q(n_T_427[541]) );
  DFFX1_LVT u_T_427_reg_22__28_ ( .D(n4394), .CLK(n4149), .Q(n_T_427[540]) );
  DFFX1_LVT u_T_427_reg_22__27_ ( .D(n4392), .CLK(n4149), .Q(n_T_427[539]) );
  DFFX1_LVT u_T_427_reg_22__26_ ( .D(n4389), .CLK(n4149), .Q(n_T_427[538]) );
  DFFX1_LVT u_T_427_reg_22__25_ ( .D(n4387), .CLK(n4149), .Q(n_T_427[537]) );
  DFFX1_LVT u_T_427_reg_22__24_ ( .D(n4384), .CLK(n4149), .Q(n_T_427[536]) );
  DFFX1_LVT u_T_427_reg_22__23_ ( .D(n4382), .CLK(n4148), .Q(n_T_427[535]) );
  DFFX1_LVT u_T_427_reg_22__22_ ( .D(n4379), .CLK(n4148), .Q(n_T_427[534]) );
  DFFX1_LVT u_T_427_reg_22__21_ ( .D(n4377), .CLK(n4148), .Q(n_T_427[533]) );
  DFFX1_LVT u_T_427_reg_22__20_ ( .D(n4374), .CLK(n4148), .Q(n_T_427[532]) );
  DFFX1_LVT u_T_427_reg_22__19_ ( .D(n4371), .CLK(n4148), .Q(n_T_427[531]) );
  DFFX1_LVT u_T_427_reg_22__18_ ( .D(n4368), .CLK(n4148), .Q(n_T_427[530]) );
  DFFX1_LVT u_T_427_reg_22__17_ ( .D(n4366), .CLK(n4148), .Q(n_T_427[529]) );
  DFFX1_LVT u_T_427_reg_22__16_ ( .D(n4363), .CLK(n4148), .Q(n_T_427[528]) );
  DFFX1_LVT u_T_427_reg_22__15_ ( .D(n4360), .CLK(n4148), .Q(n_T_427[527]) );
  DFFX1_LVT u_T_427_reg_22__14_ ( .D(n4358), .CLK(n4148), .Q(n_T_427[526]) );
  DFFX1_LVT u_T_427_reg_22__13_ ( .D(n4355), .CLK(n4148), .Q(n_T_427[525]) );
  DFFX1_LVT u_T_427_reg_22__12_ ( .D(n4353), .CLK(n4148), .Q(n_T_427[524]) );
  DFFX1_LVT u_T_427_reg_22__11_ ( .D(n4349), .CLK(n4147), .Q(n_T_427[523]) );
  DFFX1_LVT u_T_427_reg_22__10_ ( .D(n4347), .CLK(n4147), .Q(n_T_427[522]) );
  DFFX1_LVT u_T_427_reg_22__9_ ( .D(n4344), .CLK(n4147), .Q(n_T_427[521]) );
  DFFX1_LVT u_T_427_reg_22__8_ ( .D(n4341), .CLK(n4147), .Q(n_T_427[520]) );
  DFFX1_LVT u_T_427_reg_22__7_ ( .D(n4338), .CLK(n4147), .Q(n_T_427[519]) );
  DFFX1_LVT u_T_427_reg_22__6_ ( .D(n4335), .CLK(n4147), .Q(n_T_427[518]) );
  DFFX1_LVT u_T_427_reg_22__5_ ( .D(n4332), .CLK(n4147), .Q(n_T_427[517]) );
  DFFX1_LVT u_T_427_reg_22__4_ ( .D(n4329), .CLK(n4147), .Q(n_T_427[516]) );
  DFFX1_LVT u_T_427_reg_22__3_ ( .D(n4326), .CLK(n4147), .Q(n_T_427[515]) );
  DFFX1_LVT u_T_427_reg_22__2_ ( .D(n4323), .CLK(n4147), .Q(n_T_427[514]) );
  DFFX1_LVT u_T_427_reg_22__1_ ( .D(n4319), .CLK(n4147), .Q(n_T_427[513]) );
  DFFX1_LVT u_T_427_reg_22__0_ ( .D(n4316), .CLK(n4147), .Q(n_T_427[512]) );
  DFFX1_LVT u_T_427_reg_23__63_ ( .D(n4495), .CLK(n4146), .Q(n_T_427[511]) );
  DFFX1_LVT u_T_427_reg_23__62_ ( .D(n4492), .CLK(n4146), .Q(n_T_427[510]) );
  DFFX1_LVT u_T_427_reg_23__61_ ( .D(n4489), .CLK(n4146), .Q(n_T_427[509]) );
  DFFX1_LVT u_T_427_reg_23__60_ ( .D(n4486), .CLK(n4146), .Q(n_T_427[508]) );
  DFFX1_LVT u_T_427_reg_23__59_ ( .D(n4483), .CLK(n4145), .Q(n_T_427[507]) );
  DFFX1_LVT u_T_427_reg_23__58_ ( .D(n4479), .CLK(n4145), .Q(n_T_427[506]) );
  DFFX1_LVT u_T_427_reg_23__57_ ( .D(n4477), .CLK(n4145), .Q(n_T_427[505]) );
  DFFX1_LVT u_T_427_reg_23__56_ ( .D(n4473), .CLK(n4145), .Q(n_T_427[504]) );
  DFFX1_LVT u_T_427_reg_23__55_ ( .D(n4471), .CLK(n4145), .Q(n_T_427[503]) );
  DFFX1_LVT u_T_427_reg_23__54_ ( .D(n4467), .CLK(n4145), .Q(n_T_427[502]) );
  DFFX1_LVT u_T_427_reg_23__53_ ( .D(n4465), .CLK(n4145), .Q(n_T_427[501]) );
  DFFX1_LVT u_T_427_reg_23__52_ ( .D(n4461), .CLK(n4145), .Q(n_T_427[500]) );
  DFFX1_LVT u_T_427_reg_23__51_ ( .D(n4458), .CLK(n4145), .Q(n_T_427[499]) );
  DFFX1_LVT u_T_427_reg_23__50_ ( .D(n4456), .CLK(n4145), .Q(n_T_427[498]) );
  DFFX1_LVT u_T_427_reg_23__49_ ( .D(n4452), .CLK(n4145), .Q(n_T_427[497]) );
  DFFX1_LVT u_T_427_reg_23__48_ ( .D(n4450), .CLK(n4145), .Q(n_T_427[496]) );
  DFFX1_LVT u_T_427_reg_23__47_ ( .D(n4447), .CLK(n4144), .Q(n_T_427[495]) );
  DFFX1_LVT u_T_427_reg_23__46_ ( .D(n4444), .CLK(n4144), .Q(n_T_427[494]) );
  DFFX1_LVT u_T_427_reg_23__45_ ( .D(n4440), .CLK(n4144), .Q(n_T_427[493]) );
  DFFX1_LVT u_T_427_reg_23__44_ ( .D(n4438), .CLK(n4144), .Q(n_T_427[492]) );
  DFFX1_LVT u_T_427_reg_23__43_ ( .D(n4434), .CLK(n4144), .Q(n_T_427[491]) );
  DFFX1_LVT u_T_427_reg_23__42_ ( .D(n4431), .CLK(n4144), .Q(n_T_427[490]) );
  DFFX1_LVT u_T_427_reg_23__41_ ( .D(n4428), .CLK(n4144), .Q(n_T_427[489]) );
  DFFX1_LVT u_T_427_reg_23__40_ ( .D(n4426), .CLK(n4144), .Q(n_T_427[488]) );
  DFFX1_LVT u_T_427_reg_23__39_ ( .D(n4423), .CLK(n4144), .Q(n_T_427[487]) );
  DFFX1_LVT u_T_427_reg_23__38_ ( .D(n4420), .CLK(n4144), .Q(n_T_427[486]) );
  DFFX1_LVT u_T_427_reg_23__37_ ( .D(n4418), .CLK(n4144), .Q(n_T_427[485]) );
  DFFX1_LVT u_T_427_reg_23__36_ ( .D(n4414), .CLK(n4144), .Q(n_T_427[484]) );
  DFFX1_LVT u_T_427_reg_23__35_ ( .D(n4412), .CLK(n4143), .Q(n_T_427[483]) );
  DFFX1_LVT u_T_427_reg_23__34_ ( .D(n4410), .CLK(n4143), .Q(n_T_427[482]) );
  DFFX1_LVT u_T_427_reg_23__33_ ( .D(n4407), .CLK(n4143), .Q(n_T_427[481]) );
  DFFX1_LVT u_T_427_reg_23__32_ ( .D(n4405), .CLK(n4143), .Q(n_T_427[480]) );
  DFFX1_LVT u_T_427_reg_23__31_ ( .D(n4402), .CLK(n4143), .Q(n_T_427[479]) );
  DFFX1_LVT u_T_427_reg_23__30_ ( .D(n4399), .CLK(n4143), .Q(n_T_427[478]) );
  DFFX1_LVT u_T_427_reg_23__29_ ( .D(n4396), .CLK(n4143), .Q(n_T_427[477]) );
  DFFX1_LVT u_T_427_reg_23__28_ ( .D(n4394), .CLK(n4143), .Q(n_T_427[476]) );
  DFFX1_LVT u_T_427_reg_23__27_ ( .D(n4392), .CLK(n4143), .Q(n_T_427[475]) );
  DFFX1_LVT u_T_427_reg_23__26_ ( .D(n4389), .CLK(n4143), .Q(n_T_427[474]) );
  DFFX1_LVT u_T_427_reg_23__25_ ( .D(n4387), .CLK(n4143), .Q(n_T_427[473]) );
  DFFX1_LVT u_T_427_reg_23__24_ ( .D(n4384), .CLK(n4143), .Q(n_T_427[472]) );
  DFFX1_LVT u_T_427_reg_23__23_ ( .D(n4382), .CLK(n4142), .Q(n_T_427[471]) );
  DFFX1_LVT u_T_427_reg_23__22_ ( .D(n4379), .CLK(n4142), .Q(n_T_427[470]) );
  DFFX1_LVT u_T_427_reg_23__21_ ( .D(n4377), .CLK(n4142), .Q(n_T_427[469]) );
  DFFX1_LVT u_T_427_reg_23__20_ ( .D(n4374), .CLK(n4142), .Q(n_T_427[468]) );
  DFFX1_LVT u_T_427_reg_23__19_ ( .D(n4371), .CLK(n4142), .Q(n_T_427[467]) );
  DFFX1_LVT u_T_427_reg_23__18_ ( .D(n4368), .CLK(n4142), .Q(n_T_427[466]) );
  DFFX1_LVT u_T_427_reg_23__17_ ( .D(n4366), .CLK(n4142), .Q(n_T_427[465]) );
  DFFX1_LVT u_T_427_reg_23__16_ ( .D(n4363), .CLK(n4142), .Q(n_T_427[464]) );
  DFFX1_LVT u_T_427_reg_23__15_ ( .D(n4360), .CLK(n4142), .Q(n_T_427[463]) );
  DFFX1_LVT u_T_427_reg_23__14_ ( .D(n4358), .CLK(n4142), .Q(n_T_427[462]) );
  DFFX1_LVT u_T_427_reg_23__13_ ( .D(n4355), .CLK(n4142), .Q(n_T_427[461]) );
  DFFX1_LVT u_T_427_reg_23__12_ ( .D(n4353), .CLK(n4142), .Q(n_T_427[460]) );
  DFFX1_LVT u_T_427_reg_23__11_ ( .D(n4349), .CLK(n4141), .Q(n_T_427[459]) );
  DFFX1_LVT u_T_427_reg_23__10_ ( .D(n4347), .CLK(n4141), .Q(n_T_427[458]) );
  DFFX1_LVT u_T_427_reg_23__9_ ( .D(n4344), .CLK(n4141), .Q(n_T_427[457]) );
  DFFX1_LVT u_T_427_reg_23__8_ ( .D(n4341), .CLK(n4141), .Q(n_T_427[456]) );
  DFFX1_LVT u_T_427_reg_23__7_ ( .D(n4338), .CLK(n4141), .Q(n_T_427[455]) );
  DFFX1_LVT u_T_427_reg_23__6_ ( .D(n4335), .CLK(n4141), .Q(n_T_427[454]) );
  DFFX1_LVT u_T_427_reg_23__5_ ( .D(n4332), .CLK(n4141), .Q(n_T_427[453]) );
  DFFX1_LVT u_T_427_reg_23__4_ ( .D(n4329), .CLK(n4141), .Q(n_T_427[452]) );
  DFFX1_LVT u_T_427_reg_23__3_ ( .D(n4326), .CLK(n4141), .Q(n_T_427[451]) );
  DFFX1_LVT u_T_427_reg_23__2_ ( .D(n4323), .CLK(n4141), .Q(n_T_427[450]) );
  DFFX1_LVT u_T_427_reg_23__1_ ( .D(n4319), .CLK(n4141), .Q(n_T_427[449]) );
  DFFX1_LVT u_T_427_reg_23__0_ ( .D(n4316), .CLK(n4141), .Q(n_T_427[448]) );
  DFFX1_LVT u_T_427_reg_24__63_ ( .D(n4496), .CLK(n4140), .Q(n_T_427[447]) );
  DFFX1_LVT u_T_427_reg_24__62_ ( .D(n4493), .CLK(n4140), .Q(n_T_427[446]) );
  DFFX1_LVT u_T_427_reg_24__61_ ( .D(n4490), .CLK(n4140), .Q(n_T_427[445]) );
  DFFX1_LVT u_T_427_reg_24__60_ ( .D(n4487), .CLK(n4140), .Q(n_T_427[444]), 
        .QN(n3525) );
  DFFX1_LVT u_T_427_reg_24__59_ ( .D(n4484), .CLK(n4139), .Q(n_T_427[443]) );
  DFFX1_LVT u_T_427_reg_24__58_ ( .D(n4480), .CLK(n4139), .Q(n_T_427[442]) );
  DFFX1_LVT u_T_427_reg_24__57_ ( .D(n4478), .CLK(n4139), .Q(n_T_427[441]) );
  DFFX1_LVT u_T_427_reg_24__56_ ( .D(n4474), .CLK(n4139), .Q(n_T_427[440]) );
  DFFX1_LVT u_T_427_reg_24__55_ ( .D(n4472), .CLK(n4139), .Q(n_T_427[439]) );
  DFFX1_LVT u_T_427_reg_24__54_ ( .D(n4468), .CLK(n4139), .Q(n_T_427[438]) );
  DFFX1_LVT u_T_427_reg_24__53_ ( .D(n4466), .CLK(n4139), .Q(n_T_427[437]) );
  DFFX1_LVT u_T_427_reg_24__52_ ( .D(n4462), .CLK(n4139), .Q(n_T_427[436]) );
  DFFX1_LVT u_T_427_reg_24__51_ ( .D(n4459), .CLK(n4139), .Q(n_T_427[435]) );
  DFFX1_LVT u_T_427_reg_24__50_ ( .D(n4457), .CLK(n4139), .Q(n_T_427[434]) );
  DFFX1_LVT u_T_427_reg_24__49_ ( .D(n4453), .CLK(n4139), .Q(n_T_427[433]) );
  DFFX1_LVT u_T_427_reg_24__48_ ( .D(n4451), .CLK(n4139), .Q(n_T_427[432]) );
  DFFX1_LVT u_T_427_reg_24__47_ ( .D(n4448), .CLK(n4138), .Q(n_T_427[431]) );
  DFFX1_LVT u_T_427_reg_24__46_ ( .D(n4445), .CLK(n4138), .Q(n_T_427[430]) );
  DFFX1_LVT u_T_427_reg_24__45_ ( .D(n4441), .CLK(n4138), .Q(n_T_427[429]) );
  DFFX1_LVT u_T_427_reg_24__44_ ( .D(n4439), .CLK(n4138), .Q(n_T_427[428]) );
  DFFX1_LVT u_T_427_reg_24__43_ ( .D(n4435), .CLK(n4138), .Q(n_T_427[427]) );
  DFFX1_LVT u_T_427_reg_24__42_ ( .D(n4432), .CLK(n4138), .Q(n_T_427[426]) );
  DFFX1_LVT u_T_427_reg_24__41_ ( .D(n4429), .CLK(n4138), .Q(n_T_427[425]) );
  DFFX1_LVT u_T_427_reg_24__40_ ( .D(n4427), .CLK(n4138), .Q(n_T_427[424]) );
  DFFX1_LVT u_T_427_reg_24__39_ ( .D(n4424), .CLK(n4138), .Q(n_T_427[423]) );
  DFFX1_LVT u_T_427_reg_24__38_ ( .D(n4421), .CLK(n4138), .Q(n_T_427[422]) );
  DFFX1_LVT u_T_427_reg_24__37_ ( .D(n4419), .CLK(n4138), .Q(n_T_427[421]) );
  DFFX1_LVT u_T_427_reg_24__36_ ( .D(n4415), .CLK(n4138), .Q(n_T_427[420]) );
  DFFX1_LVT u_T_427_reg_24__35_ ( .D(n4413), .CLK(n4137), .Q(n_T_427[419]) );
  DFFX1_LVT u_T_427_reg_24__34_ ( .D(n4411), .CLK(n4137), .Q(n_T_427[418]), 
        .QN(n3527) );
  DFFX1_LVT u_T_427_reg_24__33_ ( .D(n4408), .CLK(n4137), .Q(n_T_427[417]) );
  DFFX1_LVT u_T_427_reg_24__32_ ( .D(n4406), .CLK(n4137), .Q(n_T_427[416]) );
  DFFX1_LVT u_T_427_reg_24__31_ ( .D(n4403), .CLK(n4137), .Q(n_T_427[415]) );
  DFFX1_LVT u_T_427_reg_24__30_ ( .D(n4400), .CLK(n4137), .Q(n_T_427[414]) );
  DFFX1_LVT u_T_427_reg_24__29_ ( .D(n4397), .CLK(n4137), .Q(n_T_427[413]) );
  DFFX1_LVT u_T_427_reg_24__28_ ( .D(n4395), .CLK(n4137), .Q(n_T_427[412]) );
  DFFX1_LVT u_T_427_reg_24__27_ ( .D(n4393), .CLK(n4137), .Q(n_T_427[411]) );
  DFFX1_LVT u_T_427_reg_24__26_ ( .D(n4390), .CLK(n4137), .Q(n_T_427[410]) );
  DFFX1_LVT u_T_427_reg_24__25_ ( .D(n4388), .CLK(n4137), .Q(n_T_427[409]) );
  DFFX1_LVT u_T_427_reg_24__24_ ( .D(n4385), .CLK(n4137), .Q(n_T_427[408]) );
  DFFX1_LVT u_T_427_reg_24__23_ ( .D(n4383), .CLK(n4136), .Q(n_T_427[407]) );
  DFFX1_LVT u_T_427_reg_24__22_ ( .D(n4380), .CLK(n4136), .Q(n_T_427[406]) );
  DFFX1_LVT u_T_427_reg_24__21_ ( .D(n4378), .CLK(n4136), .Q(n_T_427[405]) );
  DFFX1_LVT u_T_427_reg_24__20_ ( .D(n4375), .CLK(n4136), .Q(n_T_427[404]) );
  DFFX1_LVT u_T_427_reg_24__19_ ( .D(n4372), .CLK(n4136), .Q(n_T_427[403]) );
  DFFX1_LVT u_T_427_reg_24__18_ ( .D(n4369), .CLK(n4136), .Q(n_T_427[402]) );
  DFFX1_LVT u_T_427_reg_24__17_ ( .D(n4367), .CLK(n4136), .Q(n_T_427[401]) );
  DFFX1_LVT u_T_427_reg_24__16_ ( .D(n4364), .CLK(n4136), .Q(n_T_427[400]) );
  DFFX1_LVT u_T_427_reg_24__15_ ( .D(n4361), .CLK(n4136), .Q(n_T_427[399]) );
  DFFX1_LVT u_T_427_reg_24__14_ ( .D(n4359), .CLK(n4136), .Q(n_T_427[398]) );
  DFFX1_LVT u_T_427_reg_24__13_ ( .D(n4356), .CLK(n4136), .Q(n_T_427[397]) );
  DFFX1_LVT u_T_427_reg_24__12_ ( .D(n4354), .CLK(n4136), .Q(n_T_427[396]) );
  DFFX1_LVT u_T_427_reg_24__11_ ( .D(n4349), .CLK(n4135), .Q(n_T_427[395]) );
  DFFX1_LVT u_T_427_reg_24__10_ ( .D(n4348), .CLK(n4135), .Q(n_T_427[394]) );
  DFFX1_LVT u_T_427_reg_24__9_ ( .D(n4345), .CLK(n4135), .Q(n_T_427[393]) );
  DFFX1_LVT u_T_427_reg_24__8_ ( .D(n4342), .CLK(n4135), .Q(n_T_427[392]) );
  DFFX1_LVT u_T_427_reg_24__7_ ( .D(n4339), .CLK(n4135), .Q(n_T_427[391]) );
  DFFX1_LVT u_T_427_reg_24__6_ ( .D(n4336), .CLK(n4135), .Q(n_T_427[390]) );
  DFFX1_LVT u_T_427_reg_24__5_ ( .D(n4333), .CLK(n4135), .Q(n_T_427[389]) );
  DFFX1_LVT u_T_427_reg_24__4_ ( .D(n4330), .CLK(n4135), .Q(n_T_427[388]) );
  DFFX1_LVT u_T_427_reg_24__3_ ( .D(n4327), .CLK(n4135), .Q(n_T_427[387]) );
  DFFX1_LVT u_T_427_reg_24__2_ ( .D(n4324), .CLK(n4135), .Q(n_T_427[386]) );
  DFFX1_LVT u_T_427_reg_24__1_ ( .D(n4320), .CLK(n4135), .Q(n_T_427[385]) );
  DFFX1_LVT u_T_427_reg_24__0_ ( .D(n4317), .CLK(n4135), .Q(n_T_427[384]) );
  DFFX1_LVT u_T_427_reg_25__63_ ( .D(n4496), .CLK(n4134), .Q(n_T_427[383]) );
  DFFX1_LVT u_T_427_reg_25__62_ ( .D(n4493), .CLK(n4134), .Q(n_T_427[382]) );
  DFFX1_LVT u_T_427_reg_25__61_ ( .D(n4490), .CLK(n4134), .Q(n_T_427[381]) );
  DFFX1_LVT u_T_427_reg_25__60_ ( .D(n4487), .CLK(n4134), .Q(n_T_427[380]), 
        .QN(n3172) );
  DFFX1_LVT u_T_427_reg_25__59_ ( .D(n4484), .CLK(n4133), .Q(n_T_427[379]) );
  DFFX1_LVT u_T_427_reg_25__58_ ( .D(n4479), .CLK(n4133), .Q(n_T_427[378]) );
  DFFX1_LVT u_T_427_reg_25__57_ ( .D(n4478), .CLK(n4133), .Q(n_T_427[377]) );
  DFFX1_LVT u_T_427_reg_25__56_ ( .D(n4473), .CLK(n4133), .Q(n_T_427[376]) );
  DFFX1_LVT u_T_427_reg_25__55_ ( .D(n4472), .CLK(n4133), .Q(n_T_427[375]) );
  DFFX1_LVT u_T_427_reg_25__54_ ( .D(n4467), .CLK(n4133), .Q(n_T_427[374]) );
  DFFX1_LVT u_T_427_reg_25__53_ ( .D(n4466), .CLK(n4133), .Q(n_T_427[373]) );
  DFFX1_LVT u_T_427_reg_25__52_ ( .D(n4461), .CLK(n4133), .Q(n_T_427[372]) );
  DFFX1_LVT u_T_427_reg_25__51_ ( .D(n4458), .CLK(n4133), .Q(n_T_427[371]) );
  DFFX1_LVT u_T_427_reg_25__50_ ( .D(n4457), .CLK(n4133), .Q(n_T_427[370]) );
  DFFX1_LVT u_T_427_reg_25__49_ ( .D(n4452), .CLK(n4133), .Q(n_T_427[369]) );
  DFFX1_LVT u_T_427_reg_25__48_ ( .D(n4451), .CLK(n4133), .Q(n_T_427[368]) );
  DFFX1_LVT u_T_427_reg_25__47_ ( .D(n4448), .CLK(n4132), .Q(n_T_427[367]) );
  DFFX1_LVT u_T_427_reg_25__46_ ( .D(n4445), .CLK(n4132), .Q(n_T_427[366]) );
  DFFX1_LVT u_T_427_reg_25__45_ ( .D(n4440), .CLK(n4132), .Q(n_T_427[365]) );
  DFFX1_LVT u_T_427_reg_25__44_ ( .D(n4439), .CLK(n4132), .Q(n_T_427[364]) );
  DFFX1_LVT u_T_427_reg_25__43_ ( .D(n4434), .CLK(n4132), .Q(n_T_427[363]) );
  DFFX1_LVT u_T_427_reg_25__42_ ( .D(n4431), .CLK(n4132), .Q(n_T_427[362]) );
  DFFX1_LVT u_T_427_reg_25__41_ ( .D(n4428), .CLK(n4132), .Q(n_T_427[361]) );
  DFFX1_LVT u_T_427_reg_25__40_ ( .D(n4427), .CLK(n4132), .Q(n_T_427[360]) );
  DFFX1_LVT u_T_427_reg_25__39_ ( .D(n4424), .CLK(n4132), .Q(n_T_427[359]) );
  DFFX1_LVT u_T_427_reg_25__38_ ( .D(n4421), .CLK(n4132), .Q(n_T_427[358]) );
  DFFX1_LVT u_T_427_reg_25__37_ ( .D(n4419), .CLK(n4132), .Q(n_T_427[357]) );
  DFFX1_LVT u_T_427_reg_25__36_ ( .D(n4414), .CLK(n4132), .Q(n_T_427[356]) );
  DFFX1_LVT u_T_427_reg_25__35_ ( .D(n4413), .CLK(n4131), .Q(n_T_427[355]) );
  DFFX1_LVT u_T_427_reg_25__34_ ( .D(n4411), .CLK(n4131), .Q(n_T_427[354]) );
  DFFX1_LVT u_T_427_reg_25__33_ ( .D(n4408), .CLK(n4131), .Q(n_T_427[353]) );
  DFFX1_LVT u_T_427_reg_25__32_ ( .D(n4406), .CLK(n4131), .Q(n_T_427[352]) );
  DFFX1_LVT u_T_427_reg_25__31_ ( .D(n4403), .CLK(n4131), .Q(n_T_427[351]) );
  DFFX1_LVT u_T_427_reg_25__30_ ( .D(n4399), .CLK(n4131), .Q(n_T_427[350]) );
  DFFX1_LVT u_T_427_reg_25__29_ ( .D(n4396), .CLK(n4131), .Q(n_T_427[349]) );
  DFFX1_LVT u_T_427_reg_25__28_ ( .D(n4395), .CLK(n4131), .Q(n_T_427[348]) );
  DFFX1_LVT u_T_427_reg_25__27_ ( .D(n4393), .CLK(n4131), .Q(n_T_427[347]) );
  DFFX1_LVT u_T_427_reg_25__26_ ( .D(n4390), .CLK(n4131), .Q(n_T_427[346]) );
  DFFX1_LVT u_T_427_reg_25__25_ ( .D(n4388), .CLK(n4131), .Q(n_T_427[345]) );
  DFFX1_LVT u_T_427_reg_25__24_ ( .D(n4384), .CLK(n4131), .Q(n_T_427[344]) );
  DFFX1_LVT u_T_427_reg_25__23_ ( .D(n4383), .CLK(n4130), .Q(n_T_427[343]) );
  DFFX1_LVT u_T_427_reg_25__22_ ( .D(n4380), .CLK(n4130), .Q(n_T_427[342]) );
  DFFX1_LVT u_T_427_reg_25__21_ ( .D(n4378), .CLK(n4130), .Q(n_T_427[341]) );
  DFFX1_LVT u_T_427_reg_25__20_ ( .D(n4374), .CLK(n4130), .Q(n_T_427[340]) );
  DFFX1_LVT u_T_427_reg_25__19_ ( .D(n4371), .CLK(n4130), .Q(n_T_427[339]) );
  DFFX1_LVT u_T_427_reg_25__18_ ( .D(n4368), .CLK(n4130), .Q(n_T_427[338]) );
  DFFX1_LVT u_T_427_reg_25__17_ ( .D(n4367), .CLK(n4130), .Q(n_T_427[337]) );
  DFFX1_LVT u_T_427_reg_25__16_ ( .D(n4364), .CLK(n4130), .Q(n_T_427[336]) );
  DFFX1_LVT u_T_427_reg_25__15_ ( .D(n4361), .CLK(n4130), .Q(n_T_427[335]) );
  DFFX1_LVT u_T_427_reg_25__14_ ( .D(n4359), .CLK(n4130), .Q(n_T_427[334]) );
  DFFX1_LVT u_T_427_reg_25__13_ ( .D(n4356), .CLK(n4130), .Q(n_T_427[333]) );
  DFFX1_LVT u_T_427_reg_25__12_ ( .D(n4354), .CLK(n4130), .Q(n_T_427[332]) );
  DFFX1_LVT u_T_427_reg_25__11_ ( .D(n4349), .CLK(n4129), .Q(n_T_427[331]) );
  DFFX1_LVT u_T_427_reg_25__10_ ( .D(n4348), .CLK(n4129), .Q(n_T_427[330]) );
  DFFX1_LVT u_T_427_reg_25__9_ ( .D(n4345), .CLK(n4129), .Q(n_T_427[329]) );
  DFFX1_LVT u_T_427_reg_25__8_ ( .D(n4342), .CLK(n4129), .Q(n_T_427[328]) );
  DFFX1_LVT u_T_427_reg_25__7_ ( .D(n4339), .CLK(n4129), .Q(n_T_427[327]) );
  DFFX1_LVT u_T_427_reg_25__6_ ( .D(n4336), .CLK(n4129), .Q(n_T_427[326]) );
  DFFX1_LVT u_T_427_reg_25__5_ ( .D(n4333), .CLK(n4129), .Q(n_T_427[325]) );
  DFFX1_LVT u_T_427_reg_25__4_ ( .D(n4330), .CLK(n4129), .Q(n_T_427[324]), 
        .QN(n3520) );
  DFFX1_LVT u_T_427_reg_25__3_ ( .D(n4327), .CLK(n4129), .Q(n_T_427[323]) );
  DFFX1_LVT u_T_427_reg_25__2_ ( .D(n4324), .CLK(n4129), .Q(n_T_427[322]), 
        .QN(n3519) );
  DFFX1_LVT u_T_427_reg_25__1_ ( .D(n4319), .CLK(n4129), .Q(n_T_427[321]) );
  DFFX1_LVT u_T_427_reg_25__0_ ( .D(n4316), .CLK(n4129), .Q(n_T_427[320]) );
  DFFX1_LVT u_T_427_reg_26__63_ ( .D(n4496), .CLK(n4128), .Q(n_T_427[319]) );
  DFFX1_LVT u_T_427_reg_26__62_ ( .D(n4493), .CLK(n4128), .Q(n_T_427[318]) );
  DFFX1_LVT u_T_427_reg_26__61_ ( .D(n4490), .CLK(n4128), .Q(n_T_427[317]) );
  DFFX1_LVT u_T_427_reg_26__60_ ( .D(n4487), .CLK(n4128), .Q(n_T_427[316]) );
  DFFX1_LVT u_T_427_reg_26__59_ ( .D(n4484), .CLK(n4127), .Q(n_T_427[315]) );
  DFFX1_LVT u_T_427_reg_26__58_ ( .D(n4479), .CLK(n4127), .Q(n_T_427[314]) );
  DFFX1_LVT u_T_427_reg_26__57_ ( .D(n4478), .CLK(n4127), .Q(n_T_427[313]) );
  DFFX1_LVT u_T_427_reg_26__56_ ( .D(n4473), .CLK(n4127), .Q(n_T_427[312]) );
  DFFX1_LVT u_T_427_reg_26__55_ ( .D(n4472), .CLK(n4127), .Q(n_T_427[311]) );
  DFFX1_LVT u_T_427_reg_26__54_ ( .D(n4467), .CLK(n4127), .Q(n_T_427[310]) );
  DFFX1_LVT u_T_427_reg_26__53_ ( .D(n4466), .CLK(n4127), .Q(n_T_427[309]) );
  DFFX1_LVT u_T_427_reg_26__52_ ( .D(n4461), .CLK(n4127), .Q(n_T_427[308]) );
  DFFX1_LVT u_T_427_reg_26__51_ ( .D(n4458), .CLK(n4127), .Q(n_T_427[307]) );
  DFFX1_LVT u_T_427_reg_26__50_ ( .D(n4457), .CLK(n4127), .Q(n_T_427[306]) );
  DFFX1_LVT u_T_427_reg_26__49_ ( .D(n4452), .CLK(n4127), .Q(n_T_427[305]) );
  DFFX1_LVT u_T_427_reg_26__48_ ( .D(n4451), .CLK(n4127), .Q(n_T_427[304]) );
  DFFX1_LVT u_T_427_reg_26__47_ ( .D(n4448), .CLK(n4126), .Q(n_T_427[303]) );
  DFFX1_LVT u_T_427_reg_26__46_ ( .D(n4445), .CLK(n4126), .Q(n_T_427[302]) );
  DFFX1_LVT u_T_427_reg_26__45_ ( .D(n4440), .CLK(n4126), .Q(n_T_427[301]) );
  DFFX1_LVT u_T_427_reg_26__44_ ( .D(n4439), .CLK(n4126), .Q(n_T_427[300]) );
  DFFX1_LVT u_T_427_reg_26__43_ ( .D(n4434), .CLK(n4126), .Q(n_T_427[299]) );
  DFFX1_LVT u_T_427_reg_26__42_ ( .D(n4431), .CLK(n4126), .Q(n_T_427[298]) );
  DFFX1_LVT u_T_427_reg_26__41_ ( .D(n4428), .CLK(n4126), .Q(n_T_427[297]) );
  DFFX1_LVT u_T_427_reg_26__40_ ( .D(n4427), .CLK(n4126), .Q(n_T_427[296]) );
  DFFX1_LVT u_T_427_reg_26__39_ ( .D(n4424), .CLK(n4126), .Q(n_T_427[295]) );
  DFFX1_LVT u_T_427_reg_26__38_ ( .D(n4421), .CLK(n4126), .Q(n_T_427[294]) );
  DFFX1_LVT u_T_427_reg_26__37_ ( .D(n4419), .CLK(n4126), .Q(n_T_427[293]) );
  DFFX1_LVT u_T_427_reg_26__36_ ( .D(n4414), .CLK(n4126), .Q(n_T_427[292]) );
  DFFX1_LVT u_T_427_reg_26__35_ ( .D(n4413), .CLK(n4125), .Q(n_T_427[291]) );
  DFFX1_LVT u_T_427_reg_26__34_ ( .D(n4411), .CLK(n4125), .Q(n_T_427[290]) );
  DFFX1_LVT u_T_427_reg_26__33_ ( .D(n4408), .CLK(n4125), .Q(n_T_427[289]) );
  DFFX1_LVT u_T_427_reg_26__32_ ( .D(n4406), .CLK(n4125), .Q(n_T_427[288]) );
  DFFX1_LVT u_T_427_reg_26__31_ ( .D(n4403), .CLK(n4125), .Q(n_T_427[287]) );
  DFFX1_LVT u_T_427_reg_26__30_ ( .D(n4399), .CLK(n4125), .Q(n_T_427[286]) );
  DFFX1_LVT u_T_427_reg_26__29_ ( .D(n4396), .CLK(n4125), .Q(n_T_427[285]) );
  DFFX1_LVT u_T_427_reg_26__28_ ( .D(n4395), .CLK(n4125), .Q(n_T_427[284]) );
  DFFX1_LVT u_T_427_reg_26__27_ ( .D(n4393), .CLK(n4125), .Q(n_T_427[283]) );
  DFFX1_LVT u_T_427_reg_26__26_ ( .D(n4390), .CLK(n4125), .Q(n_T_427[282]) );
  DFFX1_LVT u_T_427_reg_26__25_ ( .D(n4388), .CLK(n4125), .Q(n_T_427[281]) );
  DFFX1_LVT u_T_427_reg_26__24_ ( .D(n4384), .CLK(n4125), .Q(n_T_427[280]) );
  DFFX1_LVT u_T_427_reg_26__23_ ( .D(n4383), .CLK(n4124), .Q(n_T_427[279]) );
  DFFX1_LVT u_T_427_reg_26__22_ ( .D(n4380), .CLK(n4124), .Q(n_T_427[278]) );
  DFFX1_LVT u_T_427_reg_26__21_ ( .D(n4378), .CLK(n4124), .Q(n_T_427[277]) );
  DFFX1_LVT u_T_427_reg_26__20_ ( .D(n4374), .CLK(n4124), .Q(n_T_427[276]) );
  DFFX1_LVT u_T_427_reg_26__19_ ( .D(n4371), .CLK(n4124), .Q(n_T_427[275]) );
  DFFX1_LVT u_T_427_reg_26__18_ ( .D(n4368), .CLK(n4124), .Q(n_T_427[274]) );
  DFFX1_LVT u_T_427_reg_26__17_ ( .D(n4367), .CLK(n4124), .Q(n_T_427[273]) );
  DFFX1_LVT u_T_427_reg_26__16_ ( .D(n4364), .CLK(n4124), .Q(n_T_427[272]) );
  DFFX1_LVT u_T_427_reg_26__15_ ( .D(n4361), .CLK(n4124), .Q(n_T_427[271]) );
  DFFX1_LVT u_T_427_reg_26__14_ ( .D(n4359), .CLK(n4124), .Q(n_T_427[270]) );
  DFFX1_LVT u_T_427_reg_26__13_ ( .D(n4356), .CLK(n4124), .Q(n_T_427[269]) );
  DFFX1_LVT u_T_427_reg_26__12_ ( .D(n4354), .CLK(n4124), .Q(n_T_427[268]) );
  DFFX1_LVT u_T_427_reg_26__11_ ( .D(n4349), .CLK(n4123), .Q(n_T_427[267]) );
  DFFX1_LVT u_T_427_reg_26__10_ ( .D(n4348), .CLK(n4123), .Q(n_T_427[266]) );
  DFFX1_LVT u_T_427_reg_26__9_ ( .D(n4345), .CLK(n4123), .Q(n_T_427[265]) );
  DFFX1_LVT u_T_427_reg_26__8_ ( .D(n4342), .CLK(n4123), .Q(n_T_427[264]) );
  DFFX1_LVT u_T_427_reg_26__7_ ( .D(n4339), .CLK(n4123), .Q(n_T_427[263]) );
  DFFX1_LVT u_T_427_reg_26__6_ ( .D(n4336), .CLK(n4123), .Q(n_T_427[262]) );
  DFFX1_LVT u_T_427_reg_26__5_ ( .D(n4333), .CLK(n4123), .Q(n_T_427[261]) );
  DFFX1_LVT u_T_427_reg_26__4_ ( .D(n4330), .CLK(n4123), .Q(n_T_427[260]) );
  DFFX1_LVT u_T_427_reg_26__3_ ( .D(n4327), .CLK(n4123), .Q(n_T_427[259]) );
  DFFX1_LVT u_T_427_reg_26__2_ ( .D(n4324), .CLK(n4123), .Q(n_T_427[258]) );
  DFFX1_LVT u_T_427_reg_26__1_ ( .D(n4319), .CLK(n4123), .Q(n_T_427[257]) );
  DFFX1_LVT u_T_427_reg_26__0_ ( .D(n4316), .CLK(n4123), .Q(n_T_427[256]) );
  DFFX1_LVT u_T_427_reg_27__63_ ( .D(n4496), .CLK(n4122), .Q(n_T_427[255]) );
  DFFX1_LVT u_T_427_reg_27__62_ ( .D(n4493), .CLK(n4122), .Q(n_T_427[254]) );
  DFFX1_LVT u_T_427_reg_27__61_ ( .D(n4490), .CLK(n4122), .Q(n_T_427[253]) );
  DFFX1_LVT u_T_427_reg_27__60_ ( .D(n4487), .CLK(n4122), .Q(n_T_427[252]) );
  DFFX1_LVT u_T_427_reg_27__59_ ( .D(n4484), .CLK(n4121), .Q(n_T_427[251]) );
  DFFX1_LVT u_T_427_reg_27__58_ ( .D(n4479), .CLK(n4121), .Q(n_T_427[250]) );
  DFFX1_LVT u_T_427_reg_27__57_ ( .D(n4478), .CLK(n4121), .Q(n_T_427[249]) );
  DFFX1_LVT u_T_427_reg_27__56_ ( .D(n4473), .CLK(n4121), .Q(n_T_427[248]) );
  DFFX1_LVT u_T_427_reg_27__55_ ( .D(n4472), .CLK(n4121), .Q(n_T_427[247]) );
  DFFX1_LVT u_T_427_reg_27__54_ ( .D(n4467), .CLK(n4121), .Q(n_T_427[246]) );
  DFFX1_LVT u_T_427_reg_27__53_ ( .D(n4466), .CLK(n4121), .Q(n_T_427[245]) );
  DFFX1_LVT u_T_427_reg_27__52_ ( .D(n4461), .CLK(n4121), .Q(n_T_427[244]) );
  DFFX1_LVT u_T_427_reg_27__51_ ( .D(n4458), .CLK(n4121), .Q(n_T_427[243]) );
  DFFX1_LVT u_T_427_reg_27__50_ ( .D(n4457), .CLK(n4121), .Q(n_T_427[242]) );
  DFFX1_LVT u_T_427_reg_27__49_ ( .D(n4452), .CLK(n4121), .Q(n_T_427[241]) );
  DFFX1_LVT u_T_427_reg_27__48_ ( .D(n4451), .CLK(n4121), .Q(n_T_427[240]) );
  DFFX1_LVT u_T_427_reg_27__47_ ( .D(n4448), .CLK(n4120), .Q(n_T_427[239]) );
  DFFX1_LVT u_T_427_reg_27__46_ ( .D(n4445), .CLK(n4120), .Q(n_T_427[238]), 
        .QN(n3522) );
  DFFX1_LVT u_T_427_reg_27__45_ ( .D(n4440), .CLK(n4120), .Q(n_T_427[237]) );
  DFFX1_LVT u_T_427_reg_27__44_ ( .D(n4439), .CLK(n4120), .Q(n_T_427[236]) );
  DFFX1_LVT u_T_427_reg_27__43_ ( .D(n4434), .CLK(n4120), .Q(n_T_427[235]) );
  DFFX1_LVT u_T_427_reg_27__42_ ( .D(n4431), .CLK(n4120), .Q(n_T_427[234]) );
  DFFX1_LVT u_T_427_reg_27__41_ ( .D(n4428), .CLK(n4120), .Q(n_T_427[233]) );
  DFFX1_LVT u_T_427_reg_27__40_ ( .D(n4427), .CLK(n4120), .Q(n_T_427[232]) );
  DFFX1_LVT u_T_427_reg_27__39_ ( .D(n4424), .CLK(n4120), .Q(n_T_427[231]), 
        .QN(n3523) );
  DFFX1_LVT u_T_427_reg_27__38_ ( .D(n4421), .CLK(n4120), .Q(n_T_427[230]) );
  DFFX1_LVT u_T_427_reg_27__37_ ( .D(n4419), .CLK(n4120), .Q(n_T_427[229]) );
  DFFX1_LVT u_T_427_reg_27__36_ ( .D(n4414), .CLK(n4120), .Q(n_T_427[228]) );
  DFFX1_LVT u_T_427_reg_27__35_ ( .D(n4413), .CLK(n4119), .Q(n_T_427[227]) );
  DFFX1_LVT u_T_427_reg_27__34_ ( .D(n4411), .CLK(n4119), .Q(n_T_427[226]) );
  DFFX1_LVT u_T_427_reg_27__33_ ( .D(n4408), .CLK(n4119), .Q(n_T_427[225]) );
  DFFX1_LVT u_T_427_reg_27__32_ ( .D(n4406), .CLK(n4119), .Q(n_T_427[224]) );
  DFFX1_LVT u_T_427_reg_27__31_ ( .D(n4403), .CLK(n4119), .Q(n_T_427[223]) );
  DFFX1_LVT u_T_427_reg_27__30_ ( .D(n4399), .CLK(n4119), .Q(n_T_427[222]) );
  DFFX1_LVT u_T_427_reg_27__29_ ( .D(n4396), .CLK(n4119), .Q(n_T_427[221]) );
  DFFX1_LVT u_T_427_reg_27__28_ ( .D(n4395), .CLK(n4119), .Q(n_T_427[220]) );
  DFFX1_LVT u_T_427_reg_27__27_ ( .D(n4393), .CLK(n4119), .Q(n_T_427[219]) );
  DFFX1_LVT u_T_427_reg_27__26_ ( .D(n4390), .CLK(n4119), .Q(n_T_427[218]) );
  DFFX1_LVT u_T_427_reg_27__25_ ( .D(n4388), .CLK(n4119), .Q(n_T_427[217]) );
  DFFX1_LVT u_T_427_reg_27__24_ ( .D(n4384), .CLK(n4119), .Q(n_T_427[216]) );
  DFFX1_LVT u_T_427_reg_27__23_ ( .D(n4383), .CLK(n4118), .Q(n_T_427[215]) );
  DFFX1_LVT u_T_427_reg_27__22_ ( .D(n4380), .CLK(n4118), .Q(n_T_427[214]) );
  DFFX1_LVT u_T_427_reg_27__21_ ( .D(n4378), .CLK(n4118), .Q(n_T_427[213]) );
  DFFX1_LVT u_T_427_reg_27__20_ ( .D(n4374), .CLK(n4118), .Q(n_T_427[212]) );
  DFFX1_LVT u_T_427_reg_27__19_ ( .D(n4371), .CLK(n4118), .Q(n_T_427[211]) );
  DFFX1_LVT u_T_427_reg_27__18_ ( .D(n4368), .CLK(n4118), .Q(n_T_427[210]) );
  DFFX1_LVT u_T_427_reg_27__17_ ( .D(n4367), .CLK(n4118), .Q(n_T_427[209]) );
  DFFX1_LVT u_T_427_reg_27__16_ ( .D(n4364), .CLK(n4118), .Q(n_T_427[208]), 
        .QN(n3521) );
  DFFX1_LVT u_T_427_reg_27__15_ ( .D(n4361), .CLK(n4118), .Q(n_T_427[207]) );
  DFFX1_LVT u_T_427_reg_27__14_ ( .D(n4359), .CLK(n4118), .Q(n_T_427[206]) );
  DFFX1_LVT u_T_427_reg_27__13_ ( .D(n4356), .CLK(n4118), .Q(n_T_427[205]) );
  DFFX1_LVT u_T_427_reg_27__12_ ( .D(n4354), .CLK(n4118), .Q(n_T_427[204]) );
  DFFX1_LVT u_T_427_reg_27__11_ ( .D(n4349), .CLK(n4117), .Q(n_T_427[203]) );
  DFFX1_LVT u_T_427_reg_27__10_ ( .D(n4348), .CLK(n4117), .Q(n_T_427[202]) );
  DFFX1_LVT u_T_427_reg_27__9_ ( .D(n4345), .CLK(n4117), .Q(n_T_427[201]) );
  DFFX1_LVT u_T_427_reg_27__8_ ( .D(n4342), .CLK(n4117), .Q(n_T_427[200]) );
  DFFX1_LVT u_T_427_reg_27__7_ ( .D(n4339), .CLK(n4117), .Q(n_T_427[199]) );
  DFFX1_LVT u_T_427_reg_27__6_ ( .D(n4336), .CLK(n4117), .Q(n_T_427[198]) );
  DFFX1_LVT u_T_427_reg_27__5_ ( .D(n4333), .CLK(n4117), .Q(n_T_427[197]) );
  DFFX1_LVT u_T_427_reg_27__4_ ( .D(n4330), .CLK(n4117), .Q(n_T_427[196]) );
  DFFX1_LVT u_T_427_reg_27__3_ ( .D(n4327), .CLK(n4117), .Q(n_T_427[195]) );
  DFFX1_LVT u_T_427_reg_27__2_ ( .D(n4324), .CLK(n4117), .Q(n_T_427[194]) );
  DFFX1_LVT u_T_427_reg_27__1_ ( .D(n4319), .CLK(n4117), .Q(n_T_427[193]) );
  DFFX1_LVT u_T_427_reg_27__0_ ( .D(n4316), .CLK(n4117), .Q(n_T_427[192]) );
  DFFX1_LVT u_T_427_reg_28__63_ ( .D(n4496), .CLK(n4116), .Q(n_T_427[191]) );
  DFFX1_LVT u_T_427_reg_28__62_ ( .D(n4493), .CLK(n4116), .Q(n_T_427[190]) );
  DFFX1_LVT u_T_427_reg_28__61_ ( .D(n4490), .CLK(n4116), .Q(n_T_427[189]) );
  DFFX1_LVT u_T_427_reg_28__60_ ( .D(n4487), .CLK(n4116), .Q(n_T_427[188]) );
  DFFX1_LVT u_T_427_reg_28__59_ ( .D(n4484), .CLK(n4115), .Q(n_T_427[187]) );
  DFFX1_LVT u_T_427_reg_28__58_ ( .D(n4479), .CLK(n4115), .Q(n_T_427[186]) );
  DFFX1_LVT u_T_427_reg_28__57_ ( .D(n4478), .CLK(n4115), .Q(n_T_427[185]) );
  DFFX1_LVT u_T_427_reg_28__56_ ( .D(n4473), .CLK(n4115), .Q(n_T_427[184]) );
  DFFX1_LVT u_T_427_reg_28__55_ ( .D(n4472), .CLK(n4115), .Q(n_T_427[183]) );
  DFFX1_LVT u_T_427_reg_28__54_ ( .D(n4467), .CLK(n4115), .Q(n_T_427[182]) );
  DFFX1_LVT u_T_427_reg_28__53_ ( .D(n4466), .CLK(n4115), .Q(n_T_427[181]) );
  DFFX1_LVT u_T_427_reg_28__52_ ( .D(n4461), .CLK(n4115), .Q(n_T_427[180]) );
  DFFX1_LVT u_T_427_reg_28__51_ ( .D(n4458), .CLK(n4115), .Q(n_T_427[179]) );
  DFFX1_LVT u_T_427_reg_28__50_ ( .D(n4457), .CLK(n4115), .Q(n_T_427[178]) );
  DFFX1_LVT u_T_427_reg_28__49_ ( .D(n4452), .CLK(n4115), .Q(n_T_427[177]) );
  DFFX1_LVT u_T_427_reg_28__48_ ( .D(n4451), .CLK(n4115), .Q(n_T_427[176]) );
  DFFX1_LVT u_T_427_reg_28__47_ ( .D(n4448), .CLK(n4114), .Q(n_T_427[175]) );
  DFFX1_LVT u_T_427_reg_28__46_ ( .D(n4445), .CLK(n4114), .Q(n_T_427[174]) );
  DFFX1_LVT u_T_427_reg_28__45_ ( .D(n4440), .CLK(n4114), .Q(n_T_427[173]) );
  DFFX1_LVT u_T_427_reg_28__44_ ( .D(n4439), .CLK(n4114), .Q(n_T_427[172]) );
  DFFX1_LVT u_T_427_reg_28__43_ ( .D(n4434), .CLK(n4114), .Q(n_T_427[171]) );
  DFFX1_LVT u_T_427_reg_28__42_ ( .D(n4431), .CLK(n4114), .Q(n_T_427[170]) );
  DFFX1_LVT u_T_427_reg_28__41_ ( .D(n4428), .CLK(n4114), .Q(n_T_427[169]) );
  DFFX1_LVT u_T_427_reg_28__40_ ( .D(n4427), .CLK(n4114), .Q(n_T_427[168]) );
  DFFX1_LVT u_T_427_reg_28__39_ ( .D(n4424), .CLK(n4114), .Q(n_T_427[167]) );
  DFFX1_LVT u_T_427_reg_28__38_ ( .D(n4421), .CLK(n4114), .Q(n_T_427[166]) );
  DFFX1_LVT u_T_427_reg_28__37_ ( .D(n4419), .CLK(n4114), .Q(n_T_427[165]) );
  DFFX1_LVT u_T_427_reg_28__36_ ( .D(n4414), .CLK(n4114), .Q(n_T_427[164]) );
  DFFX1_LVT u_T_427_reg_28__35_ ( .D(n4413), .CLK(n4113), .Q(n_T_427[163]) );
  DFFX1_LVT u_T_427_reg_28__34_ ( .D(n4411), .CLK(n4113), .Q(n_T_427[162]) );
  DFFX1_LVT u_T_427_reg_28__33_ ( .D(n4408), .CLK(n4113), .Q(n_T_427[161]) );
  DFFX1_LVT u_T_427_reg_28__32_ ( .D(n4406), .CLK(n4113), .Q(n_T_427[160]) );
  DFFX1_LVT u_T_427_reg_28__31_ ( .D(n4403), .CLK(n4113), .Q(n_T_427[159]) );
  DFFX1_LVT u_T_427_reg_28__30_ ( .D(n4399), .CLK(n4113), .Q(n_T_427[158]) );
  DFFX1_LVT u_T_427_reg_28__29_ ( .D(n4396), .CLK(n4113), .Q(n_T_427[157]) );
  DFFX1_LVT u_T_427_reg_28__28_ ( .D(n4395), .CLK(n4113), .Q(n_T_427[156]) );
  DFFX1_LVT u_T_427_reg_28__27_ ( .D(n4393), .CLK(n4113), .Q(n_T_427[155]) );
  DFFX1_LVT u_T_427_reg_28__26_ ( .D(n4390), .CLK(n4113), .Q(n_T_427[154]) );
  DFFX1_LVT u_T_427_reg_28__25_ ( .D(n4388), .CLK(n4113), .Q(n_T_427[153]) );
  DFFX1_LVT u_T_427_reg_28__24_ ( .D(n4384), .CLK(n4113), .Q(n_T_427[152]) );
  DFFX1_LVT u_T_427_reg_28__23_ ( .D(n4383), .CLK(n4112), .Q(n_T_427[151]), 
        .QN(n3526) );
  DFFX1_LVT u_T_427_reg_28__22_ ( .D(n4380), .CLK(n4112), .Q(n_T_427[150]) );
  DFFX1_LVT u_T_427_reg_28__21_ ( .D(n4378), .CLK(n4112), .Q(n_T_427[149]) );
  DFFX1_LVT u_T_427_reg_28__20_ ( .D(n4374), .CLK(n4112), .Q(n_T_427[148]) );
  DFFX1_LVT u_T_427_reg_28__19_ ( .D(n4371), .CLK(n4112), .Q(n_T_427[147]) );
  DFFX1_LVT u_T_427_reg_28__18_ ( .D(n4368), .CLK(n4112), .Q(n_T_427[146]) );
  DFFX1_LVT u_T_427_reg_28__17_ ( .D(n4367), .CLK(n4112), .Q(n_T_427[145]) );
  DFFX1_LVT u_T_427_reg_28__16_ ( .D(n4364), .CLK(n4112), .Q(n_T_427[144]) );
  DFFX1_LVT u_T_427_reg_28__15_ ( .D(n4361), .CLK(n4112), .Q(n_T_427[143]) );
  DFFX1_LVT u_T_427_reg_28__14_ ( .D(n4359), .CLK(n4112), .Q(n_T_427[142]) );
  DFFX1_LVT u_T_427_reg_28__13_ ( .D(n4356), .CLK(n4112), .Q(n_T_427[141]) );
  DFFX1_LVT u_T_427_reg_28__12_ ( .D(n4354), .CLK(n4112), .Q(n_T_427[140]) );
  DFFX1_LVT u_T_427_reg_28__11_ ( .D(n4349), .CLK(n4111), .Q(n_T_427[139]) );
  DFFX1_LVT u_T_427_reg_28__10_ ( .D(n4348), .CLK(n4111), .Q(n_T_427[138]) );
  DFFX1_LVT u_T_427_reg_28__9_ ( .D(n4345), .CLK(n4111), .Q(n_T_427[137]) );
  DFFX1_LVT u_T_427_reg_28__8_ ( .D(n4342), .CLK(n4111), .Q(n_T_427[136]) );
  DFFX1_LVT u_T_427_reg_28__7_ ( .D(n4339), .CLK(n4111), .Q(n_T_427[135]) );
  DFFX1_LVT u_T_427_reg_28__6_ ( .D(n4336), .CLK(n4111), .Q(n_T_427[134]) );
  DFFX1_LVT u_T_427_reg_28__5_ ( .D(n4333), .CLK(n4111), .Q(n_T_427[133]) );
  DFFX1_LVT u_T_427_reg_28__4_ ( .D(n4330), .CLK(n4111), .Q(n_T_427[132]) );
  DFFX1_LVT u_T_427_reg_28__3_ ( .D(n4327), .CLK(n4111), .Q(n_T_427[131]) );
  DFFX1_LVT u_T_427_reg_28__2_ ( .D(n4324), .CLK(n4111), .Q(n_T_427[130]) );
  DFFX1_LVT u_T_427_reg_28__1_ ( .D(n4319), .CLK(n4111), .Q(n_T_427[129]) );
  DFFX1_LVT u_T_427_reg_28__0_ ( .D(n4316), .CLK(n4111), .Q(n_T_427[128]) );
  DFFX1_LVT u_T_427_reg_29__63_ ( .D(n4496), .CLK(n4110), .Q(n_T_427[127]) );
  DFFX1_LVT u_T_427_reg_29__62_ ( .D(n4493), .CLK(n4110), .Q(n_T_427[126]) );
  DFFX1_LVT u_T_427_reg_29__61_ ( .D(n4490), .CLK(n4110), .Q(n_T_427[125]) );
  DFFX1_LVT u_T_427_reg_29__60_ ( .D(n4487), .CLK(n4110), .Q(n_T_427[124]) );
  DFFX1_LVT u_T_427_reg_29__59_ ( .D(n4484), .CLK(n4109), .Q(n_T_427[123]) );
  DFFX1_LVT u_T_427_reg_29__58_ ( .D(n4479), .CLK(n4109), .Q(n_T_427[122]) );
  DFFX1_LVT u_T_427_reg_29__57_ ( .D(n4478), .CLK(n4109), .Q(n_T_427[121]) );
  DFFX1_LVT u_T_427_reg_29__56_ ( .D(n4473), .CLK(n4109), .Q(n_T_427[120]) );
  DFFX1_LVT u_T_427_reg_29__55_ ( .D(n4472), .CLK(n4109), .Q(n_T_427[119]) );
  DFFX1_LVT u_T_427_reg_29__54_ ( .D(n4467), .CLK(n4109), .Q(n_T_427[118]) );
  DFFX1_LVT u_T_427_reg_29__53_ ( .D(n4466), .CLK(n4109), .Q(n_T_427[117]) );
  DFFX1_LVT u_T_427_reg_29__52_ ( .D(n4461), .CLK(n4109), .Q(n_T_427[116]) );
  DFFX1_LVT u_T_427_reg_29__51_ ( .D(n4458), .CLK(n4109), .Q(n_T_427[115]) );
  DFFX1_LVT u_T_427_reg_29__50_ ( .D(n4457), .CLK(n4109), .Q(n_T_427[114]) );
  DFFX1_LVT u_T_427_reg_29__49_ ( .D(n4452), .CLK(n4109), .Q(n_T_427[113]) );
  DFFX1_LVT u_T_427_reg_29__48_ ( .D(n4451), .CLK(n4109), .Q(n_T_427[112]) );
  DFFX1_LVT u_T_427_reg_29__47_ ( .D(n4448), .CLK(n4108), .Q(n_T_427[111]) );
  DFFX1_LVT u_T_427_reg_29__46_ ( .D(n4445), .CLK(n4108), .Q(n_T_427[110]), 
        .QN(n3176) );
  DFFX1_LVT u_T_427_reg_29__45_ ( .D(n4440), .CLK(n4108), .Q(n_T_427[109]) );
  DFFX1_LVT u_T_427_reg_29__44_ ( .D(n4439), .CLK(n4108), .Q(n_T_427[108]) );
  DFFX1_LVT u_T_427_reg_29__43_ ( .D(n4434), .CLK(n4108), .Q(n_T_427[107]) );
  DFFX1_LVT u_T_427_reg_29__42_ ( .D(n4431), .CLK(n4108), .Q(n_T_427[106]) );
  DFFX1_LVT u_T_427_reg_29__41_ ( .D(n4428), .CLK(n4108), .Q(n_T_427[105]) );
  DFFX1_LVT u_T_427_reg_29__40_ ( .D(n4427), .CLK(n4108), .Q(n_T_427[104]) );
  DFFX1_LVT u_T_427_reg_29__39_ ( .D(n4424), .CLK(n4108), .Q(n_T_427[103]) );
  DFFX1_LVT u_T_427_reg_29__38_ ( .D(n4421), .CLK(n4108), .Q(n_T_427[102]) );
  DFFX1_LVT u_T_427_reg_29__37_ ( .D(n4419), .CLK(n4108), .Q(n_T_427[101]) );
  DFFX1_LVT u_T_427_reg_29__36_ ( .D(n4414), .CLK(n4108), .Q(n_T_427[100]) );
  DFFX1_LVT u_T_427_reg_29__35_ ( .D(n4413), .CLK(n4107), .Q(n_T_427[99]) );
  DFFX1_LVT u_T_427_reg_29__34_ ( .D(n4411), .CLK(n4107), .Q(n_T_427[98]) );
  DFFX1_LVT u_T_427_reg_29__33_ ( .D(n4408), .CLK(n4107), .Q(n_T_427[97]) );
  DFFX1_LVT u_T_427_reg_29__32_ ( .D(n4406), .CLK(n4107), .Q(n_T_427[96]) );
  DFFX1_LVT u_T_427_reg_29__31_ ( .D(n4403), .CLK(n4107), .Q(n_T_427[95]) );
  DFFX1_LVT u_T_427_reg_29__30_ ( .D(n4399), .CLK(n4107), .Q(n_T_427[94]) );
  DFFX1_LVT u_T_427_reg_29__29_ ( .D(n4396), .CLK(n4107), .Q(n_T_427[93]) );
  DFFX1_LVT u_T_427_reg_29__28_ ( .D(n4395), .CLK(n4107), .Q(n_T_427[92]) );
  DFFX1_LVT u_T_427_reg_29__27_ ( .D(n4393), .CLK(n4107), .Q(n_T_427[91]) );
  DFFX1_LVT u_T_427_reg_29__26_ ( .D(n4390), .CLK(n4107), .Q(n_T_427[90]) );
  DFFX1_LVT u_T_427_reg_29__25_ ( .D(n4388), .CLK(n4107), .Q(n_T_427[89]) );
  DFFX1_LVT u_T_427_reg_29__24_ ( .D(n4384), .CLK(n4107), .Q(n_T_427[88]) );
  DFFX1_LVT u_T_427_reg_29__23_ ( .D(n4383), .CLK(n4106), .Q(n_T_427[87]) );
  DFFX1_LVT u_T_427_reg_29__22_ ( .D(n4380), .CLK(n4106), .Q(n_T_427[86]) );
  DFFX1_LVT u_T_427_reg_29__21_ ( .D(n4378), .CLK(n4106), .Q(n_T_427[85]) );
  DFFX1_LVT u_T_427_reg_29__20_ ( .D(n4374), .CLK(n4106), .Q(n_T_427[84]) );
  DFFX1_LVT u_T_427_reg_29__19_ ( .D(n4371), .CLK(n4106), .Q(n_T_427[83]) );
  DFFX1_LVT u_T_427_reg_29__18_ ( .D(n4368), .CLK(n4106), .Q(n_T_427[82]) );
  DFFX1_LVT u_T_427_reg_29__17_ ( .D(n4367), .CLK(n4106), .Q(n_T_427[81]) );
  DFFX1_LVT u_T_427_reg_29__16_ ( .D(n4364), .CLK(n4106), .Q(n_T_427[80]), 
        .QN(n3175) );
  DFFX1_LVT u_T_427_reg_29__15_ ( .D(n4361), .CLK(n4106), .Q(n_T_427[79]) );
  DFFX1_LVT u_T_427_reg_29__14_ ( .D(n4359), .CLK(n4106), .Q(n_T_427[78]) );
  DFFX1_LVT u_T_427_reg_29__13_ ( .D(n4356), .CLK(n4106), .Q(n_T_427[77]) );
  DFFX1_LVT u_T_427_reg_29__12_ ( .D(n4354), .CLK(n4106), .Q(n_T_427[76]) );
  DFFX1_LVT u_T_427_reg_29__11_ ( .D(n4349), .CLK(n4105), .Q(n_T_427[75]) );
  DFFX1_LVT u_T_427_reg_29__10_ ( .D(n4348), .CLK(n4105), .Q(n_T_427[74]) );
  DFFX1_LVT u_T_427_reg_29__9_ ( .D(n4345), .CLK(n4105), .Q(n_T_427[73]) );
  DFFX1_LVT u_T_427_reg_29__8_ ( .D(n4342), .CLK(n4105), .Q(n_T_427[72]) );
  DFFX1_LVT u_T_427_reg_29__7_ ( .D(n4339), .CLK(n4105), .Q(n_T_427[71]) );
  DFFX1_LVT u_T_427_reg_29__6_ ( .D(n4336), .CLK(n4105), .Q(n_T_427[70]) );
  DFFX1_LVT u_T_427_reg_29__5_ ( .D(n4333), .CLK(n4105), .Q(n_T_427[69]) );
  DFFX1_LVT u_T_427_reg_29__4_ ( .D(n4330), .CLK(n4105), .Q(n_T_427[68]) );
  DFFX1_LVT u_T_427_reg_29__3_ ( .D(n4327), .CLK(n4105), .Q(n_T_427[67]) );
  DFFX1_LVT u_T_427_reg_29__2_ ( .D(n4324), .CLK(n4105), .Q(n_T_427[66]) );
  DFFX1_LVT u_T_427_reg_29__1_ ( .D(n4319), .CLK(n4105), .Q(n_T_427[65]) );
  DFFX1_LVT u_T_427_reg_29__0_ ( .D(n4316), .CLK(n4105), .Q(n_T_427[64]) );
  DFFX1_LVT u_T_427_reg_30__63_ ( .D(n4496), .CLK(n4104), .Q(n_T_427[63]) );
  DFFX1_LVT u_T_427_reg_30__62_ ( .D(n4493), .CLK(n4104), .Q(n_T_427[62]) );
  DFFX1_LVT u_T_427_reg_30__61_ ( .D(n4490), .CLK(n4104), .Q(n_T_427[61]) );
  DFFX1_LVT u_T_427_reg_30__60_ ( .D(n4487), .CLK(n4104), .Q(n_T_427[60]) );
  DFFX1_LVT u_T_427_reg_30__59_ ( .D(n4484), .CLK(n4103), .Q(n_T_427[59]) );
  DFFX1_LVT u_T_427_reg_30__58_ ( .D(n4479), .CLK(n4103), .Q(n_T_427[58]) );
  DFFX1_LVT u_T_427_reg_30__57_ ( .D(n4478), .CLK(n4103), .Q(n_T_427[57]) );
  DFFX1_LVT u_T_427_reg_30__56_ ( .D(n4473), .CLK(n4103), .Q(n_T_427[56]) );
  DFFX1_LVT u_T_427_reg_30__55_ ( .D(n4472), .CLK(n4103), .Q(n_T_427[55]) );
  DFFX1_LVT u_T_427_reg_30__54_ ( .D(n4467), .CLK(n4103), .Q(n_T_427[54]) );
  DFFX1_LVT u_T_427_reg_30__53_ ( .D(n4466), .CLK(n4103), .Q(n_T_427[53]) );
  DFFX1_LVT u_T_427_reg_30__52_ ( .D(n4461), .CLK(n4103), .Q(n_T_427[52]) );
  DFFX1_LVT u_T_427_reg_30__51_ ( .D(n4458), .CLK(n4103), .Q(n_T_427[51]) );
  DFFX1_LVT u_T_427_reg_30__50_ ( .D(n4457), .CLK(n4103), .Q(n_T_427[50]) );
  DFFX1_LVT u_T_427_reg_30__49_ ( .D(n4452), .CLK(n4103), .Q(n_T_427[49]) );
  DFFX1_LVT u_T_427_reg_30__48_ ( .D(n4451), .CLK(n4103), .Q(n_T_427[48]) );
  DFFX1_LVT u_T_427_reg_30__47_ ( .D(n4448), .CLK(n4102), .Q(n_T_427[47]) );
  DFFX1_LVT u_T_427_reg_30__46_ ( .D(n4445), .CLK(n4102), .Q(n_T_427[46]) );
  DFFX1_LVT u_T_427_reg_30__45_ ( .D(n4440), .CLK(n4102), .Q(n_T_427[45]) );
  DFFX1_LVT u_T_427_reg_30__44_ ( .D(n4439), .CLK(n4102), .Q(n_T_427[44]) );
  DFFX1_LVT u_T_427_reg_30__43_ ( .D(n4434), .CLK(n4102), .Q(n_T_427[43]) );
  DFFX1_LVT u_T_427_reg_30__42_ ( .D(n4431), .CLK(n4102), .Q(n_T_427[42]) );
  DFFX1_LVT u_T_427_reg_30__41_ ( .D(n4428), .CLK(n4102), .Q(n_T_427[41]) );
  DFFX1_LVT u_T_427_reg_30__40_ ( .D(n4427), .CLK(n4102), .Q(n_T_427[40]) );
  DFFX1_LVT u_T_427_reg_30__39_ ( .D(n4424), .CLK(n4102), .Q(n_T_427[39]) );
  DFFX1_LVT u_T_427_reg_30__38_ ( .D(n4421), .CLK(n4102), .Q(n_T_427[38]) );
  DFFX1_LVT u_T_427_reg_30__37_ ( .D(n4419), .CLK(n4102), .Q(n_T_427[37]) );
  DFFX1_LVT u_T_427_reg_30__36_ ( .D(n4414), .CLK(n4102), .Q(n_T_427[36]) );
  DFFX1_LVT u_T_427_reg_30__35_ ( .D(n4413), .CLK(n4101), .Q(n_T_427[35]) );
  DFFX1_LVT u_T_427_reg_30__34_ ( .D(n4411), .CLK(n4101), .Q(n_T_427[34]) );
  DFFX1_LVT u_T_427_reg_30__33_ ( .D(n4408), .CLK(n4101), .Q(n_T_427[33]) );
  DFFX1_LVT u_T_427_reg_30__32_ ( .D(n4406), .CLK(n4101), .Q(n_T_427[32]) );
  DFFX1_LVT u_T_427_reg_30__31_ ( .D(n4403), .CLK(n4101), .Q(n_T_427[31]) );
  DFFX1_LVT u_T_427_reg_30__30_ ( .D(n4399), .CLK(n4101), .Q(n_T_427[30]) );
  DFFX1_LVT u_T_427_reg_30__29_ ( .D(n4396), .CLK(n4101), .Q(n_T_427[29]) );
  DFFX1_LVT u_T_427_reg_30__28_ ( .D(n4395), .CLK(n4101), .Q(n_T_427[28]) );
  DFFX1_LVT u_T_427_reg_30__27_ ( .D(n4393), .CLK(n4101), .Q(n_T_427[27]) );
  DFFX1_LVT u_T_427_reg_30__26_ ( .D(n4390), .CLK(n4101), .Q(n_T_427[26]) );
  DFFX1_LVT u_T_427_reg_30__25_ ( .D(n4388), .CLK(n4101), .Q(n_T_427[25]) );
  DFFX1_LVT u_T_427_reg_30__24_ ( .D(n4384), .CLK(n4101), .Q(n_T_427[24]) );
  DFFX1_LVT u_T_427_reg_30__23_ ( .D(n4383), .CLK(n4100), .Q(n_T_427[23]), 
        .QN(n3177) );
  DFFX1_LVT u_T_427_reg_30__22_ ( .D(n4380), .CLK(n4100), .Q(n_T_427[22]) );
  DFFX1_LVT u_T_427_reg_30__21_ ( .D(n4378), .CLK(n4100), .Q(n_T_427[21]) );
  DFFX1_LVT u_T_427_reg_30__20_ ( .D(n4374), .CLK(n4100), .Q(n_T_427[20]) );
  DFFX1_LVT u_T_427_reg_30__19_ ( .D(n4371), .CLK(n4100), .Q(n_T_427[19]) );
  DFFX1_LVT u_T_427_reg_30__18_ ( .D(n4368), .CLK(n4100), .Q(n_T_427[18]) );
  DFFX1_LVT u_T_427_reg_30__17_ ( .D(n4367), .CLK(n4100), .Q(n_T_427[17]) );
  DFFX1_LVT u_T_427_reg_30__16_ ( .D(n4364), .CLK(n4100), .Q(n_T_427[16]) );
  DFFX1_LVT u_T_427_reg_30__15_ ( .D(n4361), .CLK(n4100), .Q(n_T_427[15]) );
  DFFX1_LVT u_T_427_reg_30__14_ ( .D(n4359), .CLK(n4100), .Q(n_T_427[14]) );
  DFFX1_LVT u_T_427_reg_30__13_ ( .D(n4356), .CLK(n4100), .Q(n_T_427[13]) );
  DFFX1_LVT u_T_427_reg_30__12_ ( .D(n4354), .CLK(n4100), .Q(n_T_427[12]) );
  DFFX1_LVT u_T_427_reg_30__11_ ( .D(n4349), .CLK(n4099), .Q(n_T_427[11]) );
  DFFX1_LVT u_T_427_reg_30__10_ ( .D(n4348), .CLK(n4099), .Q(n_T_427[10]) );
  DFFX1_LVT u_T_427_reg_30__9_ ( .D(n4345), .CLK(n4099), .Q(n_T_427[9]) );
  DFFX1_LVT u_T_427_reg_30__8_ ( .D(n4342), .CLK(n4099), .Q(n_T_427[8]) );
  DFFX1_LVT u_T_427_reg_30__7_ ( .D(n4339), .CLK(n4099), .Q(n_T_427[7]) );
  DFFX1_LVT u_T_427_reg_30__6_ ( .D(n4336), .CLK(n4099), .Q(n_T_427[6]) );
  DFFX1_LVT u_T_427_reg_30__5_ ( .D(n4333), .CLK(n4099), .Q(n_T_427[5]) );
  DFFX1_LVT u_T_427_reg_30__4_ ( .D(n4330), .CLK(n4099), .Q(n_T_427[4]) );
  DFFX1_LVT u_T_427_reg_30__3_ ( .D(n4327), .CLK(n4099), .Q(n_T_427[3]) );
  DFFX1_LVT u_T_427_reg_30__2_ ( .D(n4324), .CLK(n4099), .Q(n_T_427[2]) );
  DFFX1_LVT u_T_427_reg_30__1_ ( .D(n4319), .CLK(n4099), .Q(n_T_427[1]) );
  DFFX1_LVT u_T_427_reg_30__0_ ( .D(n4316), .CLK(n4099), .Q(n_T_427[0]) );
  DFFX1_LVT u_T_1185_reg_31_ ( .D(N777), .CLK(n4071), .Q(n_T_1187[31]), .QN(
        n3267) );
  DFFX1_LVT u_T_1185_reg_30_ ( .D(N776), .CLK(n4071), .Q(n_T_1187[30]) );
  DFFX1_LVT u_T_1185_reg_29_ ( .D(N775), .CLK(n4071), .Q(n_T_1187[29]), .QN(
        n3131) );
  DFFX1_LVT u_T_1185_reg_28_ ( .D(N774), .CLK(n4071), .Q(n_T_1187[28]), .QN(
        n3274) );
  DFFX1_LVT u_T_1185_reg_26_ ( .D(N772), .CLK(n4071), .Q(n_T_1187[26]), .QN(
        n3265) );
  DFFX1_LVT u_T_1185_reg_25_ ( .D(N771), .CLK(n4071), .Q(n_T_1187[25]), .QN(
        n3089) );
  DFFX1_LVT u_T_1185_reg_24_ ( .D(N770), .CLK(n4071), .Q(n_T_1187[24]), .QN(
        n3275) );
  DFFX1_LVT u_T_1185_reg_23_ ( .D(N769), .CLK(n4071), .Q(n_T_1187[23]), .QN(
        n3268) );
  DFFX1_LVT u_T_1185_reg_22_ ( .D(N768), .CLK(n4071), .Q(n_T_1187[22]) );
  DFFX1_LVT u_T_1185_reg_21_ ( .D(N767), .CLK(n4071), .Q(n_T_1187[21]), .QN(
        n3130) );
  DFFX1_LVT u_T_1185_reg_20_ ( .D(N766), .CLK(n4071), .Q(n_T_1187[20]), .QN(
        n3273) );
  DFFX1_LVT u_T_1185_reg_19_ ( .D(N765), .CLK(n4072), .Q(n_T_1187[19]), .QN(
        n3258) );
  DFFX1_LVT u_T_1185_reg_18_ ( .D(N764), .CLK(n4072), .Q(n_T_1187[18]), .QN(
        n3263) );
  DFFX1_LVT u_T_1185_reg_17_ ( .D(N763), .CLK(n4072), .Q(n_T_1187[17]), .QN(
        n3113) );
  DFFX1_LVT u_T_1185_reg_16_ ( .D(N762), .CLK(n4072), .Q(n_T_1187[16]), .QN(
        n3261) );
  DFFX1_LVT u_T_1185_reg_15_ ( .D(N761), .CLK(n4072), .Q(n_T_1187[15]), .QN(
        n3266) );
  DFFX1_LVT u_T_1185_reg_14_ ( .D(N760), .CLK(n4072), .Q(n_T_1187[14]), .QN(
        n3127) );
  DFFX1_LVT u_T_1185_reg_13_ ( .D(N759), .CLK(n4072), .Q(n_T_1187[13]), .QN(
        n3272) );
  DFFX1_LVT u_T_1185_reg_12_ ( .D(N758), .CLK(n4072), .Q(n_T_1187[12]), .QN(
        n3260) );
  DFFX1_LVT u_T_1185_reg_11_ ( .D(N757), .CLK(n4072), .Q(n_T_1187[11]), .QN(
        n3259) );
  DFFX1_LVT u_T_1185_reg_10_ ( .D(N756), .CLK(n4072), .Q(n_T_1187[10]), .QN(
        n3129) );
  DFFX1_LVT u_T_1185_reg_9_ ( .D(N755), .CLK(n4072), .Q(n_T_1187[9]), .QN(
        n3133) );
  DFFX1_LVT u_T_1185_reg_8_ ( .D(N754), .CLK(n4072), .Q(n_T_1187[8]), .QN(
        n3134) );
  DFFX1_LVT u_T_1185_reg_7_ ( .D(N753), .CLK(n4073), .Q(n_T_1187[7]), .QN(
        n3270) );
  DFFX1_LVT u_T_1185_reg_6_ ( .D(N752), .CLK(n4073), .Q(n_T_1187[6]), .QN(
        n3136) );
  DFFX1_LVT u_T_1185_reg_5_ ( .D(N751), .CLK(n4073), .Q(n_T_1187[5]), .QN(
        n3271) );
  DFFX1_LVT u_T_1185_reg_4_ ( .D(N750), .CLK(n4073), .Q(n_T_1187[4]), .QN(
        n3132) );
  DFFX1_LVT u_T_1185_reg_3_ ( .D(N749), .CLK(n4073), .Q(n_T_1187[3]), .QN(
        n3269) );
  DFFX1_LVT u_T_1185_reg_2_ ( .D(N748), .CLK(n4073), .Q(n_T_1187[2]), .QN(
        n3264) );
  DFFX1_LVT u_T_1185_reg_1_ ( .D(N747), .CLK(n4073), .Q(n_T_1187[1]), .QN(
        n3128) );
  DFFX1_LVT u_T_1298_reg_31_ ( .D(N810), .CLK(n4068), .Q(n_T_1298[31]), .QN(
        n3241) );
  DFFX1_LVT u_T_1298_reg_30_ ( .D(N809), .CLK(n4068), .Q(n_T_1298[30]), .QN(
        n3118) );
  DFFX1_LVT u_T_1298_reg_29_ ( .D(N808), .CLK(n4068), .Q(n_T_1298[29]), .QN(
        n3084) );
  DFFX1_LVT u_T_1298_reg_28_ ( .D(N807), .CLK(n4068), .Q(n_T_1298[28]), .QN(
        n3123) );
  DFFX1_LVT u_T_1298_reg_27_ ( .D(N806), .CLK(n4068), .Q(n_T_1298[27]), .QN(
        n3085) );
  DFFX1_LVT u_T_1298_reg_26_ ( .D(N805), .CLK(n4068), .Q(n_T_1298[26]), .QN(
        n3232) );
  DFFX1_LVT u_T_1298_reg_25_ ( .D(N804), .CLK(n4068), .Q(n_T_1298[25]), .QN(
        n3116) );
  DFFX1_LVT u_T_1298_reg_24_ ( .D(N803), .CLK(n4068), .Q(n_T_1298[24]), .QN(
        n3237) );
  DFFX1_LVT u_T_1298_reg_23_ ( .D(N802), .CLK(n4068), .Q(n_T_1298[23]), .QN(
        n3239) );
  DFFX1_LVT u_T_1298_reg_22_ ( .D(N801), .CLK(n4068), .Q(n_T_1298[22]), .QN(
        n3117) );
  DFFX1_LVT u_T_1298_reg_21_ ( .D(N800), .CLK(n4068), .Q(n_T_1298[21]), .QN(
        n3114) );
  DFFX1_LVT u_T_1298_reg_20_ ( .D(N799), .CLK(n4068), .Q(n_T_1298[20]), .QN(
        n3238) );
  DFFX1_LVT u_T_1298_reg_19_ ( .D(N798), .CLK(n4069), .Q(n_T_1298[19]), .QN(
        n3126) );
  DFFX1_LVT u_T_1298_reg_18_ ( .D(N797), .CLK(n4069), .Q(n_T_1298[18]), .QN(
        n3250) );
  DFFX1_LVT u_T_1298_reg_17_ ( .D(N796), .CLK(n4069), .Q(n_T_1298[17]), .QN(
        n3087) );
  DFFX1_LVT u_T_1298_reg_16_ ( .D(N795), .CLK(n4069), .Q(n_T_1298[16]), .QN(
        n3252) );
  DFFX1_LVT u_T_1298_reg_15_ ( .D(N794), .CLK(n4069), .Q(n_T_1298[15]), .QN(
        n3236) );
  DFFX1_LVT u_T_1298_reg_14_ ( .D(N793), .CLK(n4069), .Q(n_T_1298[14]), .QN(
        n3121) );
  DFFX1_LVT u_T_1298_reg_13_ ( .D(N792), .CLK(n4069), .Q(n_T_1298[13]), .QN(
        n3120) );
  DFFX1_LVT u_T_1298_reg_12_ ( .D(N791), .CLK(n4069), .Q(n_T_1298[12]), .QN(
        n3235) );
  DFFX1_LVT u_T_1298_reg_11_ ( .D(N790), .CLK(n4069), .Q(n_T_1298[11]), .QN(
        n3240) );
  DFFX1_LVT u_T_1298_reg_10_ ( .D(N789), .CLK(n4069), .Q(n_T_1298[10]), .QN(
        n3115) );
  DFFX1_LVT u_T_1298_reg_9_ ( .D(N788), .CLK(n4069), .Q(n_T_1298[9]), .QN(
        n3119) );
  DFFX1_LVT u_T_1298_reg_8_ ( .D(N787), .CLK(n4069), .Q(n_T_1298[8]), .QN(
        n3242) );
  DFFX1_LVT u_T_1298_reg_7_ ( .D(N786), .CLK(n4070), .Q(n_T_1298[7]), .QN(
        n3125) );
  DFFX1_LVT u_T_1298_reg_6_ ( .D(N785), .CLK(n4070), .Q(n_T_1298[6]), .QN(
        n3248) );
  DFFX1_LVT u_T_1298_reg_5_ ( .D(N784), .CLK(n4070), .Q(n_T_1298[5]), .QN(
        n3088) );
  DFFX1_LVT u_T_1298_reg_4_ ( .D(N783), .CLK(n4070), .Q(n_T_1298[4]), .QN(
        n3253) );
  DFFX1_LVT u_T_1298_reg_3_ ( .D(N782), .CLK(n4070), .Q(n_T_1298[3]), .QN(
        n3124) );
  DFFX1_LVT u_T_1298_reg_2_ ( .D(N781), .CLK(n4070), .Q(n_T_1298[2]), .QN(
        n3247) );
  DFFX1_LVT u_T_1298_reg_1_ ( .D(N780), .CLK(n4070), .Q(n_T_1298[1]), .QN(
        n3086) );
  DFFX1_LVT u_T_1298_reg_0_ ( .D(N779), .CLK(n4070), .Q(n_T_1298[0]), .QN(
        n3254) );
  AO22X1_LVT U613 ( .A1(csr_io_pc[0]), .A2(n4062), .A3(1'b0), .A4(n4065), .Y(
        io_imem_req_bits_pc[0]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_61_ ( .D(N743), .CLK(n4085), .Q(n_T_628[63])
         );
  DFFX1_LVT ex_reg_mem_size_reg_1_ ( .D(N370), .CLK(n4314), .Q(
        io_dmem_req_bits_size[1]), .QN(n586) );
  DFFX1_LVT u_T_427_reg_0__50_ ( .D(n4455), .CLK(n4283), .QN(n3277) );
  DFFX1_LVT u_T_427_reg_0__32_ ( .D(n4404), .CLK(n4281), .QN(n3276) );
  DFFX1_LVT u_T_427_reg_19__34_ ( .D(n4410), .CLK(n4167), .QN(n3141) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_39_ ( .D(N721), .CLK(n4083), .Q(n_T_628[41])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_53_ ( .D(N735), .CLK(n4084), .Q(n_T_628[55])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_33_ ( .D(N715), .CLK(n4082), .Q(n_T_628[35])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_56_ ( .D(N738), .CLK(n4084), .Q(n_T_628[58])
         );
  DFFX1_LVT u_T_427_reg_0__55_ ( .D(n4470), .CLK(n4283), .Q(n_T_427[1934]), 
        .QN(n3563) );
  DFFX1_LVT u_T_427_reg_0__53_ ( .D(n4464), .CLK(n4283), .Q(n_T_427[1932]), 
        .QN(n3561) );
  DFFX1_LVT u_T_427_reg_0__48_ ( .D(n4449), .CLK(n4283), .Q(n_T_427[1928]), 
        .QN(n3557) );
  DFFX1_LVT u_T_427_reg_0__47_ ( .D(n4446), .CLK(n4282), .Q(n_T_427[1927]), 
        .QN(n3556) );
  DFFX1_LVT u_T_427_reg_0__40_ ( .D(n4425), .CLK(n4282), .Q(n_T_427[1920]), 
        .QN(n3551) );
  DFFX1_LVT u_T_427_reg_0__37_ ( .D(n4417), .CLK(n4282), .Q(n_T_427[1917]), 
        .QN(n3550) );
  DFFX1_LVT u_T_427_reg_3__17_ ( .D(n4365), .CLK(n4262), .Q(n_T_427[1744]), 
        .QN(n3541) );
  DFFX1_LVT u_T_427_reg_0__17_ ( .D(n4365), .CLK(n4280), .Q(n_T_427[1898]), 
        .QN(n3540) );
  DFFX1_LVT u_T_427_reg_0__15_ ( .D(n4360), .CLK(n4280), .Q(n_T_427[1896]), 
        .QN(n3539) );
  DFFX1_LVT u_T_427_reg_0__13_ ( .D(n4355), .CLK(n4280), .Q(n_T_427[1894]), 
        .QN(n3538) );
  DFFX1_LVT u_T_427_reg_0__12_ ( .D(n4352), .CLK(n4280), .Q(n_T_427[1893]), 
        .QN(n3537) );
  DFFX1_LVT u_T_427_reg_0__10_ ( .D(n4346), .CLK(n4279), .Q(n_T_427[1891]), 
        .QN(n3536) );
  DFFX1_LVT u_T_427_reg_0__9_ ( .D(n4343), .CLK(n4279), .Q(n_T_427[1890]), 
        .QN(n3535) );
  DFFX1_LVT u_T_427_reg_0__8_ ( .D(n4340), .CLK(n4279), .Q(n_T_427[1889]), 
        .QN(n3534) );
  DFFX1_LVT u_T_427_reg_0__7_ ( .D(n4337), .CLK(n4279), .Q(n_T_427[1888]), 
        .QN(n3533) );
  DFFX1_LVT u_T_427_reg_0__6_ ( .D(n4334), .CLK(n4279), .Q(n_T_427[1887]), 
        .QN(n3532) );
  DFFX1_LVT u_T_427_reg_0__3_ ( .D(n4325), .CLK(n4279), .QN(n3531) );
  DFFX1_LVT u_T_427_reg_0__1_ ( .D(n4319), .CLK(n4279), .Q(n_T_427[1883]), 
        .QN(n3530) );
  DFFX1_LVT u_T_427_reg_4__59_ ( .D(n4482), .CLK(n4259), .Q(n_T_427[1722]), 
        .QN(n3518) );
  DFFX1_LVT u_T_427_reg_3__59_ ( .D(n4482), .CLK(n4265), .Q(n_T_427[1786]), 
        .QN(n3517) );
  DFFX1_LVT u_T_427_reg_3__57_ ( .D(n4476), .CLK(n4265), .Q(n_T_427[1784]), 
        .QN(n3515) );
  DFFX1_LVT u_T_427_reg_4__55_ ( .D(n4470), .CLK(n4259), .Q(n_T_427[1718]), 
        .QN(n3513) );
  DFFX1_LVT u_T_427_reg_3__55_ ( .D(n4470), .CLK(n4265), .Q(n_T_427[1782]), 
        .QN(n3512) );
  DFFX1_LVT u_T_427_reg_3__53_ ( .D(n4464), .CLK(n4265), .Q(n_T_427[1780]), 
        .QN(n3510) );
  DFFX1_LVT u_T_427_reg_3__50_ ( .D(n4455), .CLK(n4265), .Q(n_T_427[1777]), 
        .QN(n3507) );
  DFFX1_LVT u_T_427_reg_3__48_ ( .D(n4449), .CLK(n4265), .Q(n_T_427[1775]), 
        .QN(n3505) );
  DFFX1_LVT u_T_427_reg_3__47_ ( .D(n4446), .CLK(n4264), .Q(n_T_427[1774]), 
        .QN(n3504) );
  DFFX1_LVT u_T_427_reg_3__40_ ( .D(n4425), .CLK(n4264), .Q(n_T_427[1767]), 
        .QN(n3499) );
  DFFX1_LVT u_T_427_reg_3__37_ ( .D(n4417), .CLK(n4264), .Q(n_T_427[1764]), 
        .QN(n3498) );
  DFFX1_LVT u_T_427_reg_4__32_ ( .D(n4404), .CLK(n4257), .Q(n_T_427[1695]), 
        .QN(n3496) );
  DFFX1_LVT u_T_427_reg_3__32_ ( .D(n4404), .CLK(n4263), .Q(n_T_427[1759]), 
        .QN(n3495) );
  DFFX1_LVT u_T_427_reg_4__17_ ( .D(n4365), .CLK(n4256), .Q(n_T_427[1680]), 
        .QN(n3494) );
  DFFX1_LVT u_T_427_reg_0__59_ ( .D(n4482), .CLK(n4283), .Q(n_T_427[1938]), 
        .QN(n3493) );
  DFFX1_LVT u_T_427_reg_0__57_ ( .D(n4476), .CLK(n4283), .Q(n_T_427[1936]), 
        .QN(n3491) );
  DFFX1_LVT u_T_427_reg_20__47_ ( .D(n4447), .CLK(n4162), .Q(n_T_427[687]), 
        .QN(n3482) );
  DFFX1_LVT u_T_427_reg_1__38_ ( .D(n4420), .CLK(n4276), .Q(n_T_427[1877]), 
        .QN(n3481) );
  DFFX1_LVT u_T_427_reg_1__35_ ( .D(n4412), .CLK(n4275), .Q(n_T_427[1876]), 
        .QN(n3480) );
  DFFX1_LVT u_T_427_reg_1__33_ ( .D(n4407), .CLK(n4275), .Q(n_T_427[1874]), 
        .QN(n3479) );
  DFFX1_LVT u_T_427_reg_1__31_ ( .D(n4402), .CLK(n4275), .Q(n_T_427[1873]), 
        .QN(n3376) );
  DFFX1_LVT u_T_427_reg_1__28_ ( .D(n4394), .CLK(n4275), .Q(n_T_427[1871]), 
        .QN(n3374) );
  DFFX1_LVT u_T_427_reg_1__26_ ( .D(n4389), .CLK(n4275), .Q(n_T_427[1869]), 
        .QN(n3373) );
  DFFX1_LVT u_T_427_reg_1__25_ ( .D(n4387), .CLK(n4275), .Q(n_T_427[1868]), 
        .QN(n3372) );
  DFFX1_LVT u_T_427_reg_1__22_ ( .D(n4379), .CLK(n4274), .QN(n3371) );
  DFFX1_LVT u_T_427_reg_1__21_ ( .D(n4377), .CLK(n4274), .Q(n_T_427[1866]), 
        .QN(n3370) );
  DFFX1_LVT u_T_427_reg_4__38_ ( .D(n4420), .CLK(n4258), .Q(n_T_427[1701]), 
        .QN(n3685) );
  DFFX1_LVT u_T_427_reg_4__33_ ( .D(n4407), .CLK(n4257), .Q(n_T_427[1696]), 
        .QN(n3655) );
  DFFX1_LVT u_T_427_reg_2__47_ ( .D(n4446), .CLK(n4270), .Q(n_T_427[1835]), 
        .QN(n3477) );
  DFFX1_LVT u_T_427_reg_2__50_ ( .D(n4455), .CLK(n4271), .Q(n_T_427[1838]), 
        .QN(n3476) );
  DFFX1_LVT u_T_427_reg_2__57_ ( .D(n4476), .CLK(n4271), .Q(n_T_427[1844]), 
        .QN(n3473) );
  DFFX1_LVT u_T_427_reg_2__53_ ( .D(n4464), .CLK(n4271), .Q(n_T_427[1841]), 
        .QN(n3470) );
  DFFX1_LVT u_T_427_reg_2__46_ ( .D(n4443), .CLK(n4270), .Q(n_T_427[1834]), 
        .QN(n3467) );
  DFFX1_LVT u_T_427_reg_1__46_ ( .D(n4443), .CLK(n4276), .Q(n_T_427[1880]), 
        .QN(n3466) );
  DFFX1_LVT u_T_427_reg_1__44_ ( .D(n4437), .CLK(n4276), .Q(n_T_427[1879]), 
        .QN(n3465) );
  DFFX1_LVT u_T_427_reg_19__40_ ( .D(n4426), .CLK(n4168), .Q(n_T_427[743]), 
        .QN(n3461) );
  DFFX1_LVT u_T_427_reg_2__40_ ( .D(n4425), .CLK(n4270), .Q(n_T_427[1828]), 
        .QN(n3460) );
  DFFX1_LVT u_T_427_reg_7__39_ ( .D(n4422), .CLK(n4240), .Q(n_T_427[1510]), 
        .QN(n3459) );
  DFFX1_LVT u_T_427_reg_2__39_ ( .D(n4422), .CLK(n4270), .Q(n_T_427[1827]), 
        .QN(n3458) );
  DFFX1_LVT u_T_427_reg_1__39_ ( .D(n4422), .CLK(n4276), .Q(n_T_427[1878]), 
        .QN(n3457) );
  DFFX1_LVT u_T_427_reg_2__37_ ( .D(n4417), .CLK(n4270), .Q(n_T_427[1825]), 
        .QN(n3456) );
  DFFX1_LVT u_T_427_reg_2__34_ ( .D(n4409), .CLK(n4269), .Q(n_T_427[1822]), 
        .QN(n3453) );
  DFFX1_LVT u_T_427_reg_1__34_ ( .D(n4409), .CLK(n4275), .Q(n_T_427[1875]), 
        .QN(n3452) );
  DFFX1_LVT u_T_427_reg_2__23_ ( .D(n4381), .CLK(n4268), .Q(n_T_427[1812]), 
        .QN(n3448) );
  DFFX1_LVT u_T_427_reg_2__16_ ( .D(n4362), .CLK(n4268), .Q(n_T_427[1806]), 
        .QN(n3444) );
  DFFX1_LVT u_T_427_reg_12__15_ ( .D(n4360), .CLK(n4208), .Q(n_T_427[1166]), 
        .QN(n3443) );
  DFFX1_LVT u_T_427_reg_7__15_ ( .D(n4360), .CLK(n4238), .Q(n_T_427[1486]), 
        .QN(n3442) );
  DFFX1_LVT u_T_427_reg_12__14_ ( .D(n4358), .CLK(n4208), .Q(n_T_427[1165]), 
        .QN(n3441) );
  DFFX1_LVT u_T_427_reg_7__14_ ( .D(n4357), .CLK(n4238), .Q(n_T_427[1485]), 
        .QN(n3440) );
  DFFX1_LVT u_T_427_reg_12__13_ ( .D(n4355), .CLK(n4208), .Q(n_T_427[1164]), 
        .QN(n3439) );
  DFFX1_LVT u_T_427_reg_7__13_ ( .D(n4355), .CLK(n4238), .Q(n_T_427[1484]), 
        .QN(n3438) );
  DFFX1_LVT u_T_427_reg_12__12_ ( .D(n4353), .CLK(n4208), .Q(n_T_427[1163]), 
        .QN(n3437) );
  DFFX1_LVT u_T_427_reg_7__12_ ( .D(n4352), .CLK(n4238), .Q(n_T_427[1483]), 
        .QN(n3436) );
  DFFX1_LVT u_T_427_reg_12__10_ ( .D(n4347), .CLK(n4207), .Q(n_T_427[1161]), 
        .QN(n3434) );
  DFFX1_LVT u_T_427_reg_7__10_ ( .D(n4346), .CLK(n4237), .Q(n_T_427[1481]), 
        .QN(n3433) );
  DFFX1_LVT u_T_427_reg_12__9_ ( .D(n4344), .CLK(n4207), .Q(n_T_427[1160]), 
        .QN(n3432) );
  DFFX1_LVT u_T_427_reg_7__9_ ( .D(n4343), .CLK(n4237), .Q(n_T_427[1480]), 
        .QN(n3431) );
  DFFX1_LVT u_T_427_reg_12__8_ ( .D(n4341), .CLK(n4207), .Q(n_T_427[1159]), 
        .QN(n3430) );
  DFFX1_LVT u_T_427_reg_7__8_ ( .D(n4340), .CLK(n4237), .Q(n_T_427[1479]), 
        .QN(n3429) );
  DFFX1_LVT u_T_427_reg_12__7_ ( .D(n4338), .CLK(n4207), .Q(n_T_427[1158]), 
        .QN(n3428) );
  DFFX1_LVT u_T_427_reg_7__7_ ( .D(n4337), .CLK(n4237), .Q(n_T_427[1478]), 
        .QN(n3427) );
  DFFX1_LVT u_T_427_reg_12__6_ ( .D(n4335), .CLK(n4207), .Q(n_T_427[1157]), 
        .QN(n3426) );
  DFFX1_LVT u_T_427_reg_7__6_ ( .D(n4334), .CLK(n4237), .Q(n_T_427[1477]), 
        .QN(n3425) );
  DFFX1_LVT u_T_427_reg_12__5_ ( .D(n4332), .CLK(n4207), .Q(n_T_427[1156]), 
        .QN(n3424) );
  DFFX1_LVT u_T_427_reg_7__5_ ( .D(n4331), .CLK(n4237), .Q(n_T_427[1476]), 
        .QN(n3423) );
  DFFX1_LVT u_T_427_reg_12__4_ ( .D(n4329), .CLK(n4207), .Q(n_T_427[1155]) );
  DFFX1_LVT u_T_427_reg_7__4_ ( .D(n4328), .CLK(n4237), .Q(n_T_427[1475]), 
        .QN(n3422) );
  DFFX1_LVT u_T_427_reg_12__3_ ( .D(n4326), .CLK(n4207), .Q(n_T_427[1154]), 
        .QN(n3421) );
  DFFX1_LVT u_T_427_reg_7__3_ ( .D(n4325), .CLK(n4237), .Q(n_T_427[1474]), 
        .QN(n3420) );
  DFFX1_LVT u_T_427_reg_12__2_ ( .D(n4323), .CLK(n4207), .Q(n_T_427[1153]), 
        .QN(n3419) );
  DFFX1_LVT u_T_427_reg_7__2_ ( .D(n4322), .CLK(n4237), .Q(n_T_427[1473]), 
        .QN(n3418) );
  DFFX1_LVT u_T_427_reg_2__44_ ( .D(n4437), .CLK(n4270), .Q(n_T_427[1832]), 
        .QN(n3415) );
  DFFX1_LVT u_T_427_reg_2__48_ ( .D(n4449), .CLK(n4271), .Q(n_T_427[1836]), 
        .QN(n3414) );
  DFFX1_LVT u_T_427_reg_14__59_ ( .D(n4483), .CLK(n4199), .Q(n_T_427[1082]), 
        .QN(n3368) );
  DFFX1_LVT u_T_427_reg_12__59_ ( .D(n4483), .CLK(n4211), .Q(n_T_427[1210]), 
        .QN(n3367) );
  DFFX1_LVT u_T_427_reg_14__57_ ( .D(n4477), .CLK(n4199), .Q(n_T_427[1080]), 
        .QN(n3364) );
  DFFX1_LVT u_T_427_reg_12__57_ ( .D(n4477), .CLK(n4211), .Q(n_T_427[1208]), 
        .QN(n3363) );
  DFFX1_LVT u_T_427_reg_12__55_ ( .D(n4471), .CLK(n4211), .Q(n_T_427[1206]), 
        .QN(n3361) );
  DFFX1_LVT u_T_427_reg_12__53_ ( .D(n4465), .CLK(n4211), .Q(n_T_427[1204]), 
        .QN(n3358) );
  DFFX1_LVT u_T_427_reg_14__53_ ( .D(n4465), .CLK(n4199), .Q(n_T_427[1076]), 
        .QN(n3357) );
  DFFX1_LVT u_T_427_reg_12__50_ ( .D(n4456), .CLK(n4211), .Q(n_T_427[1201]), 
        .QN(n3352) );
  DFFX1_LVT u_T_427_reg_14__50_ ( .D(n4456), .CLK(n4199), .Q(n_T_427[1073]), 
        .QN(n3351) );
  DFFX1_LVT u_T_427_reg_12__48_ ( .D(n4450), .CLK(n4211), .Q(n_T_427[1199]), 
        .QN(n3348) );
  DFFX1_LVT u_T_427_reg_14__47_ ( .D(n4447), .CLK(n4198), .Q(n_T_427[1070]), 
        .QN(n3347) );
  DFFX1_LVT u_T_427_reg_12__47_ ( .D(n4447), .CLK(n4210), .Q(n_T_427[1198]), 
        .QN(n3346) );
  DFFX1_LVT u_T_427_reg_12__46_ ( .D(n4444), .CLK(n4210), .Q(n_T_427[1197]), 
        .QN(n3345) );
  DFFX1_LVT u_T_427_reg_12__44_ ( .D(n4438), .CLK(n4210), .Q(n_T_427[1195]), 
        .QN(n3342) );
  DFFX1_LVT u_T_427_reg_14__40_ ( .D(n4426), .CLK(n4198), .Q(n_T_427[1063]), 
        .QN(n3338) );
  DFFX1_LVT u_T_427_reg_12__40_ ( .D(n4426), .CLK(n4210), .Q(n_T_427[1191]), 
        .QN(n3337) );
  DFFX1_LVT u_T_427_reg_12__37_ ( .D(n4418), .CLK(n4210), .Q(n_T_427[1188]), 
        .QN(n3336) );
  DFFX1_LVT u_T_427_reg_12__34_ ( .D(n4410), .CLK(n4209), .Q(n_T_427[1185]), 
        .QN(n3335) );
  DFFX1_LVT u_T_427_reg_12__32_ ( .D(n4405), .CLK(n4209), .Q(n_T_427[1183]), 
        .QN(n3334) );
  DFFX1_LVT u_T_427_reg_14__32_ ( .D(n4405), .CLK(n4197), .Q(n_T_427[1055]), 
        .QN(n3333) );
  DFFX1_LVT u_T_427_reg_1__23_ ( .D(n4381), .CLK(n4274), .Q(n_T_427[1867]), 
        .QN(n3325) );
  DFFX1_LVT u_T_427_reg_14__23_ ( .D(n4382), .CLK(n4196), .Q(n_T_427[1046]), 
        .QN(n3324) );
  DFFX1_LVT u_T_427_reg_12__23_ ( .D(n4382), .CLK(n4208), .Q(n_T_427[1174]), 
        .QN(n3323) );
  DFFX1_LVT u_T_427_reg_12__17_ ( .D(n4366), .CLK(n4208), .Q(n_T_427[1168]), 
        .QN(n3313) );
  DFFX1_LVT u_T_427_reg_12__16_ ( .D(n4363), .CLK(n4208), .Q(n_T_427[1167]), 
        .QN(n3312) );
  DFFX1_LVT u_T_427_reg_20__39_ ( .D(n4423), .CLK(n4162), .Q(n_T_427[679]), 
        .QN(n3179) );
  DFFX1_LVT u_T_427_reg_0__16_ ( .D(n4362), .CLK(n4280), .Q(n_T_427[1897]), 
        .QN(n3524) );
  DFFX1_LVT u_T_427_reg_19__50_ ( .D(n4456), .CLK(n4169), .Q(n_T_427[753]), 
        .QN(n3407) );
  DFFX1_LVT u_T_427_reg_19__46_ ( .D(n4444), .CLK(n4168), .Q(n_T_427[749]), 
        .QN(n3406) );
  DFFX1_LVT u_T_427_reg_7__38_ ( .D(n4420), .CLK(n4240), .Q(n_T_427[1509]), 
        .QN(n3403) );
  DFFX1_LVT u_T_427_reg_2__38_ ( .D(n4420), .CLK(n4270), .Q(n_T_427[1826]), 
        .QN(n3402) );
  DFFX1_LVT u_T_427_reg_2__35_ ( .D(n4412), .CLK(n4269), .Q(n_T_427[1823]), 
        .QN(n3401) );
  DFFX1_LVT u_T_427_reg_19__35_ ( .D(n4412), .CLK(n4167), .Q(n_T_427[738]), 
        .QN(n3400) );
  DFFX1_LVT u_T_427_reg_2__33_ ( .D(n4407), .CLK(n4269), .Q(n_T_427[1821]), 
        .QN(n3399) );
  DFFX1_LVT u_T_427_reg_19__32_ ( .D(n4405), .CLK(n4167), .Q(n_T_427[736]), 
        .QN(n3398) );
  DFFX1_LVT u_T_427_reg_2__31_ ( .D(n4402), .CLK(n4269), .Q(n_T_427[1820]), 
        .QN(n3397) );
  DFFX1_LVT u_T_427_reg_2__28_ ( .D(n4394), .CLK(n4269), .Q(n_T_427[1817]), 
        .QN(n3395) );
  DFFX1_LVT u_T_427_reg_2__26_ ( .D(n4389), .CLK(n4269), .Q(n_T_427[1815]), 
        .QN(n3394) );
  DFFX1_LVT u_T_427_reg_2__25_ ( .D(n4387), .CLK(n4269), .Q(n_T_427[1814]), 
        .QN(n3393) );
  DFFX1_LVT u_T_427_reg_2__22_ ( .D(n4379), .CLK(n4268), .Q(n_T_427[1811]), 
        .QN(n3392) );
  DFFX1_LVT u_T_427_reg_2__21_ ( .D(n4377), .CLK(n4268), .Q(n_T_427[1810]), 
        .QN(n3391) );
  DFFX1_LVT u_T_427_reg_4__15_ ( .D(n4360), .CLK(n4256), .Q(n_T_427[1678]), 
        .QN(n3390) );
  DFFX1_LVT u_T_427_reg_4__14_ ( .D(n4357), .CLK(n4256), .Q(n_T_427[1677]), 
        .QN(n3389) );
  DFFX1_LVT u_T_427_reg_4__13_ ( .D(n4355), .CLK(n4256), .Q(n_T_427[1676]), 
        .QN(n3388) );
  DFFX1_LVT u_T_427_reg_4__12_ ( .D(n4352), .CLK(n4256), .Q(n_T_427[1675]), 
        .QN(n3387) );
  DFFX1_LVT u_T_427_reg_12__11_ ( .D(n4350), .CLK(n4207), .Q(n_T_427[1162]) );
  DFFX1_LVT u_T_427_reg_7__11_ ( .D(n4350), .CLK(n4237), .Q(n_T_427[1482]), 
        .QN(n3386) );
  DFFX1_LVT u_T_427_reg_4__10_ ( .D(n4346), .CLK(n4255), .Q(n_T_427[1673]), 
        .QN(n3385) );
  DFFX1_LVT u_T_427_reg_4__9_ ( .D(n4343), .CLK(n4255), .Q(n_T_427[1672]), 
        .QN(n3384) );
  DFFX1_LVT u_T_427_reg_4__8_ ( .D(n4340), .CLK(n4255), .Q(n_T_427[1671]), 
        .QN(n3383) );
  DFFX1_LVT u_T_427_reg_4__7_ ( .D(n4337), .CLK(n4255), .Q(n_T_427[1670]), 
        .QN(n3382) );
  DFFX1_LVT u_T_427_reg_4__6_ ( .D(n4334), .CLK(n4255), .Q(n_T_427[1669]), 
        .QN(n3381) );
  DFFX1_LVT u_T_427_reg_4__5_ ( .D(n4331), .CLK(n4255), .Q(n_T_427[1668]), 
        .QN(n3380) );
  DFFX1_LVT u_T_427_reg_4__4_ ( .D(n4328), .CLK(n4255), .Q(n_T_427[1667]), 
        .QN(n3379) );
  DFFX1_LVT u_T_427_reg_4__3_ ( .D(n4325), .CLK(n4255), .Q(n_T_427[1666]), 
        .QN(n3378) );
  DFFX1_LVT u_T_427_reg_4__2_ ( .D(n4322), .CLK(n4255), .Q(n_T_427[1665]), 
        .QN(n3377) );
  DFFX1_LVT u_T_427_reg_19__57_ ( .D(n4477), .CLK(n4169), .Q(n_T_427[760]), 
        .QN(n3302) );
  DFFX1_LVT u_T_427_reg_19__55_ ( .D(n4471), .CLK(n4169), .Q(n_T_427[758]), 
        .QN(n3301) );
  DFFX1_LVT u_T_427_reg_14__46_ ( .D(n4444), .CLK(n4198), .Q(n_T_427[1069]), 
        .QN(n3300) );
  DFFX1_LVT u_T_427_reg_12__35_ ( .D(n4412), .CLK(n4209), .Q(n_T_427[1186]), 
        .QN(n3299) );
  DFFX1_LVT u_T_427_reg_12__33_ ( .D(n4407), .CLK(n4209), .Q(n_T_427[1184]), 
        .QN(n3298) );
  DFFX1_LVT u_T_427_reg_14__31_ ( .D(n4402), .CLK(n4197), .Q(n_T_427[1054]), 
        .QN(n3297) );
  DFFX1_LVT u_T_427_reg_12__31_ ( .D(n4402), .CLK(n4209), .Q(n_T_427[1182]), 
        .QN(n3296) );
  DFFX1_LVT u_T_427_reg_14__28_ ( .D(n4394), .CLK(n4197), .Q(n_T_427[1051]), 
        .QN(n3293) );
  DFFX1_LVT u_T_427_reg_12__28_ ( .D(n4394), .CLK(n4209), .Q(n_T_427[1179]), 
        .QN(n3292) );
  DFFX1_LVT u_T_427_reg_14__26_ ( .D(n4389), .CLK(n4197), .Q(n_T_427[1049]), 
        .QN(n3291) );
  DFFX1_LVT u_T_427_reg_12__26_ ( .D(n4389), .CLK(n4209), .Q(n_T_427[1177]), 
        .QN(n3290) );
  DFFX1_LVT u_T_427_reg_14__25_ ( .D(n4387), .CLK(n4197), .Q(n_T_427[1048]), 
        .QN(n3289) );
  DFFX1_LVT u_T_427_reg_12__25_ ( .D(n4387), .CLK(n4209), .Q(n_T_427[1176]), 
        .QN(n3288) );
  DFFX1_LVT u_T_427_reg_14__22_ ( .D(n4379), .CLK(n4196), .Q(n_T_427[1045]), 
        .QN(n3287) );
  DFFX1_LVT u_T_427_reg_12__22_ ( .D(n4379), .CLK(n4208), .Q(n_T_427[1173]), 
        .QN(n3286) );
  DFFX1_LVT u_T_427_reg_14__21_ ( .D(n4377), .CLK(n4196), .Q(n_T_427[1044]), 
        .QN(n3285) );
  DFFX1_LVT u_T_427_reg_12__21_ ( .D(n4377), .CLK(n4208), .Q(n_T_427[1172]), 
        .QN(n3284) );
  DFFX1_LVT u_T_427_reg_14__17_ ( .D(n4366), .CLK(n4196), .Q(n_T_427[1040]), 
        .QN(n3283) );
  DFFX1_LVT u_T_427_reg_14__16_ ( .D(n4363), .CLK(n4196), .Q(n_T_427[1039]), 
        .QN(n3282) );
  DFFX1_LVT u_T_427_reg_20__35_ ( .D(n4413), .CLK(n4161), .Q(n_T_427[675]), 
        .QN(n3369) );
  DFFX1_LVT u_T_427_reg_20__4_ ( .D(n4329), .CLK(n4159), .Q(n_T_427[644]), 
        .QN(n3174) );
  DFFX1_LVT u_T_427_reg_20__2_ ( .D(n4323), .CLK(n4159), .Q(n_T_427[642]), 
        .QN(n3173) );
  DFFX2_LVT ex_ctrl_alu_fn_reg_2_ ( .D(N283), .CLK(n4313), .Q(alu_io_fn[2]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_50_ ( .D(N732), .CLK(net34650), .Q(n_T_628[52]) );
  DFFX1_LVT mem_reg_sfence_reg ( .D(n2525), .CLK(clock), .Q(n326), .QN(
        mem_reg_sfence) );
  DFFX1_LVT u_T_1057_reg ( .D(n2524), .CLK(n4499), .Q(n_T_1057) );
  DFFASX1_LVT imem_might_request_reg_reg ( .D(N271), .CLK(clock), .SETB(1'b1), 
        .Q(io_imem_might_request) );
  DFFASX1_LVT wb_reg_inst_reg_8_ ( .D(n_T_849[1]), .CLK(n4311), .SETB(1'b1), 
        .Q(wb_waddr[1]), .QN(n3103) );
  OA21X1_LVT wb_reg_cause_reg_63__U2 ( .A1(mem_reg_xcpt_interrupt), .A2(
        mem_reg_xcpt), .A3(mem_reg_cause[63]), .Y(n2521) );
  DFFASX1_LVT wb_reg_cause_reg_63_ ( .D(n2521), .CLK(n4311), .SETB(1'b1), .Q(
        wb_reg_cause[63]) );
  DFFASX1_LVT mem_reg_cause_reg_63_ ( .D(n308), .CLK(net34480), .SETB(1'b1), 
        .QN(mem_reg_cause[63]) );
  OA21X1_LVT wb_reg_cause_reg_1__U2 ( .A1(n5168), .A2(n63), .A3(n1281), .Y(
        n2518) );
  DFFASX1_LVT wb_reg_cause_reg_1_ ( .D(n2518), .CLK(n4300), .SETB(1'b1), .QN(
        wb_reg_cause[1]) );
  INVX0_LVT mem_reg_slow_bypass_reg_U4 ( .A(io_dmem_req_bits_size[1]), .Y(
        n2515) );
  DFFX1_LVT mem_reg_slow_bypass_reg ( .D(n2516), .CLK(n4285), .Q(
        mem_reg_slow_bypass) );
  OA21X1_LVT mem_reg_flush_pipe_reg_U2 ( .A1(n2495), .A2(n9516), .A3(n309), 
        .Y(n2514) );
  DFFX1_LVT mem_reg_flush_pipe_reg ( .D(n2514), .CLK(n4285), .Q(n64), .QN(
        mem_reg_flush_pipe) );
  DFFSSRX1_LVT ex_reg_rvc_reg ( .D(n9430), .SETB(1'b1), .RSTB(n4497), .CLK(
        net34469), .Q(n3215), .QN(ex_reg_rvc) );
  DFFSSRX1_LVT ex_ctrl_fp_reg ( .D(1'b0), .SETB(1'b0), .RSTB(n2512), .CLK(
        n4312), .Q(n322), .QN(io_dmem_req_bits_tag[0]) );
  DFFSSRX1_LVT ex_ctrl_mem_reg ( .D(1'b0), .SETB(1'b0), .RSTB(n2510), .CLK(
        n4312), .Q(n312), .QN(ex_ctrl_mem) );
  DFFX1_LVT ex_reg_cause_reg_63_ ( .D(csr_io_interrupt), .CLK(net34640), .QN(
        n308) );
  DFFSSRX1_LVT wb_reg_valid_reg ( .D(io_dmem_s1_kill), .SETB(n9425), .RSTB(
        1'b1), .CLK(n4499), .Q(n3203), .QN(wb_reg_valid) );
  DFFSSRX1_LVT ex_ctrl_mem_cmd_reg_1_ ( .D(n9520), .SETB(n9435), .RSTB(n1853), 
        .CLK(net34469), .Q(io_dmem_req_bits_cmd[1]), .QN(n559) );
  DFFASX1_LVT ex_reg_cause_reg_3_ ( .D(n2507), .CLK(net34640), .SETB(1'b1), 
        .Q(n75) );
  DFFSSRX1_LVT u_T_1185_reg_27_ ( .D(n5310), .SETB(1'b1), .RSTB(n5309), .CLK(
        net34660), .Q(n3135), .QN(n_T_1187[27]) );
  DFFSSRX1_LVT wb_reg_flush_pipe_reg ( .D(n64), .SETB(n1829), .RSTB(1'b1), 
        .CLK(clock), .QN(wb_reg_flush_pipe) );
  DFFSSRX1_LVT ex_reg_rs_bypass_0_reg ( .D(n9412), .SETB(1'b1), .RSTB(n1262), 
        .CLK(net34469), .Q(n3101), .QN(n2493) );
  DFFSSRX1_LVT ex_ctrl_mem_cmd_reg_3_ ( .D(1'b0), .SETB(n3578), .RSTB(n5138), 
        .CLK(net34469), .Q(io_dmem_req_bits_cmd[3]), .QN(n3122) );
  DFFSSRX1_LVT ex_ctrl_sel_alu1_reg_1_ ( .D(1'b0), .SETB(n2675), .RSTB(n9100), 
        .CLK(net34469), .Q(n561) );
  DFFSSRX1_LVT mem_reg_xcpt_reg ( .D(n2501), .SETB(n98), .RSTB(n407), .CLK(
        clock), .Q(mem_reg_xcpt), .QN(n3251) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_38_ ( .D(N720), .CLK(n4083), .Q(n_T_628[40])
         );
  DFFSSRX1_LVT ex_reg_xcpt_reg ( .D(n2874), .SETB(n1431), .RSTB(1'b1), .CLK(
        n4499), .QN(n2501) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_59_ ( .D(N741), .CLK(n4084), .Q(n_T_628[61])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_32_ ( .D(N714), .CLK(n4082), .Q(n_T_628[34])
         );
  AO221X1_LVT U2645 ( .A1(1'b1), .A2(n2234), .A3(n9158), .A4(n_T_642[3]), .A5(
        n2236), .Y(alu_io_in2[3]) );
  OA221X1_LVT U2646 ( .A1(1'b0), .A2(n1628), .A3(n9090), .A4(n2238), .A5(n2239), .Y(n2241) );
  OA221X1_LVT U2647 ( .A1(1'b0), .A2(n2199), .A3(n9512), .A4(n_T_698[1]), .A5(
        n2200), .Y(n2202) );
  OA221X1_LVT U2648 ( .A1(1'b0), .A2(n2208), .A3(n_T_698[13]), .A4(n9500), 
        .A5(n2209), .Y(n2210) );
  OA221X1_LVT U2649 ( .A1(1'b0), .A2(n2196), .A3(n9488), .A4(n_T_698[23]), 
        .A5(n2210), .Y(n2211) );
  OA21X1_LVT U2650 ( .A1(n3195), .A2(n3596), .A3(n2035), .Y(n2337) );
  IBUFFX2_LVT U2651 ( .A(n9517), .Y(n9434) );
  NAND3X4_LVT U2652 ( .A1(n3078), .A2(n9519), .A3(n9434), .Y(n5072) );
  AND2X1_LVT U2653 ( .A1(n3573), .A2(n3572), .Y(n1832) );
  AND2X1_LVT U2654 ( .A1(n6914), .A2(n1832), .Y(n6965) );
  AND2X1_LVT U2655 ( .A1(n6906), .A2(n1832), .Y(n5124) );
  AND4X1_LVT U2656 ( .A1(n2623), .A2(n2624), .A3(n5161), .A4(n5162), .Y(n2170)
         );
  NAND3X0_LVT U2657 ( .A1(n5147), .A2(n5173), .A3(n1833), .Y(n5162) );
  NAND3X0_LVT U2658 ( .A1(n5145), .A2(n3079), .A3(n1834), .Y(n1833) );
  AO21X1_LVT U2659 ( .A1(n2528), .A2(n9434), .A3(n5143), .Y(n1834) );
  NAND2X0_LVT U2660 ( .A1(n2138), .A2(n1835), .Y(n5174) );
  INVX1_LVT U2661 ( .A(io_fpu_inst[28]), .Y(n1835) );
  NOR2X0_LVT U2662 ( .A1(n3783), .A2(n2139), .Y(n2138) );
  NAND3X0_LVT U2663 ( .A1(n5107), .A2(n1837), .A3(n5106), .Y(n5108) );
  OR2X1_LVT U2664 ( .A1(n1836), .A2(n1431), .Y(n9229) );
  OR2X1_LVT U2665 ( .A1(n1837), .A2(n9092), .Y(n1836) );
  AND2X1_LVT U2666 ( .A1(io_fpu_inst[5]), .A2(n9522), .Y(n1837) );
  NAND2X0_LVT U2667 ( .A1(n1838), .A2(n5173), .Y(n5135) );
  INVX1_LVT U2668 ( .A(io_fpu_inst[13]), .Y(n1838) );
  OA22X1_LVT U2669 ( .A1(n9079), .A2(n1839), .A3(n3079), .A4(n5133), .Y(n2642)
         );
  INVX1_LVT U2670 ( .A(n5173), .Y(n1839) );
  AND2X1_LVT U2671 ( .A1(n9105), .A2(n3593), .Y(n5173) );
  OA21X1_LVT U2672 ( .A1(n4504), .A2(n1840), .A3(n4506), .Y(n4512) );
  OR3X1_LVT U2673 ( .A1(n2553), .A2(n5099), .A3(n4509), .Y(n1840) );
  AOI22X1_LVT U2674 ( .A1(n2648), .A2(n2649), .A3(n5173), .A4(n2647), .Y(n2658) );
  NAND4X0_LVT U2675 ( .A1(n3723), .A2(n3724), .A3(n8914), .A4(n1841), .Y(n8924) );
  AND2X1_LVT U2676 ( .A1(n8913), .A2(n8912), .Y(n1841) );
  AND3X1_LVT U2677 ( .A1(n3590), .A2(io_fpu_inst[6]), .A3(n9529), .Y(n2649) );
  INVX0_LVT U2678 ( .A(n9113), .Y(n3582) );
  AND3X1_LVT U2679 ( .A1(n5075), .A2(io_fpu_inst[5]), .A3(n3597), .Y(n5119) );
  IBUFFX2_LVT U2680 ( .A(n3708), .Y(n3771) );
  NAND2X1_LVT U2681 ( .A1(n3771), .A2(n_T_427[763]), .Y(n8910) );
  NAND3X1_LVT U2682 ( .A1(n7105), .A2(n7104), .A3(n7103), .Y(n7106) );
  NAND3X0_LVT U2683 ( .A1(n2166), .A2(n8125), .A3(n1842), .Y(N718) );
  AND3X1_LVT U2684 ( .A1(n2165), .A2(n8126), .A3(n8124), .Y(n1842) );
  NAND3X1_LVT U2685 ( .A1(n7087), .A2(n7086), .A3(n7085), .Y(n7109) );
  AND2X1_LVT U2686 ( .A1(n2552), .A2(n3590), .Y(n5074) );
  AOI22X2_LVT U2687 ( .A1(n1844), .A2(n1843), .A3(n_T_427[1016]), .A4(n3755), 
        .Y(n1855) );
  IBUFFX2_LVT U2688 ( .A(n3364), .Y(n1843) );
  IBUFFX2_LVT U2689 ( .A(n4013), .Y(n1844) );
  NAND2X1_LVT U2690 ( .A1(n2882), .A2(n_T_427[1916]), .Y(n8046) );
  NAND3X1_LVT U2691 ( .A1(n7083), .A2(n7082), .A3(n7081), .Y(n7110) );
  NAND2X4_LVT U2692 ( .A1(n9105), .A2(n3593), .Y(n3039) );
  NAND4X1_LVT U2693 ( .A1(n8312), .A2(n8310), .A3(n8311), .A4(n2608), .Y(n8313) );
  NOR2X0_LVT U2694 ( .A1(n8314), .A2(n8313), .Y(n3035) );
  NAND3X0_LVT U2695 ( .A1(n8051), .A2(n8049), .A3(n8050), .Y(n8080) );
  OA21X1_LVT U2696 ( .A1(n2657), .A2(n2637), .A3(n2633), .Y(n5110) );
  NAND2X0_LVT U2697 ( .A1(n2169), .A2(n2170), .Y(n2144) );
  NAND4X0_LVT U2698 ( .A1(n2894), .A2(n1892), .A3(n2893), .A4(n1845), .Y(N689)
         );
  AND3X1_LVT U2699 ( .A1(n2937), .A2(n1900), .A3(n1846), .Y(n1845) );
  AND2X1_LVT U2700 ( .A1(n7245), .A2(n7244), .Y(n1846) );
  NAND2X0_LVT U2701 ( .A1(n_T_427[1650]), .A2(n3652), .Y(n8596) );
  AND2X1_LVT U2702 ( .A1(n2933), .A2(n2934), .Y(n1888) );
  NAND2X0_LVT U2703 ( .A1(n_T_427[1662]), .A2(n3643), .Y(n9023) );
  NBUFFX2_LVT U2704 ( .A(n5116), .Y(n1847) );
  NAND2X0_LVT U2705 ( .A1(n_T_427[810]), .A2(n9056), .Y(n8323) );
  NAND2X0_LVT U2706 ( .A1(n_T_427[826]), .A2(n9056), .Y(n8884) );
  IBUFFX32_LVT U2707 ( .A(n3137), .Y(n1848) );
  NAND2X0_LVT U2708 ( .A1(n1848), .A2(n3692), .Y(n3569) );
  NAND2X0_LVT U2709 ( .A1(n_T_427[1400]), .A2(n3610), .Y(n8781) );
  IBUFFX2_LVT U2710 ( .A(n9095), .Y(n2570) );
  NAND3X4_LVT U2711 ( .A1(n5101), .A2(n2570), .A3(n9097), .Y(n5104) );
  AND2X1_LVT U2712 ( .A1(n2561), .A2(n3765), .Y(n3772) );
  AND3X1_LVT U2713 ( .A1(n4511), .A2(n4513), .A3(n4512), .Y(n9432) );
  NAND4X0_LVT U2714 ( .A1(n2917), .A2(n2916), .A3(n2958), .A4(n1849), .Y(N693)
         );
  AND2X1_LVT U2715 ( .A1(n2959), .A2(n2960), .Y(n1849) );
  AND2X4_LVT U2716 ( .A1(n7911), .A2(n7910), .Y(n8105) );
  IBUFFX2_LVT U2717 ( .A(n2984), .Y(n4013) );
  IBUFFX4_LVT U2718 ( .A(n4013), .Y(n1875) );
  OA21X1_LVT U2719 ( .A1(n3163), .A2(n3987), .A3(n8781), .Y(n8784) );
  NOR2X0_LVT U2720 ( .A1(io_fpu_inst[6]), .A2(n3590), .Y(n5164) );
  AND3X1_LVT U2721 ( .A1(n8896), .A2(n8894), .A3(n1850), .Y(n8899) );
  OA21X1_LVT U2722 ( .A1(n3409), .A2(n2969), .A3(n8895), .Y(n1850) );
  NAND2X0_LVT U2723 ( .A1(n9529), .A2(n5071), .Y(n4504) );
  AND2X1_LVT U2724 ( .A1(n3590), .A2(n9524), .Y(n5071) );
  AND3X1_LVT U2725 ( .A1(n8590), .A2(n8589), .A3(n1851), .Y(n3725) );
  AOI22X1_LVT U2726 ( .A1(n_T_427[1010]), .A2(n3759), .A3(n1875), .A4(n1884), 
        .Y(n1851) );
  NAND3X0_LVT U2727 ( .A1(n2571), .A2(n3587), .A3(n1852), .Y(n4500) );
  AND3X1_LVT U2728 ( .A1(n3590), .A2(n9445), .A3(n9435), .Y(n1852) );
  NBUFFX2_LVT U2729 ( .A(n3077), .Y(n1853) );
  NBUFFX2_LVT U2730 ( .A(n3078), .Y(io_fpu_inst[30]) );
  NAND3X2_LVT U2731 ( .A1(n3773), .A2(n6954), .A3(n2068), .Y(n9014) );
  NAND3X0_LVT U2732 ( .A1(n8796), .A2(n8795), .A3(n1855), .Y(n8797) );
  NAND3X0_LVT U2733 ( .A1(n8194), .A2(n8195), .A3(n1856), .Y(n8196) );
  OA21X1_LVT U2734 ( .A1(n3460), .A2(n3751), .A3(n8193), .Y(n1856) );
  NBUFFX2_LVT U2735 ( .A(n3076), .Y(io_fpu_inst[3]) );
  NOR4X1_LVT U2736 ( .A1(n8797), .A2(n8789), .A3(n8790), .A4(n8798), .Y(n2365)
         );
  NAND4X1_LVT U2737 ( .A1(n9061), .A2(n9060), .A3(n2619), .A4(n9057), .Y(n2600) );
  NOR3X2_LVT U2738 ( .A1(n2600), .A2(n9063), .A3(n9062), .Y(n3750) );
  NAND3X2_LVT U2739 ( .A1(n5109), .A2(n5110), .A3(n9432), .Y(n6906) );
  AND2X1_LVT U2740 ( .A1(n3593), .A2(io_fpu_inst[4]), .Y(n3597) );
  OR3X1_LVT U2741 ( .A1(n7106), .A2(n1858), .A3(n7107), .Y(n7108) );
  NAND4X0_LVT U2742 ( .A1(n7102), .A2(n2587), .A3(n2588), .A4(n7101), .Y(n1858) );
  NBUFFX2_LVT U2743 ( .A(ibuf_io_inst_0_bits_raw[30]), .Y(n1859) );
  IBUFFX2_LVT U2744 ( .A(io_fpu_inst[31]), .Y(n2139) );
  AOI22X2_LVT U2745 ( .A1(n1861), .A2(n1860), .A3(n3606), .A4(n_T_427[1379]), 
        .Y(n8054) );
  IBUFFX2_LVT U2746 ( .A(n9006), .Y(n1860) );
  IBUFFX2_LVT U2747 ( .A(n3145), .Y(n1861) );
  AND3X1_LVT U2748 ( .A1(n4510), .A2(n2620), .A3(n5149), .Y(n2145) );
  NAND2X0_LVT U2749 ( .A1(n3582), .A2(n1862), .Y(n4506) );
  AND2X1_LVT U2750 ( .A1(n4505), .A2(n5086), .Y(n1862) );
  NBUFFX2_LVT U2751 ( .A(n2553), .Y(n1863) );
  AND3X2_LVT U2752 ( .A1(n2988), .A2(n2989), .A3(n8946), .Y(n1883) );
  NAND4X1_LVT U2753 ( .A1(n3634), .A2(n1883), .A3(n2530), .A4(n2987), .Y(N741)
         );
  IBUFFX32_LVT U2754 ( .A(n_T_427[1187]), .Y(n1864) );
  OR2X1_LVT U2755 ( .A1(n3663), .A2(n1864), .Y(n8076) );
  IBUFFX2_LVT U2756 ( .A(n3783), .Y(n2553) );
  NAND3X0_LVT U2757 ( .A1(n3766), .A2(n2925), .A3(n1865), .Y(N714) );
  AND3X1_LVT U2758 ( .A1(n3762), .A2(n2923), .A3(n2924), .Y(n1865) );
  AND3X1_LVT U2759 ( .A1(n2911), .A2(n8729), .A3(n1866), .Y(n2581) );
  AND2X1_LVT U2760 ( .A1(n8727), .A2(n8728), .Y(n1866) );
  IBUFFX2_LVT U2761 ( .A(n3692), .Y(n3987) );
  NAND2X0_LVT U2762 ( .A1(n2602), .A2(n8220), .Y(n2601) );
  OA22X1_LVT U2763 ( .A1(n2641), .A2(n2642), .A3(n5158), .A4(n5141), .Y(n2623)
         );
  NBUFFX2_LVT U2764 ( .A(n9104), .Y(n1867) );
  NAND2X0_LVT U2765 ( .A1(n8848), .A2(n1868), .Y(n2147) );
  NAND2X0_LVT U2766 ( .A1(n_T_427[825]), .A2(n9056), .Y(n1868) );
  NBUFFX2_LVT U2767 ( .A(n9022), .Y(n3643) );
  AND3X1_LVT U2768 ( .A1(n6966), .A2(n6965), .A3(n2548), .Y(n7911) );
  NBUFFX2_LVT U2769 ( .A(n9022), .Y(n3649) );
  NAND2X0_LVT U2770 ( .A1(n_T_427[228]), .A2(n3745), .Y(n8048) );
  NOR2X0_LVT U2771 ( .A1(n1869), .A2(n7974), .Y(n2129) );
  NAND3X0_LVT U2772 ( .A1(n7971), .A2(n7973), .A3(n7972), .Y(n1869) );
  AND2X1_LVT U2773 ( .A1(n7248), .A2(n1870), .Y(n1893) );
  NAND2X0_LVT U2774 ( .A1(n_T_427[1352]), .A2(n3603), .Y(n1870) );
  NAND2X0_LVT U2775 ( .A1(n_T_427[1717]), .A2(n3689), .Y(n8697) );
  AOI22X1_LVT U2776 ( .A1(n1872), .A2(n1871), .A3(n3628), .A4(n_T_427[1420]), 
        .Y(n7360) );
  INVX1_LVT U2777 ( .A(n2090), .Y(n1871) );
  INVX1_LVT U2778 ( .A(n3092), .Y(n1872) );
  NAND3X0_LVT U2779 ( .A1(n2884), .A2(n2898), .A3(n1873), .Y(N672) );
  AND3X1_LVT U2780 ( .A1(n2883), .A2(n2900), .A3(n2899), .Y(n1873) );
  NAND3X1_LVT U2781 ( .A1(n5075), .A2(io_fpu_inst[5]), .A3(n3597), .Y(n5076)
         );
  NAND2X0_LVT U2782 ( .A1(n_T_427[1647]), .A2(n3643), .Y(n8493) );
  AOI22X2_LVT U2783 ( .A1(n1875), .A2(n1874), .A3(n3761), .A4(n_T_427[989]), 
        .Y(n7859) );
  IBUFFX2_LVT U2784 ( .A(n3332), .Y(n1874) );
  NAND2X0_LVT U2785 ( .A1(n_T_427[298]), .A2(n3789), .Y(n8289) );
  NOR3X0_LVT U2786 ( .A1(n3076), .A2(n9111), .A3(io_fpu_inst[11]), .Y(n4503)
         );
  NAND2X0_LVT U2787 ( .A1(n_T_427[1657]), .A2(n3649), .Y(n8829) );
  NBUFFX2_LVT U2788 ( .A(n9522), .Y(io_fpu_inst[25]) );
  NAND4X0_LVT U2789 ( .A1(n2892), .A2(n2584), .A3(n2891), .A4(n1877), .Y(N690)
         );
  AND2X1_LVT U2790 ( .A1(n7273), .A2(n2936), .Y(n1877) );
  NAND3X0_LVT U2791 ( .A1(n2905), .A2(n2971), .A3(n1878), .Y(N694) );
  AND3X1_LVT U2792 ( .A1(n2970), .A2(n2972), .A3(n2904), .Y(n1878) );
  NAND2X0_LVT U2793 ( .A1(n5119), .A2(n1879), .Y(n5111) );
  AND2X1_LVT U2794 ( .A1(n9089), .A2(csr_io_decode_0_write_illegal), .Y(n1879)
         );
  NAND4X0_LVT U2795 ( .A1(n3008), .A2(n3071), .A3(n3007), .A4(n1880), .Y(N698)
         );
  AND2X1_LVT U2796 ( .A1(n3070), .A2(n3069), .Y(n1880) );
  NAND3X0_LVT U2797 ( .A1(n2907), .A2(n2976), .A3(n1881), .Y(N686) );
  AND3X1_LVT U2798 ( .A1(n2975), .A2(n2906), .A3(n2977), .Y(n1881) );
  NBUFFX2_LVT U2799 ( .A(n9525), .Y(io_fpu_inst[6]) );
  NBUFFX2_LVT U2800 ( .A(n9528), .Y(n3077) );
  OR4X2_LVT U2801 ( .A1(n5099), .A2(n3077), .A3(n2537), .A4(io_fpu_inst[6]), 
        .Y(n2634) );
  IBUFFX2_LVT U2802 ( .A(n9528), .Y(n3578) );
  NAND4X0_LVT U2803 ( .A1(n8834), .A2(n8832), .A3(n8833), .A4(n1882), .Y(n8835) );
  OR2X1_LVT U2804 ( .A1(n3366), .A2(n4011), .Y(n1882) );
  AND2X1_LVT U2805 ( .A1(n3765), .A2(n6923), .Y(n2983) );
  NAND2X0_LVT U2806 ( .A1(n_T_427[1641]), .A2(n3649), .Y(n8272) );
  IBUFFX2_LVT U2807 ( .A(n3353), .Y(n1884) );
  OA21X1_LVT U2808 ( .A1(n3584), .A2(n1885), .A3(n5076), .Y(n3072) );
  AND2X1_LVT U2809 ( .A1(n9076), .A2(n3585), .Y(n1885) );
  NAND3X0_LVT U2810 ( .A1(n3014), .A2(n3694), .A3(n1886), .Y(N705) );
  AND3X1_LVT U2811 ( .A1(n3013), .A2(n3693), .A3(n3695), .Y(n1886) );
  NAND3X0_LVT U2812 ( .A1(n3016), .A2(n3699), .A3(n1887), .Y(N706) );
  AND3X1_LVT U2813 ( .A1(n3015), .A2(n3698), .A3(n3700), .Y(n1887) );
  NBUFFX2_LVT U2814 ( .A(n9528), .Y(n3076) );
  NAND4X1_LVT U2815 ( .A1(n2167), .A2(n2168), .A3(n2932), .A4(n1888), .Y(N722)
         );
  NAND4X0_LVT U2816 ( .A1(n2896), .A2(n2942), .A3(n2895), .A4(n1889), .Y(N683)
         );
  AND2X1_LVT U2817 ( .A1(n2943), .A2(n2944), .Y(n1889) );
  NAND4X0_LVT U2818 ( .A1(n2890), .A2(n2939), .A3(n2889), .A4(n1890), .Y(N692)
         );
  AND2X1_LVT U2819 ( .A1(n2941), .A2(n2940), .Y(n1890) );
  NBUFFX2_LVT U2820 ( .A(n3593), .Y(n1891) );
  AND2X1_LVT U2821 ( .A1(n2561), .A2(n6922), .Y(n3709) );
  AND3X1_LVT U2822 ( .A1(n7247), .A2(n7246), .A3(n1893), .Y(n1892) );
  OA21X1_LVT U2823 ( .A1(n3305), .A2(n1894), .A3(n8955), .Y(n8958) );
  IBUFFX4_LVT U2824 ( .A(n3768), .Y(n1894) );
  OA21X1_LVT U2825 ( .A1(n3339), .A2(n1894), .A3(n8250), .Y(n8253) );
  OA21X1_LVT U2826 ( .A1(n3346), .A2(n1894), .A3(n8446), .Y(n8449) );
  OA21X1_LVT U2827 ( .A1(n3365), .A2(n1894), .A3(n8828), .Y(n8831) );
  OA21X2_LVT U2828 ( .A1(n3349), .A2(n1894), .A3(n8510), .Y(n8513) );
  AND3X1_LVT U2829 ( .A1(n2962), .A2(n2961), .A3(n1895), .Y(n2945) );
  AND3X1_LVT U2830 ( .A1(n8480), .A2(n8479), .A3(n1896), .Y(n1895) );
  AOI22X1_LVT U2831 ( .A1(n_T_427[1135]), .A2(n3668), .A3(n3635), .A4(
        n_T_427[1263]), .Y(n1896) );
  AND4X1_LVT U2832 ( .A1(n7132), .A2(n1899), .A3(n7134), .A4(n7133), .Y(n1898)
         );
  IBUFFX32_LVT U2833 ( .A(n3424), .Y(n1897) );
  AND2X1_LVT U2834 ( .A1(n3599), .A2(n1898), .Y(n1901) );
  NAND2X0_LVT U2835 ( .A1(n1897), .A2(n3768), .Y(n1899) );
  IBUFFX4_LVT U2836 ( .A(n3768), .Y(n4010) );
  OA22X1_LVT U2837 ( .A1(n3189), .A2(n4016), .A3(n3432), .A4(n2081), .Y(n1900)
         );
  NAND4X0_LVT U2838 ( .A1(n2886), .A2(n2885), .A3(n3598), .A4(n1901), .Y(N685)
         );
  NAND2X0_LVT U2839 ( .A1(n1902), .A2(n2909), .Y(N682) );
  AND3X1_LVT U2840 ( .A1(n2978), .A2(n2908), .A3(n1903), .Y(n1902) );
  AND3X1_LVT U2841 ( .A1(n2979), .A2(n7044), .A3(n1904), .Y(n1903) );
  AND2X1_LVT U2842 ( .A1(n7046), .A2(n1905), .Y(n1904) );
  OA21X1_LVT U2843 ( .A1(n3419), .A2(n3663), .A3(n7045), .Y(n1905) );
  NAND4X0_LVT U2844 ( .A1(n3778), .A2(n1907), .A3(n2949), .A4(n1906), .Y(N721)
         );
  AND2X1_LVT U2845 ( .A1(n2948), .A2(n3754), .Y(n1906) );
  AND4X1_LVT U2846 ( .A1(n1909), .A2(n8255), .A3(n1908), .A4(n8256), .Y(n1907)
         );
  AND2X1_LVT U2847 ( .A1(n8254), .A2(n8252), .Y(n1908) );
  AND2X1_LVT U2848 ( .A1(n8251), .A2(n8253), .Y(n1909) );
  NAND4X0_LVT U2849 ( .A1(n2888), .A2(n2887), .A3(n2938), .A4(n1910), .Y(N695)
         );
  AND2X1_LVT U2850 ( .A1(n1912), .A2(n1911), .Y(n1910) );
  AND4X1_LVT U2851 ( .A1(n7411), .A2(n1913), .A3(n7414), .A4(n7412), .Y(n1911)
         );
  AND3X1_LVT U2852 ( .A1(n7416), .A2(n7415), .A3(n7413), .Y(n1912) );
  OA22X1_LVT U2853 ( .A1(n4016), .A2(n3093), .A3(n3443), .A4(n4009), .Y(n1913)
         );
  AND3X2_LVT U2854 ( .A1(n2677), .A2(io_fpu_inst[14]), .A3(n9231), .Y(n9087)
         );
  AND3X2_LVT U2855 ( .A1(n9412), .A2(n9099), .A3(n5167), .Y(n2677) );
  NAND4X0_LVT U2856 ( .A1(n4765), .A2(n6924), .A3(n4764), .A4(n4763), .Y(n4766) );
  NAND3X0_LVT U2857 ( .A1(n1914), .A2(n1915), .A3(n1916), .Y(n4852) );
  OR4X1_LVT U2858 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .Y(n1914)
         );
  OR4X1_LVT U2859 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .Y(n1915)
         );
  AND4X1_LVT U2860 ( .A1(n4780), .A2(io_fpu_dec_ren1), .A3(n4779), .A4(n9286), 
        .Y(n1916) );
  NAND4X1_LVT U2861 ( .A1(n4954), .A2(n4955), .A3(n4953), .A4(n4952), .Y(n1917) );
  NBUFFX2_LVT U2862 ( .A(n6810), .Y(n1918) );
  NBUFFX2_LVT U2863 ( .A(n6810), .Y(n1919) );
  AND2X1_LVT U2864 ( .A1(n2981), .A2(n3864), .Y(n6829) );
  OR2X2_LVT U2865 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(
        ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n4814) );
  OA22X1_LVT U2866 ( .A1(n3162), .A2(n1994), .A3(n3514), .A4(n3800), .Y(n6676)
         );
  AND4X1_LVT U2867 ( .A1(n1920), .A2(n1921), .A3(n1922), .A4(n1923), .Y(n6458)
         );
  AOI22X2_LVT U2868 ( .A1(n3829), .A2(n_T_427[1835]), .A3(n_T_427[1710]), .A4(
        n3825), .Y(n1920) );
  AOI22X2_LVT U2869 ( .A1(n3893), .A2(n_T_427[1582]), .A3(n_T_427[1646]), .A4(
        n3887), .Y(n1921) );
  AOI22X2_LVT U2870 ( .A1(n3925), .A2(n_T_427[1518]), .A3(n_T_427[1390]), .A4(
        n3919), .Y(n1922) );
  AOI22X2_LVT U2871 ( .A1(n3935), .A2(n_T_427[1454]), .A3(n_T_427[1326]), .A4(
        n3930), .Y(n1923) );
  AND4X1_LVT U2872 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .Y(n6317)
         );
  AOI22X2_LVT U2873 ( .A1(n3830), .A2(n_T_427[1829]), .A3(n_T_427[1704]), .A4(
        n3825), .Y(n1924) );
  AOI22X2_LVT U2874 ( .A1(n3892), .A2(n_T_427[1576]), .A3(n_T_427[1640]), .A4(
        n3887), .Y(n1925) );
  AOI22X2_LVT U2875 ( .A1(n3925), .A2(n_T_427[1512]), .A3(n_T_427[1384]), .A4(
        n3919), .Y(n1926) );
  AOI22X2_LVT U2876 ( .A1(n3935), .A2(n_T_427[1448]), .A3(n_T_427[1320]), .A4(
        n3929), .Y(n1927) );
  AND4X1_LVT U2877 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .Y(n6204)
         );
  AOI22X2_LVT U2878 ( .A1(n3829), .A2(n_T_427[1824]), .A3(n_T_427[1699]), .A4(
        n3825), .Y(n1928) );
  AOI22X1_LVT U2879 ( .A1(n3892), .A2(n_T_427[1571]), .A3(n_T_427[1635]), .A4(
        n3886), .Y(n1929) );
  AOI22X1_LVT U2880 ( .A1(n3924), .A2(n_T_427[1507]), .A3(n_T_427[1379]), .A4(
        n3919), .Y(n1930) );
  AOI22X1_LVT U2881 ( .A1(n3934), .A2(n_T_427[1443]), .A3(n_T_427[1315]), .A4(
        n3929), .Y(n1931) );
  AND4X1_LVT U2882 ( .A1(n1932), .A2(n1933), .A3(n1934), .A4(n1935), .Y(n6409)
         );
  AOI22X2_LVT U2883 ( .A1(n3830), .A2(n_T_427[1833]), .A3(n_T_427[1708]), .A4(
        n3825), .Y(n1932) );
  AOI22X2_LVT U2884 ( .A1(n3893), .A2(n_T_427[1580]), .A3(n_T_427[1644]), .A4(
        n3888), .Y(n1933) );
  AOI22X2_LVT U2885 ( .A1(n3925), .A2(n_T_427[1516]), .A3(n_T_427[1388]), .A4(
        n3919), .Y(n1934) );
  AOI22X2_LVT U2886 ( .A1(n3935), .A2(n_T_427[1452]), .A3(n_T_427[1324]), .A4(
        n3930), .Y(n1935) );
  AND4X1_LVT U2887 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .Y(n6363)
         );
  AOI22X2_LVT U2888 ( .A1(n3829), .A2(n_T_427[1831]), .A3(n_T_427[1706]), .A4(
        n3825), .Y(n1936) );
  AOI22X2_LVT U2889 ( .A1(n3893), .A2(n_T_427[1578]), .A3(n_T_427[1642]), .A4(
        n3887), .Y(n1937) );
  AOI22X2_LVT U2890 ( .A1(n3925), .A2(n_T_427[1514]), .A3(n_T_427[1386]), .A4(
        n3920), .Y(n1938) );
  AOI22X2_LVT U2891 ( .A1(n3935), .A2(n_T_427[1450]), .A3(n_T_427[1322]), .A4(
        n3929), .Y(n1939) );
  AND4X1_LVT U2892 ( .A1(n1940), .A2(n1941), .A3(n1942), .A4(n1943), .Y(n6225)
         );
  AOI22X2_LVT U2893 ( .A1(n3829), .A2(n_T_427[1825]), .A3(n_T_427[1700]), .A4(
        n3825), .Y(n1940) );
  AOI22X2_LVT U2894 ( .A1(n3892), .A2(n_T_427[1572]), .A3(n_T_427[1636]), .A4(
        n3887), .Y(n1941) );
  AOI22X1_LVT U2895 ( .A1(n3924), .A2(n_T_427[1508]), .A3(n_T_427[1380]), .A4(
        n3919), .Y(n1942) );
  AOI22X1_LVT U2896 ( .A1(n3934), .A2(n_T_427[1444]), .A3(n_T_427[1316]), .A4(
        n3929), .Y(n1943) );
  AOI22X1_LVT U2897 ( .A1(n3801), .A2(n_T_427[1864]), .A3(n_T_427[1746]), .A4(
        n2866), .Y(n1988) );
  AND4X1_LVT U2898 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(n1947), .Y(n6012)
         );
  AOI22X1_LVT U2899 ( .A1(n1918), .A2(n_T_427[347]), .A3(n_T_427[539]), .A4(
        n3819), .Y(n1944) );
  AOI22X1_LVT U2900 ( .A1(n3912), .A2(n_T_427[475]), .A3(n_T_427[922]), .A4(
        n3896), .Y(n1945) );
  AOI22X1_LVT U2901 ( .A1(n3914), .A2(n_T_427[27]), .A3(n_T_427[155]), .A4(
        n2863), .Y(n1946) );
  AND3X1_LVT U2902 ( .A1(n6005), .A2(n6004), .A3(n6003), .Y(n1947) );
  AND4X1_LVT U2903 ( .A1(n1948), .A2(n1949), .A3(n1950), .A4(n1951), .Y(n6532)
         );
  AOI22X1_LVT U2904 ( .A1(n2765), .A2(n_T_427[1838]), .A3(n_T_427[1713]), .A4(
        n3824), .Y(n1948) );
  AOI22X2_LVT U2905 ( .A1(n3893), .A2(n_T_427[1585]), .A3(n_T_427[1649]), .A4(
        n3887), .Y(n1949) );
  AOI22X2_LVT U2906 ( .A1(n3925), .A2(n_T_427[1521]), .A3(n_T_427[1393]), .A4(
        n3920), .Y(n1950) );
  AOI22X2_LVT U2907 ( .A1(n3935), .A2(n_T_427[1457]), .A3(n_T_427[1329]), .A4(
        n3929), .Y(n1951) );
  AND4X1_LVT U2908 ( .A1(n1952), .A2(n1953), .A3(n1954), .A4(n1955), .Y(n6609)
         );
  AOI22X1_LVT U2909 ( .A1(n2765), .A2(n_T_427[1841]), .A3(n_T_427[1716]), .A4(
        n3824), .Y(n1952) );
  AOI22X2_LVT U2910 ( .A1(n3893), .A2(n_T_427[1588]), .A3(n_T_427[1652]), .A4(
        n3888), .Y(n1953) );
  AOI22X2_LVT U2911 ( .A1(n3926), .A2(n_T_427[1524]), .A3(n_T_427[1396]), .A4(
        n3920), .Y(n1954) );
  AOI22X2_LVT U2912 ( .A1(n3936), .A2(n_T_427[1460]), .A3(n_T_427[1332]), .A4(
        n3930), .Y(n1955) );
  AND4X1_LVT U2913 ( .A1(n1956), .A2(n1957), .A3(n1958), .A4(n1959), .Y(n6702)
         );
  AOI22X1_LVT U2914 ( .A1(n2765), .A2(n_T_427[1844]), .A3(n_T_427[1720]), .A4(
        n3824), .Y(n1956) );
  AOI22X2_LVT U2915 ( .A1(n3893), .A2(n_T_427[1592]), .A3(n_T_427[1656]), .A4(
        n3888), .Y(n1957) );
  AOI22X2_LVT U2916 ( .A1(n3926), .A2(n_T_427[1528]), .A3(n_T_427[1400]), .A4(
        n3921), .Y(n1958) );
  AOI22X2_LVT U2917 ( .A1(n3936), .A2(n_T_427[1464]), .A3(n_T_427[1336]), .A4(
        n3930), .Y(n1959) );
  AND4X1_LVT U2918 ( .A1(n1960), .A2(n1961), .A3(n1962), .A4(n1963), .Y(n6850)
         );
  AOI22X1_LVT U2919 ( .A1(n2765), .A2(n_T_427[1847]), .A3(n_T_427[1725]), .A4(
        n3827), .Y(n1960) );
  AOI22X2_LVT U2920 ( .A1(n3894), .A2(n_T_427[1597]), .A3(n_T_427[1661]), .A4(
        n3888), .Y(n1961) );
  AOI22X2_LVT U2921 ( .A1(n3926), .A2(n_T_427[1533]), .A3(n_T_427[1405]), .A4(
        n3920), .Y(n1962) );
  AOI22X2_LVT U2922 ( .A1(n3936), .A2(n_T_427[1469]), .A3(n_T_427[1341]), .A4(
        n3929), .Y(n1963) );
  AND4X1_LVT U2923 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .Y(n5947)
         );
  AOI22X1_LVT U2924 ( .A1(n2765), .A2(n_T_427[1813]), .A3(n_T_427[1687]), .A4(
        n3826), .Y(n1964) );
  AOI22X2_LVT U2925 ( .A1(n3892), .A2(n_T_427[1559]), .A3(n_T_427[1623]), .A4(
        n3887), .Y(n1965) );
  AOI22X2_LVT U2926 ( .A1(n3924), .A2(n_T_427[1495]), .A3(n_T_427[1367]), .A4(
        n3918), .Y(n1966) );
  AOI22X2_LVT U2927 ( .A1(n3934), .A2(n_T_427[1431]), .A3(n_T_427[1303]), .A4(
        n3928), .Y(n1967) );
  AND4X1_LVT U2928 ( .A1(n1968), .A2(n1969), .A3(n1970), .A4(n1971), .Y(n6292)
         );
  AOI22X1_LVT U2929 ( .A1(n2765), .A2(n_T_427[1828]), .A3(n_T_427[1703]), .A4(
        n3825), .Y(n1968) );
  AOI22X2_LVT U2930 ( .A1(n3892), .A2(n_T_427[1575]), .A3(n_T_427[1639]), .A4(
        n3887), .Y(n1969) );
  AOI22X2_LVT U2931 ( .A1(n3925), .A2(n_T_427[1511]), .A3(n_T_427[1383]), .A4(
        n3919), .Y(n1970) );
  AOI22X2_LVT U2932 ( .A1(n3935), .A2(n_T_427[1447]), .A3(n_T_427[1319]), .A4(
        n3929), .Y(n1971) );
  AND4X1_LVT U2933 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .Y(n6629)
         );
  AOI22X1_LVT U2934 ( .A1(n2765), .A2(n_T_427[1842]), .A3(n_T_427[1717]), .A4(
        n3824), .Y(n1972) );
  AOI22X2_LVT U2935 ( .A1(n3893), .A2(n_T_427[1589]), .A3(n_T_427[1653]), .A4(
        n3888), .Y(n1973) );
  AOI22X2_LVT U2936 ( .A1(n3926), .A2(n_T_427[1525]), .A3(n_T_427[1397]), .A4(
        n3921), .Y(n1974) );
  AOI22X2_LVT U2937 ( .A1(n3936), .A2(n_T_427[1461]), .A3(n_T_427[1333]), .A4(
        n3930), .Y(n1975) );
  AND4X1_LVT U2938 ( .A1(n1976), .A2(n1977), .A3(n1978), .A4(n1979), .Y(n6342)
         );
  AOI22X1_LVT U2939 ( .A1(n2765), .A2(n_T_427[1830]), .A3(n_T_427[1705]), .A4(
        n3825), .Y(n1976) );
  AOI22X2_LVT U2940 ( .A1(n3893), .A2(n_T_427[1577]), .A3(n_T_427[1641]), .A4(
        n3887), .Y(n1977) );
  AOI22X2_LVT U2941 ( .A1(n3925), .A2(n_T_427[1513]), .A3(n_T_427[1385]), .A4(
        n3920), .Y(n1978) );
  AOI22X2_LVT U2942 ( .A1(n3935), .A2(n_T_427[1449]), .A3(n_T_427[1321]), .A4(
        n3929), .Y(n1979) );
  AND4X1_LVT U2943 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .Y(n5923)
         );
  AOI22X1_LVT U2944 ( .A1(n2028), .A2(n_T_427[1867]), .A3(n_T_427[1750]), .A4(
        n2868), .Y(n1980) );
  AOI22X1_LVT U2945 ( .A1(n2765), .A2(n_T_427[1812]), .A3(n_T_427[1686]), .A4(
        n3825), .Y(n1981) );
  AOI22X1_LVT U2946 ( .A1(n3891), .A2(n_T_427[1558]), .A3(n_T_427[1622]), .A4(
        n3886), .Y(n1982) );
  AOI22X2_LVT U2947 ( .A1(n5911), .A2(n6877), .A3(n_T_427[1904]), .A4(n3884), 
        .Y(n1983) );
  AND4X1_LVT U2948 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .Y(n5724)
         );
  AOI22X2_LVT U2949 ( .A1(n6764), .A2(n_T_427[1859]), .A3(n_T_427[1740]), .A4(
        n2866), .Y(n1984) );
  AOI22X2_LVT U2950 ( .A1(n3828), .A2(n_T_427[1803]), .A3(n_T_427[1676]), .A4(
        n3827), .Y(n1985) );
  AOI22X1_LVT U2951 ( .A1(n3891), .A2(n_T_427[1548]), .A3(n_T_427[1612]), .A4(
        n3885), .Y(n1986) );
  AOI22X2_LVT U2952 ( .A1(n3923), .A2(n_T_427[1484]), .A3(n_T_427[1356]), .A4(
        n3918), .Y(n1987) );
  AND4X1_LVT U2953 ( .A1(n1988), .A2(n1989), .A3(n1990), .A4(n1991), .Y(n2429)
         );
  AOI22X1_LVT U2954 ( .A1(n2765), .A2(n_T_427[1808]), .A3(n_T_427[1682]), .A4(
        n3825), .Y(n1989) );
  AOI22X2_LVT U2955 ( .A1(n3886), .A2(n_T_427[1618]), .A3(n_T_427[1554]), .A4(
        n3891), .Y(n1990) );
  AOI22X2_LVT U2956 ( .A1(n3918), .A2(n_T_427[1362]), .A3(n_T_427[1490]), .A4(
        n3924), .Y(n1991) );
  INVX1_LVT U2957 ( .A(n3586), .Y(n1992) );
  NBUFFX2_LVT U2958 ( .A(n3877), .Y(n1993) );
  AND2X1_LVT U2959 ( .A1(n5434), .A2(n6238), .Y(n2981) );
  NBUFFX2_LVT U2960 ( .A(n2875), .Y(n1994) );
  NBUFFX2_LVT U2961 ( .A(n2875), .Y(n3080) );
  AND4X1_LVT U2962 ( .A1(n1995), .A2(n1996), .A3(n1997), .A4(n1998), .Y(n6096)
         );
  AOI22X2_LVT U2963 ( .A1(n2866), .A2(n_T_427[1758]), .A3(n_T_427[1820]), .A4(
        n3830), .Y(n1995) );
  AOI22X1_LVT U2964 ( .A1(n_T_427[1873]), .A2(n3801), .A3(n3884), .A4(
        n_T_427[1912]), .Y(n1996) );
  AOI22X1_LVT U2965 ( .A1(n3826), .A2(n_T_427[1694]), .A3(n_T_427[1566]), .A4(
        n3890), .Y(n1997) );
  AOI22X1_LVT U2966 ( .A1(n3889), .A2(n_T_427[1630]), .A3(n_T_427[1502]), .A4(
        n3922), .Y(n1998) );
  AND4X1_LVT U2967 ( .A1(n1999), .A2(n2000), .A3(n2001), .A4(n2002), .Y(n5876)
         );
  AOI22X1_LVT U2968 ( .A1(n2868), .A2(n_T_427[1748]), .A3(n_T_427[1810]), .A4(
        n3829), .Y(n1999) );
  AOI22X1_LVT U2969 ( .A1(n_T_427[1866]), .A2(n6764), .A3(n3884), .A4(
        n_T_427[1902]), .Y(n2000) );
  AOI22X1_LVT U2970 ( .A1(n3827), .A2(n_T_427[1684]), .A3(n_T_427[1556]), .A4(
        n3890), .Y(n2001) );
  AOI22X2_LVT U2971 ( .A1(n3888), .A2(n_T_427[1620]), .A3(n_T_427[1492]), .A4(
        n3922), .Y(n2002) );
  AND4X1_LVT U2972 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .Y(n5991)
         );
  AOI22X2_LVT U2973 ( .A1(n2866), .A2(n_T_427[1753]), .A3(n_T_427[1815]), .A4(
        n3830), .Y(n2003) );
  AOI22X1_LVT U2974 ( .A1(n3802), .A2(n_T_427[1869]), .A3(n3884), .A4(
        n_T_427[1907]), .Y(n2004) );
  AOI22X1_LVT U2975 ( .A1(n3827), .A2(n_T_427[1689]), .A3(n_T_427[1561]), .A4(
        n3890), .Y(n2005) );
  AOI22X1_LVT U2976 ( .A1(n3889), .A2(n_T_427[1625]), .A3(n_T_427[1497]), .A4(
        n3922), .Y(n2006) );
  AND4X1_LVT U2977 ( .A1(n2007), .A2(n2008), .A3(n2009), .A4(n2010), .Y(n5763)
         );
  AOI22X1_LVT U2978 ( .A1(n3801), .A2(n_T_427[1861]), .A3(n_T_427[1742]), .A4(
        n2868), .Y(n2007) );
  AOI22X1_LVT U2979 ( .A1(n2765), .A2(n_T_427[1805]), .A3(n_T_427[1678]), .A4(
        n3824), .Y(n2008) );
  AOI22X1_LVT U2980 ( .A1(n3892), .A2(n_T_427[1550]), .A3(n_T_427[1614]), .A4(
        n3886), .Y(n2009) );
  AOI22X2_LVT U2981 ( .A1(n3924), .A2(n_T_427[1486]), .A3(n_T_427[1358]), .A4(
        n3918), .Y(n2010) );
  AND4X1_LVT U2982 ( .A1(n2011), .A2(n2012), .A3(n2013), .A4(n2014), .Y(n2290)
         );
  AOI22X2_LVT U2983 ( .A1(n2866), .A2(n_T_427[1755]), .A3(n_T_427[1817]), .A4(
        n2765), .Y(n2011) );
  AOI22X1_LVT U2984 ( .A1(n_T_427[1871]), .A2(n6764), .A3(n3884), .A4(
        n_T_427[1909]), .Y(n2012) );
  AOI22X1_LVT U2985 ( .A1(n3827), .A2(n_T_427[1691]), .A3(n_T_427[1563]), .A4(
        n3890), .Y(n2013) );
  AOI22X2_LVT U2986 ( .A1(n3922), .A2(n_T_427[1499]), .A3(n_T_427[1627]), .A4(
        n3887), .Y(n2014) );
  AND4X1_LVT U2987 ( .A1(n2015), .A2(n2016), .A3(n2017), .A4(n2018), .Y(n2229)
         );
  AOI22X1_LVT U2988 ( .A1(n3802), .A2(n_T_427[1850]), .A3(n_T_427[1731]), .A4(
        n3798), .Y(n2015) );
  AOI22X1_LVT U2989 ( .A1(n2765), .A2(n_T_427[1794]), .A3(n_T_427[1667]), .A4(
        n3826), .Y(n2016) );
  AOI22X1_LVT U2990 ( .A1(n3891), .A2(n_T_427[1539]), .A3(n_T_427[1603]), .A4(
        n3885), .Y(n2017) );
  AOI22X1_LVT U2991 ( .A1(n5534), .A2(n1992), .A3(n_T_427[1885]), .A4(n3884), 
        .Y(n2018) );
  AND4X1_LVT U2992 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .Y(n2249)
         );
  AOI22X2_LVT U2993 ( .A1(n2866), .A2(n_T_427[1765]), .A3(n_T_427[1826]), .A4(
        n2765), .Y(n2019) );
  AOI22X1_LVT U2994 ( .A1(n_T_427[1877]), .A2(n3802), .A3(n3884), .A4(
        n_T_427[1918]), .Y(n2020) );
  AOI22X1_LVT U2995 ( .A1(n3827), .A2(n_T_427[1701]), .A3(n_T_427[1573]), .A4(
        n3890), .Y(n2021) );
  AOI22X2_LVT U2996 ( .A1(n3922), .A2(n_T_427[1509]), .A3(n_T_427[1637]), .A4(
        n3889), .Y(n2022) );
  AND4X1_LVT U2997 ( .A1(n2023), .A2(n2024), .A3(n2025), .A4(n2026), .Y(n6158)
         );
  AOI22X1_LVT U2998 ( .A1(n3802), .A2(n_T_427[1875]), .A3(n_T_427[1761]), .A4(
        n2868), .Y(n2023) );
  AOI22X1_LVT U2999 ( .A1(n6146), .A2(n6877), .A3(n3884), .A4(n_T_427[1914]), 
        .Y(n2024) );
  AOI22X2_LVT U3000 ( .A1(n3829), .A2(n_T_427[1822]), .A3(n_T_427[1697]), .A4(
        n3825), .Y(n2025) );
  AOI22X1_LVT U3001 ( .A1(n3892), .A2(n_T_427[1569]), .A3(n_T_427[1633]), .A4(
        n3886), .Y(n2026) );
  NBUFFX2_LVT U3002 ( .A(n2875), .Y(n2027) );
  INVX1_LVT U3003 ( .A(n2875), .Y(n2028) );
  IBUFFX2_LVT U3004 ( .A(io_dmem_resp_bits_tag[0]), .Y(n2029) );
  NBUFFX2_LVT U3005 ( .A(io_dmem_resp_valid), .Y(n2030) );
  NAND3X0_LVT U3006 ( .A1(n9390), .A2(n2152), .A3(n2573), .Y(n9395) );
  IBUFFX2_LVT U3007 ( .A(n3883), .Y(n3881) );
  IBUFFX2_LVT U3008 ( .A(n3883), .Y(n3882) );
  AOI22X2_LVT U3009 ( .A1(n3828), .A2(n_T_427[1809]), .A3(n_T_427[1683]), .A4(
        n3827), .Y(n2800) );
  IBUFFX2_LVT U3010 ( .A(n3082), .Y(n3824) );
  IBUFFX2_LVT U3011 ( .A(n3082), .Y(n3827) );
  IBUFFX2_LVT U3012 ( .A(n4969), .Y(n4748) );
  NAND2X4_LVT U3013 ( .A1(n6238), .A2(n3579), .Y(n3803) );
  AND3X1_LVT U3014 ( .A1(n2031), .A2(n2032), .A3(n2033), .Y(n2035) );
  AOI22X1_LVT U3015 ( .A1(n3891), .A2(n_T_427[1549]), .A3(n_T_427[1613]), .A4(
        n3886), .Y(n2031) );
  AOI22X2_LVT U3016 ( .A1(n1992), .A2(n5736), .A3(n_T_427[1895]), .A4(n3884), 
        .Y(n2032) );
  AOI22X1_LVT U3017 ( .A1(n2765), .A2(n_T_427[1804]), .A3(n_T_427[1677]), .A4(
        n3826), .Y(n2033) );
  NBUFFX2_LVT U3018 ( .A(n5453), .Y(n2034) );
  AND2X1_LVT U3019 ( .A1(n4901), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5453) );
  IBUFFX2_LVT U3020 ( .A(n6898), .Y(n3596) );
  IBUFFX2_LVT U3021 ( .A(n3195), .Y(n4359) );
  AOI21X2_LVT U3022 ( .A1(n3843), .A2(csr_io_rw_rdata[14]), .A3(n5731), .Y(
        n3195) );
  AND2X4_LVT U3023 ( .A1(n4970), .A2(n4752), .Y(n6948) );
  AND2X4_LVT U3024 ( .A1(n6948), .A2(n6956), .Y(n9041) );
  AND2X4_LVT U3025 ( .A1(n6948), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n9039) );
  OR2X2_LVT U3026 ( .A1(n2877), .A2(ibuf_io_inst_0_bits_inst_rs1[0]), .Y(n4969) );
  OR2X2_LVT U3027 ( .A1(ibuf_io_inst_0_bits_inst_rs2[3]), .A2(n4880), .Y(n6423) );
  NBUFFX2_LVT U3028 ( .A(n3040), .Y(n2036) );
  AND2X4_LVT U3029 ( .A1(n2036), .A2(n2061), .Y(n9389) );
  AND2X4_LVT U3030 ( .A1(n2036), .A2(n3042), .Y(n9393) );
  IBUFFX2_LVT U3031 ( .A(n3042), .Y(n2037) );
  DELLN3X2_LVT U3032 ( .A(n2037), .Y(n2061) );
  NBUFFX2_LVT U3033 ( .A(ibuf_io_inst_0_bits_inst_rs1[2]), .Y(n2038) );
  AND2X4_LVT U3034 ( .A1(n4748), .A2(n4752), .Y(n6957) );
  AND3X1_LVT U3035 ( .A1(n2039), .A2(n2040), .A3(n2041), .Y(n2108) );
  AND4X1_LVT U3036 ( .A1(n8184), .A2(n8182), .A3(n8183), .A4(n2612), .Y(n2039)
         );
  AND2X1_LVT U3037 ( .A1(n8170), .A2(n8169), .Y(n2040) );
  AND3X1_LVT U3038 ( .A1(n8181), .A2(n8180), .A3(n8179), .Y(n2041) );
  OA21X1_LVT U3039 ( .A1(n3144), .A2(n2120), .A3(n7935), .Y(n7936) );
  AND3X1_LVT U3040 ( .A1(n2042), .A2(n2043), .A3(n2044), .Y(n3743) );
  AND3X1_LVT U3041 ( .A1(n8458), .A2(n2589), .A3(n8459), .Y(n2042) );
  AND3X1_LVT U3042 ( .A1(n8465), .A2(n8464), .A3(n8463), .Y(n2043) );
  AND2X1_LVT U3043 ( .A1(n8461), .A2(n8460), .Y(n2044) );
  OA21X1_LVT U3044 ( .A1(n3146), .A2(n3767), .A3(n8101), .Y(n8104) );
  NAND3X0_LVT U3045 ( .A1(n2045), .A2(n2046), .A3(n2047), .Y(N696) );
  AND3X1_LVT U3046 ( .A1(n2086), .A2(n2087), .A3(n2088), .Y(n2045) );
  AND3X1_LVT U3047 ( .A1(n7420), .A2(n7419), .A3(n7418), .Y(n2046) );
  AND3X1_LVT U3048 ( .A1(n7424), .A2(n7423), .A3(n7422), .Y(n2047) );
  AND2X1_LVT U3049 ( .A1(n8994), .A2(n_T_427[122]), .Y(n2149) );
  NAND3X2_LVT U3050 ( .A1(n4497), .A2(n6916), .A3(n6915), .Y(n2627) );
  AND3X1_LVT U3051 ( .A1(n2048), .A2(n2049), .A3(n2050), .Y(n2173) );
  AND4X1_LVT U3052 ( .A1(n8564), .A2(n8562), .A3(n2603), .A4(n2593), .Y(n2048)
         );
  AND3X1_LVT U3053 ( .A1(n8560), .A2(n8559), .A3(n8558), .Y(n2049) );
  AND3X1_LVT U3054 ( .A1(n8554), .A2(n8555), .A3(n8556), .Y(n2050) );
  AND2X1_LVT U3055 ( .A1(n2051), .A2(n2052), .Y(n2160) );
  AND3X1_LVT U3056 ( .A1(n8381), .A2(n8380), .A3(n8379), .Y(n2051) );
  AND3X1_LVT U3057 ( .A1(n8384), .A2(n8382), .A3(n2604), .Y(n2052) );
  AND2X1_LVT U3058 ( .A1(n2053), .A2(n2054), .Y(n2543) );
  AND3X1_LVT U3059 ( .A1(n8365), .A2(n8364), .A3(n8363), .Y(n2053) );
  AND3X1_LVT U3060 ( .A1(n8361), .A2(n8360), .A3(n8359), .Y(n2054) );
  NAND3X1_LVT U3061 ( .A1(n4497), .A2(n6915), .A3(n6916), .Y(n6962) );
  NAND3X0_LVT U3062 ( .A1(n5166), .A2(n3049), .A3(n5110), .Y(n3075) );
  AND2X1_LVT U3063 ( .A1(n1612), .A2(n3049), .Y(n2510) );
  OA21X1_LVT U3064 ( .A1(n3480), .A2(n3767), .A3(n8027), .Y(n8030) );
  AND2X1_LVT U3065 ( .A1(n2055), .A2(n2056), .Y(n2096) );
  AND3X1_LVT U3066 ( .A1(n7188), .A2(n7189), .A3(n2622), .Y(n2055) );
  AND4X1_LVT U3067 ( .A1(n7191), .A2(n7193), .A3(n7192), .A4(n2597), .Y(n2056)
         );
  OA21X1_LVT U3068 ( .A1(n3479), .A2(n2120), .A3(n7959), .Y(n7962) );
  AND4X1_LVT U3069 ( .A1(n2057), .A2(n2058), .A3(n2059), .A4(n2060), .Y(n2166)
         );
  AND2X1_LVT U3070 ( .A1(n8136), .A2(n8135), .Y(n2057) );
  AND4X1_LVT U3071 ( .A1(n8150), .A2(n8148), .A3(n8149), .A4(n2614), .Y(n2058)
         );
  AND3X1_LVT U3072 ( .A1(n8134), .A2(n8133), .A3(n8132), .Y(n2059) );
  AND3X1_LVT U3073 ( .A1(n8130), .A2(n8129), .A3(n8128), .Y(n2060) );
  AND3X1_LVT U3074 ( .A1(n2133), .A2(n2574), .A3(n2061), .Y(n2150) );
  AND3X1_LVT U3075 ( .A1(n2062), .A2(n2063), .A3(n2064), .Y(n3740) );
  AND3X1_LVT U3076 ( .A1(n8529), .A2(n8530), .A3(n8531), .Y(n2062) );
  AND2X1_LVT U3077 ( .A1(n8526), .A2(n8525), .Y(n2063) );
  AND3X1_LVT U3078 ( .A1(n8524), .A2(n8523), .A3(n8522), .Y(n2064) );
  NAND3X0_LVT U3079 ( .A1(n2065), .A2(n2066), .A3(n2067), .Y(N691) );
  AND3X1_LVT U3080 ( .A1(n2111), .A2(n2112), .A3(n2113), .Y(n2065) );
  AND3X1_LVT U3081 ( .A1(n7285), .A2(n7284), .A3(n7283), .Y(n2066) );
  AND3X1_LVT U3082 ( .A1(n7281), .A2(n7280), .A3(n7279), .Y(n2067) );
  AND2X1_LVT U3083 ( .A1(n2143), .A2(n6917), .Y(n2068) );
  NAND3X2_LVT U3084 ( .A1(n6940), .A2(n6972), .A3(n3772), .Y(n2069) );
  NAND2X4_LVT U3085 ( .A1(n5446), .A2(n5451), .Y(n3081) );
  AND2X1_LVT U3086 ( .A1(n2070), .A2(n2071), .Y(n2557) );
  AND3X1_LVT U3087 ( .A1(n8112), .A2(n8111), .A3(n8110), .Y(n2070) );
  AND3X1_LVT U3088 ( .A1(n8116), .A2(n8115), .A3(n8114), .Y(n2071) );
  NBUFFX2_LVT U3089 ( .A(ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n2072) );
  AND2X1_LVT U3090 ( .A1(n2073), .A2(n2074), .Y(n2109) );
  AND3X1_LVT U3091 ( .A1(n8168), .A2(n8167), .A3(n8166), .Y(n2073) );
  AND3X1_LVT U3092 ( .A1(n8164), .A2(n8163), .A3(n8162), .Y(n2074) );
  AND2X1_LVT U3093 ( .A1(n2075), .A2(n2076), .Y(n2095) );
  AND4X1_LVT U3094 ( .A1(n7174), .A2(n7172), .A3(n7173), .A4(n2586), .Y(n2075)
         );
  AND3X1_LVT U3095 ( .A1(n7187), .A2(n7186), .A3(n7185), .Y(n2076) );
  AND2X1_LVT U3096 ( .A1(n2077), .A2(n2078), .Y(n3742) );
  AND3X1_LVT U3097 ( .A1(n8452), .A2(n8450), .A3(n2579), .Y(n2077) );
  AND3X1_LVT U3098 ( .A1(n8449), .A2(n8448), .A3(n8447), .Y(n2078) );
  AND2X1_LVT U3099 ( .A1(n2079), .A2(n2080), .Y(n3739) );
  AND3X1_LVT U3100 ( .A1(n8516), .A2(n8514), .A3(n2580), .Y(n2079) );
  AND3X1_LVT U3101 ( .A1(n8513), .A2(n8512), .A3(n8511), .Y(n2080) );
  DELLN1X2_LVT U3102 ( .A(n8105), .Y(n2135) );
  NAND4X1_LVT U3103 ( .A1(n4954), .A2(n4955), .A3(n4953), .A4(n4952), .Y(n9282) );
  AND3X2_LVT U3104 ( .A1(n6940), .A2(n6972), .A3(n3772), .Y(n3689) );
  IBUFFX2_LVT U3105 ( .A(n3768), .Y(n2081) );
  AND2X1_LVT U3106 ( .A1(n2082), .A2(n2083), .Y(n3736) );
  AND3X1_LVT U3107 ( .A1(n8619), .A2(n8617), .A3(n2578), .Y(n2082) );
  AND3X1_LVT U3108 ( .A1(n8616), .A2(n8615), .A3(n8614), .Y(n2083) );
  AND2X1_LVT U3109 ( .A1(n2084), .A2(n2085), .Y(n2159) );
  AND3X1_LVT U3110 ( .A1(n8373), .A2(n8372), .A3(n8371), .Y(n2084) );
  AND3X1_LVT U3111 ( .A1(n8377), .A2(n8376), .A3(n8375), .Y(n2085) );
  OA21X2_LVT U3112 ( .A1(n2657), .A2(n2637), .A3(n2633), .Y(n2130) );
  AND3X1_LVT U3113 ( .A1(n7427), .A2(n7425), .A3(n2610), .Y(n2086) );
  AND3X1_LVT U3114 ( .A1(n7429), .A2(n7428), .A3(n3568), .Y(n2087) );
  AND3X1_LVT U3115 ( .A1(n7442), .A2(n7441), .A3(n7440), .Y(n2088) );
  IBUFFX2_LVT U3116 ( .A(n9036), .Y(n2089) );
  IBUFFX2_LVT U3117 ( .A(n9036), .Y(n2090) );
  AND2X4_LVT U3118 ( .A1(n6939), .A2(n6938), .Y(n9036) );
  NBUFFX2_LVT U3119 ( .A(n9016), .Y(n2091) );
  NBUFFX2_LVT U3120 ( .A(n9016), .Y(n2092) );
  NBUFFX2_LVT U3121 ( .A(n3613), .Y(n3610) );
  NBUFFX2_LVT U3122 ( .A(n9015), .Y(n2093) );
  NBUFFX2_LVT U3123 ( .A(n9015), .Y(n2094) );
  NAND3X0_LVT U3124 ( .A1(n2095), .A2(n2096), .A3(n2097), .Y(N687) );
  AND3X1_LVT U3125 ( .A1(n7171), .A2(n7170), .A3(n7169), .Y(n2097) );
  NBUFFX2_LVT U3126 ( .A(ibuf_io_inst_0_bits_inst_rs1[0]), .Y(n2098) );
  AND3X2_LVT U3127 ( .A1(n6940), .A2(n6926), .A3(n2983), .Y(n9016) );
  NAND3X0_LVT U3128 ( .A1(n2099), .A2(n2100), .A3(n2101), .Y(N726) );
  AND3X1_LVT U3129 ( .A1(n2124), .A2(n2125), .A3(n2126), .Y(n2099) );
  AND3X1_LVT U3130 ( .A1(n8408), .A2(n8407), .A3(n8406), .Y(n2100) );
  AND3X1_LVT U3131 ( .A1(n2117), .A2(n2118), .A3(n2119), .Y(n2101) );
  NAND3X0_LVT U3132 ( .A1(n2102), .A2(n2103), .A3(n2104), .Y(N742) );
  AND3X1_LVT U3133 ( .A1(n2114), .A2(n2115), .A3(n2116), .Y(n2102) );
  AND3X1_LVT U3134 ( .A1(n8974), .A2(n8973), .A3(n8972), .Y(n2103) );
  AND3X1_LVT U3135 ( .A1(n2162), .A2(n2163), .A3(n2164), .Y(n2104) );
  NAND3X0_LVT U3136 ( .A1(n2107), .A2(n2106), .A3(n2105), .Y(n2140) );
  AND2X1_LVT U3137 ( .A1(n3569), .A2(n2142), .Y(n2105) );
  AND4X1_LVT U3138 ( .A1(n7670), .A2(n7683), .A3(n7669), .A4(n2141), .Y(n2106)
         );
  AND3X1_LVT U3139 ( .A1(n7668), .A2(n2592), .A3(n7672), .Y(n2107) );
  AND3X2_LVT U3140 ( .A1(n3773), .A2(n6957), .A3(n6973), .Y(n3712) );
  AND3X2_LVT U3141 ( .A1(n6973), .A2(n6946), .A3(n2983), .Y(n9007) );
  AND3X2_LVT U3142 ( .A1(n6973), .A2(n6974), .A3(n3772), .Y(n2984) );
  AND2X4_LVT U3143 ( .A1(n2144), .A2(n6924), .Y(n6973) );
  NBUFFX2_LVT U3144 ( .A(n9026), .Y(n3760) );
  NBUFFX2_LVT U3145 ( .A(n9026), .Y(n3761) );
  AND3X2_LVT U3146 ( .A1(n6973), .A2(n6957), .A3(n2983), .Y(n9026) );
  NAND3X0_LVT U3147 ( .A1(n2108), .A2(n2109), .A3(n2110), .Y(N719) );
  AND3X1_LVT U3148 ( .A1(n8160), .A2(n8159), .A3(n8158), .Y(n2110) );
  AND3X1_LVT U3149 ( .A1(n7301), .A2(n7300), .A3(n7299), .Y(n2111) );
  AND4X1_LVT U3150 ( .A1(n2595), .A2(n7302), .A3(n7303), .A4(n7304), .Y(n2112)
         );
  AND3X1_LVT U3151 ( .A1(n7298), .A2(n7297), .A3(n7296), .Y(n2113) );
  AND3X1_LVT U3152 ( .A1(n8970), .A2(n8969), .A3(n8968), .Y(n2114) );
  AND3X1_LVT U3153 ( .A1(n8978), .A2(n8977), .A3(n8976), .Y(n2115) );
  AND4X1_LVT U3154 ( .A1(n8979), .A2(n2175), .A3(n2176), .A4(n2177), .Y(n2116)
         );
  AND3X1_LVT U3155 ( .A1(n8412), .A2(n8411), .A3(n8410), .Y(n2117) );
  AND3X1_LVT U3156 ( .A1(n8419), .A2(n8417), .A3(n2605), .Y(n2118) );
  AND3X1_LVT U3157 ( .A1(n8416), .A2(n8415), .A3(n8414), .Y(n2119) );
  NBUFFX2_LVT U3158 ( .A(n9006), .Y(n2120) );
  OR2X4_LVT U3159 ( .A1(n3140), .A2(n2120), .Y(n2668) );
  NBUFFX2_LVT U3160 ( .A(n9030), .Y(n3667) );
  NAND3X0_LVT U3161 ( .A1(n2121), .A2(n2122), .A3(n2123), .Y(N733) );
  AND3X1_LVT U3162 ( .A1(n8643), .A2(n8642), .A3(n8641), .Y(n2121) );
  AND4X1_LVT U3163 ( .A1(n3721), .A2(n3722), .A3(n8655), .A4(n8656), .Y(n2122)
         );
  NOR2X0_LVT U3164 ( .A1(n8670), .A2(n8669), .Y(n2123) );
  DELLN1X2_LVT U3165 ( .A(n5119), .Y(n2134) );
  AND3X1_LVT U3166 ( .A1(n8425), .A2(n8426), .A3(n8427), .Y(n2124) );
  AND3X1_LVT U3167 ( .A1(n8432), .A2(n8433), .A3(n8431), .Y(n2125) );
  AND2X1_LVT U3168 ( .A1(n8428), .A2(n8429), .Y(n2126) );
  AND3X1_LVT U3169 ( .A1(n4511), .A2(n4512), .A3(n4513), .Y(n3049) );
  AND3X2_LVT U3170 ( .A1(n2130), .A2(n5166), .A3(n9432), .Y(n2169) );
  OR2X2_LVT U3171 ( .A1(n3322), .A2(n2969), .Y(n2664) );
  OR2X2_LVT U3172 ( .A1(n3370), .A2(n3989), .Y(n2656) );
  NBUFFX2_LVT U3173 ( .A(n9026), .Y(n3758) );
  NBUFFX2_LVT U3174 ( .A(n9026), .Y(n3756) );
  NBUFFX2_LVT U3175 ( .A(n9026), .Y(n3759) );
  NBUFFX2_LVT U3176 ( .A(n9026), .Y(n3757) );
  NAND3X0_LVT U3177 ( .A1(n2127), .A2(n2128), .A3(n2129), .Y(N713) );
  AND3X1_LVT U3178 ( .A1(n7965), .A2(n7964), .A3(n7963), .Y(n2127) );
  AND3X1_LVT U3179 ( .A1(n2963), .A2(n2964), .A3(n2965), .Y(n2128) );
  AND2X4_LVT U3180 ( .A1(n5403), .A2(n5402), .Y(div_io_resp_ready) );
  DELLN2X2_LVT U3181 ( .A(n9381), .Y(n3046) );
  NAND3X2_LVT U3182 ( .A1(n9436), .A2(n2635), .A3(n5154), .Y(n5066) );
  NAND4X1_LVT U3183 ( .A1(n9075), .A2(n5164), .A3(io_fpu_inst[4]), .A4(n9104), 
        .Y(n2632) );
  AND2X4_LVT U3184 ( .A1(io_fpu_inst[5]), .A2(n9522), .Y(n3575) );
  AND3X4_LVT U3185 ( .A1(n3590), .A2(n3577), .A3(io_fpu_inst[6]), .Y(n5102) );
  OR3X2_LVT U3186 ( .A1(io_fpu_inst[23]), .A2(io_fpu_inst[24]), .A3(
        io_fpu_inst[22]), .Y(n5144) );
  IBUFFX2_LVT U3187 ( .A(ibuf_io_inst_0_bits_inst_rs2[4]), .Y(n5434) );
  AO21X2_LVT U3188 ( .A1(n9076), .A2(n3585), .A3(n3584), .Y(n2131) );
  NBUFFX2_LVT U3189 ( .A(n5423), .Y(n2132) );
  NBUFFX2_LVT U3190 ( .A(n9390), .Y(n2133) );
  NOR2X4_LVT U3191 ( .A1(n5306), .A2(n2132), .Y(n5356) );
  IBUFFX2_LVT U3192 ( .A(n9390), .Y(n9392) );
  AND3X2_LVT U3193 ( .A1(n3046), .A2(n2132), .A3(n5427), .Y(n5379) );
  AND2X4_LVT U3194 ( .A1(n5423), .A2(n5306), .Y(n5339) );
  DELLN1X2_LVT U3195 ( .A(n9022), .Y(n3642) );
  OR3X1_LVT U3196 ( .A1(n2461), .A2(n8078), .A3(n8080), .Y(N716) );
  AND3X1_LVT U3197 ( .A1(n7681), .A2(n7671), .A3(n7682), .Y(n2141) );
  AND2X4_LVT U3198 ( .A1(n2981), .A2(n3796), .Y(n6889) );
  AND2X4_LVT U3199 ( .A1(n2981), .A2(n3868), .Y(n6811) );
  AO21X2_LVT U3200 ( .A1(wb_ctrl_wxd), .A2(csr_io_retire), .A3(n9381), .Y(
        n9397) );
  NAND2X2_LVT U3201 ( .A1(n5415), .A2(n5403), .Y(n9381) );
  IBUFFX2_LVT U3202 ( .A(n5119), .Y(n2547) );
  NBUFFX2_LVT U3203 ( .A(n9519), .Y(io_fpu_inst[29]) );
  NBUFFX2_LVT U3204 ( .A(n2546), .Y(n2137) );
  IBUFFX4_LVT U3205 ( .A(n2546), .Y(n2537) );
  NAND2X0_LVT U3206 ( .A1(n9439), .A2(n2137), .Y(n2568) );
  NOR2X1_LVT U3207 ( .A1(n9517), .A2(n9519), .Y(n2546) );
  AO21X2_LVT U3208 ( .A1(io_fpu_inst[28]), .A2(n2138), .A3(n3039), .Y(n4843)
         );
  OR3X1_LVT U3209 ( .A1(n7684), .A2(n2140), .A3(n7685), .Y(N704) );
  OR2X2_LVT U3210 ( .A1(n9028), .A2(n3327), .Y(n2142) );
  AND3X1_LVT U3211 ( .A1(n2137), .A2(n9447), .A3(n2174), .Y(n4502) );
  NBUFFX2_LVT U3212 ( .A(n9029), .Y(n3637) );
  NAND3X2_LVT U3213 ( .A1(n5008), .A2(n5007), .A3(n5006), .Y(n3048) );
  OA21X2_LVT U3214 ( .A1(n9089), .A2(n9288), .A3(n2134), .Y(n5088) );
  NAND3X1_LVT U3215 ( .A1(n9107), .A2(n1891), .A3(io_fpu_inst[14]), .Y(n9088)
         );
  NAND3X1_LVT U3216 ( .A1(n4918), .A2(csr_io_decode_0_fp_csr), .A3(n2134), .Y(
        n4929) );
  NAND3X2_LVT U3217 ( .A1(n9288), .A2(csr_io_decode_0_write_illegal), .A3(
        n5119), .Y(n5120) );
  NAND3X2_LVT U3218 ( .A1(n5154), .A2(n3593), .A3(n9436), .Y(n5069) );
  OR2X4_LVT U3219 ( .A1(io_fpu_inst[14]), .A2(n3593), .Y(n4509) );
  DELLN1X2_LVT U3220 ( .A(n8932), .Y(n2859) );
  AND2X4_LVT U3221 ( .A1(n4749), .A2(n4752), .Y(n6974) );
  OR2X2_LVT U3222 ( .A1(n4752), .A2(n4969), .Y(n6955) );
  NAND2X0_LVT U3223 ( .A1(n2169), .A2(n2170), .Y(n2143) );
  NAND3X2_LVT U3224 ( .A1(n2533), .A2(n2532), .A3(n9388), .Y(n6935) );
  AND2X4_LVT U3225 ( .A1(n6972), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n9037) );
  AND2X4_LVT U3226 ( .A1(n6972), .A2(n6956), .Y(n8932) );
  AO21X2_LVT U3227 ( .A1(n7068), .A2(n7067), .A3(n3612), .Y(n7069) );
  AO21X2_LVT U3228 ( .A1(n7040), .A2(n7039), .A3(n3612), .Y(n7041) );
  AO21X2_LVT U3229 ( .A1(n7097), .A2(n7096), .A3(n3612), .Y(n7098) );
  AO21X2_LVT U3230 ( .A1(n6968), .A2(n6967), .A3(n3612), .Y(n6969) );
  AO21X2_LVT U3231 ( .A1(n7008), .A2(n7007), .A3(n3612), .Y(n7009) );
  NOR2X4_LVT U3232 ( .A1(n4040), .A2(n3612), .Y(n8939) );
  NOR2X4_LVT U3233 ( .A1(n3184), .A2(n9047), .Y(n8873) );
  NAND2X0_LVT U3234 ( .A1(n2145), .A2(n2146), .Y(n4511) );
  NOR3X4_LVT U3235 ( .A1(n2552), .A2(n4509), .A3(n4508), .Y(n2146) );
  NAND3X1_LVT U3236 ( .A1(n2677), .A2(n1863), .A3(io_fpu_inst[3]), .Y(n_GEN_9)
         );
  OA21X2_LVT U3237 ( .A1(n9438), .A2(n5129), .A3(n3076), .Y(n5068) );
  OR3X1_LVT U3238 ( .A1(n2147), .A2(n2148), .A3(n2149), .Y(n8849) );
  AND2X1_LVT U3239 ( .A1(n_T_427[186]), .A2(n3791), .Y(n2148) );
  DELLN1X2_LVT U3240 ( .A(n9056), .Y(n3600) );
  NBUFFX2_LVT U3241 ( .A(n9517), .Y(io_fpu_inst[31]) );
  AND3X4_LVT U3242 ( .A1(n9412), .A2(n9448), .A3(n9242), .Y(n9116) );
  NAND3X2_LVT U3243 ( .A1(n9412), .A2(n9099), .A3(n5167), .Y(n1431) );
  IBUFFX2_LVT U3244 ( .A(n3040), .Y(n2152) );
  AND2X1_LVT U3245 ( .A1(io_dmem_resp_valid), .A2(io_dmem_resp_bits_has_data), 
        .Y(n2153) );
  NOR2X4_LVT U3246 ( .A1(n9412), .A2(ibuf_io_inst_0_bits_rvc), .Y(n2529) );
  AND2X2_LVT U3247 ( .A1(n6939), .A2(n6936), .Y(n9412) );
  IBUFFX2_LVT U3248 ( .A(n3683), .Y(n2154) );
  IBUFFX2_LVT U3249 ( .A(n3683), .Y(n2155) );
  OA21X2_LVT U3250 ( .A1(n3407), .A2(n3691), .A3(n8561), .Y(n2603) );
  OA21X2_LVT U3251 ( .A1(n3405), .A2(n3708), .A3(n8323), .Y(n8326) );
  NAND3X0_LVT U3252 ( .A1(n2156), .A2(n2157), .A3(n2158), .Y(n8776) );
  AND3X1_LVT U3253 ( .A1(n8753), .A2(n8752), .A3(n2591), .Y(n2156) );
  AND4X1_LVT U3254 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n2638), .Y(n2157)
         );
  AND2X1_LVT U3255 ( .A1(n8755), .A2(n8754), .Y(n2158) );
  AO21X2_LVT U3256 ( .A1(n7588), .A2(n7587), .A3(n9047), .Y(n7589) );
  AO21X2_LVT U3257 ( .A1(n7467), .A2(n7466), .A3(n3631), .Y(n7468) );
  OR2X4_LVT U3258 ( .A1(n8457), .A2(n3612), .Y(n8458) );
  NAND3X0_LVT U3259 ( .A1(n2159), .A2(n2160), .A3(n2161), .Y(N725) );
  NOR3X0_LVT U3260 ( .A1(n8400), .A2(n8399), .A3(n8398), .Y(n2161) );
  AND3X1_LVT U3261 ( .A1(n8990), .A2(n8989), .A3(n8988), .Y(n2162) );
  AND2X1_LVT U3262 ( .A1(n8993), .A2(n8992), .Y(n2163) );
  AND3X1_LVT U3263 ( .A1(n8999), .A2(n8998), .A3(n8997), .Y(n2164) );
  AND3X1_LVT U3264 ( .A1(n8147), .A2(n8146), .A3(n8145), .Y(n2165) );
  AND3X1_LVT U3265 ( .A1(n8266), .A2(n8265), .A3(n8264), .Y(n2167) );
  NOR2X0_LVT U3266 ( .A1(n8276), .A2(n8275), .Y(n2168) );
  NAND2X0_LVT U3267 ( .A1(n2169), .A2(n2170), .Y(n6966) );
  AND3X2_LVT U3268 ( .A1(n5163), .A2(n9434), .A3(n2615), .Y(n5156) );
  NAND3X0_LVT U3269 ( .A1(n2171), .A2(n2172), .A3(n2173), .Y(N730) );
  AND3X1_LVT U3270 ( .A1(n8539), .A2(n8538), .A3(n8537), .Y(n2171) );
  AND3X1_LVT U3271 ( .A1(n8552), .A2(n8551), .A3(n8550), .Y(n2172) );
  NAND3X1_LVT U3272 ( .A1(n2553), .A2(n3079), .A3(n9434), .Y(n5114) );
  IBUFFX2_LVT U3273 ( .A(n9075), .Y(n2639) );
  AND2X1_LVT U3274 ( .A1(n2621), .A2(n6964), .Y(n2561) );
  OR3X1_LVT U3275 ( .A1(n9529), .A2(n9440), .A3(io_fpu_inst[27]), .Y(n4501) );
  OA21X1_LVT U3276 ( .A1(n3148), .A2(n3989), .A3(n8242), .Y(n8245) );
  NAND2X0_LVT U3277 ( .A1(n2527), .A2(n_T_427[447]), .Y(n2619) );
  IBUFFX2_LVT U3278 ( .A(n3715), .Y(n3994) );
  IBUFFX2_LVT U3279 ( .A(n5163), .Y(n9090) );
  OA21X1_LVT U3280 ( .A1(n3170), .A2(n2969), .A3(n9005), .Y(n9011) );
  NAND2X0_LVT U3281 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[17]), .Y(n7470)
         );
  OA21X1_LVT U3282 ( .A1(n3159), .A2(n2969), .A3(n8675), .Y(n8678) );
  NBUFFX2_LVT U3283 ( .A(n9523), .Y(io_fpu_inst[14]) );
  INVX1_LVT U3284 ( .A(n9516), .Y(io_ptw_status_debug) );
  OR2X1_LVT U3285 ( .A1(n9111), .A2(n9445), .Y(n9112) );
  IBUFFX2_LVT U3286 ( .A(io_fpu_inst[8]), .Y(n2174) );
  NAND2X0_LVT U3287 ( .A1(n_T_427[1149]), .A2(n3670), .Y(n2175) );
  OR2X1_LVT U3288 ( .A1(n4011), .A2(n3307), .Y(n2176) );
  NAND2X0_LVT U3289 ( .A1(n_T_427[1277]), .A2(n3641), .Y(n2177) );
  AO22X1_LVT U3290 ( .A1(io_fpu_dmem_resp_data[4]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[4]), .A4(n9065), .Y(n2178) );
  AO22X1_LVT U3291 ( .A1(n_T_628[4]), .A2(n2497), .A3(n_T_918[4]), .A4(n9066), 
        .Y(n2179) );
  OR2X1_LVT U3292 ( .A1(n2178), .A2(n2179), .Y(io_fpu_fromint_data[4]) );
  INVX0_LVT U3293 ( .A(n9492), .Y(n2180) );
  AO222X1_LVT U3294 ( .A1(n2180), .A2(n4060), .A3(n4063), .A4(csr_io_pc[30]), 
        .A5(csr_io_evec[30]), .A6(n4066), .Y(io_imem_req_bits_pc[30]) );
  AND4X1_LVT U3295 ( .A1(n3122), .A2(n3245), .A3(io_dmem_req_bits_cmd[1]), 
        .A4(io_dmem_req_bits_cmd[0]), .Y(n2181) );
  AO21X1_LVT U3296 ( .A1(io_dmem_req_bits_cmd[2]), .A2(n2181), .A3(n2515), .Y(
        n2516) );
  AND2X1_LVT U3297 ( .A1(n2572), .A2(n_T_1187[21]), .Y(n2182) );
  NAND2X0_LVT U3298 ( .A1(n5328), .A2(n5385), .Y(n2183) );
  AO22X1_LVT U3299 ( .A1(n5383), .A2(n5325), .A3(n2182), .A4(n2183), .Y(N767)
         );
  NAND4X0_LVT U3300 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .Y(n2184) );
  AO22X1_LVT U3301 ( .A1(n6813), .A2(n_T_427[832]), .A3(n_T_427[768]), .A4(
        n3906), .Y(n2185) );
  OA22X1_LVT U3302 ( .A1(n3081), .A2(n3138), .A3(n3530), .A4(n3880), .Y(n2186)
         );
  NAND2X0_LVT U3303 ( .A1(n4321), .A2(n3958), .Y(n2187) );
  NAND2X0_LVT U3304 ( .A1(n5479), .A2(n1992), .Y(n2188) );
  NAND4X0_LVT U3305 ( .A1(n2186), .A2(n9382), .A3(n2187), .A4(n2188), .Y(n2189) );
  OR3X1_LVT U3306 ( .A1(n2184), .A2(n2185), .A3(n2189), .Y(n2190) );
  NAND4X0_LVT U3307 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .Y(n2191) );
  INVX0_LVT U3308 ( .A(n5480), .Y(n2192) );
  OA21X1_LVT U3309 ( .A1(n2190), .A2(n2191), .A3(n2192), .Y(N679) );
  AOI22X1_LVT U3310 ( .A1(n_T_918[48]), .A2(n6855), .A3(io_fpu_toint_data[48]), 
        .A4(n6856), .Y(n2193) );
  NAND2X0_LVT U3311 ( .A1(n6857), .A2(n2193), .Y(N646) );
  INVX0_LVT U3312 ( .A(n9356), .Y(n2194) );
  INVX0_LVT U3313 ( .A(n123), .Y(n2195) );
  OA22X1_LVT U3314 ( .A1(n_T_698[18]), .A2(n9496), .A3(n_T_698[12]), .A4(n9491), .Y(n2196) );
  NAND2X0_LVT U3315 ( .A1(n9451), .A2(n9450), .Y(n2197) );
  NAND4X0_LVT U3316 ( .A1(n9453), .A2(n9471), .A3(n9472), .A4(n9452), .Y(n2198) );
  NOR4X0_LVT U3317 ( .A1(n_T_698[0]), .A2(n4599), .A3(n2197), .A4(n2198), .Y(
        n2199) );
  HADDX1_LVT U3318 ( .A0(n9334), .B0(n137), .SO(n2200) );
  OA21X1_LVT U3320 ( .A1(n_T_698[3]), .A2(n9503), .A3(n2202), .Y(n2203) );
  OA21X1_LVT U3321 ( .A1(n9495), .A2(n_T_698[4]), .A3(n2203), .Y(n2204) );
  OA21X1_LVT U3322 ( .A1(n9499), .A2(n_T_698[7]), .A3(n2204), .Y(n2205) );
  OA21X1_LVT U3323 ( .A1(n_T_698[6]), .A2(n9485), .A3(n2205), .Y(n2206) );
  OA21X1_LVT U3324 ( .A1(n_T_698[9]), .A2(n9507), .A3(n2206), .Y(n2207) );
  OA21X1_LVT U3325 ( .A1(n_T_698[8]), .A2(n9511), .A3(n2207), .Y(n2208) );
  OA22X1_LVT U3326 ( .A1(n_T_698[10]), .A2(n9509), .A3(n_T_698[14]), .A4(n9506), .Y(n2209) );
  OA221X1_LVT U3327 ( .A1(n9356), .A2(n123), .A3(n2194), .A4(n2195), .A5(n2211), .Y(n4600) );
  AO22X1_LVT U3328 ( .A1(io_fpu_dmem_resp_data[5]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[5]), .A4(n9065), .Y(n2212) );
  AO22X1_LVT U3329 ( .A1(n_T_628[5]), .A2(n2493), .A3(n_T_918[5]), .A4(n9066), 
        .Y(n2213) );
  OR2X1_LVT U3330 ( .A1(n2212), .A2(n2213), .Y(io_fpu_fromint_data[5]) );
  AO222X1_LVT U3331 ( .A1(n4065), .A2(csr_io_evec[39]), .A3(n9377), .A4(n4059), 
        .A5(n4062), .A6(csr_io_pc[39]), .Y(io_imem_req_bits_pc[39]) );
  NAND2X0_LVT U3332 ( .A1(n5357), .A2(n5356), .Y(n2214) );
  AND2X1_LVT U3333 ( .A1(n_T_1187[2]), .A2(n2214), .Y(n2215) );
  AO22X1_LVT U3334 ( .A1(n2572), .A2(n2215), .A3(n5355), .A4(n5374), .Y(N748)
         );
  AND4X1_LVT U3335 ( .A1(n2973), .A2(n7201), .A3(n7199), .A4(n7200), .Y(n2216)
         );
  AND4X1_LVT U3336 ( .A1(n7216), .A2(n7217), .A3(n7195), .A4(n7196), .Y(n2217)
         );
  AND3X1_LVT U3337 ( .A1(n7218), .A2(n7197), .A3(n2217), .Y(n2218) );
  NAND3X0_LVT U3338 ( .A1(n2974), .A2(n2216), .A3(n2218), .Y(N688) );
  AO222X1_LVT U3339 ( .A1(n9293), .A2(n2515), .A3(n_T_702[24]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[56]), .Y(N517) );
  AO22X1_LVT U3340 ( .A1(n2872), .A2(n_T_427[68]), .A3(n_T_427[1027]), .A4(
        n3900), .Y(n2219) );
  AO22X1_LVT U3341 ( .A1(n2865), .A2(n_T_427[388]), .A3(n_T_427[771]), .A4(
        n3907), .Y(n2220) );
  AO22X1_LVT U3342 ( .A1(n3909), .A2(n_T_427[132]), .A3(n_T_427[452]), .A4(
        n3912), .Y(n2221) );
  AO22X1_LVT U3343 ( .A1(n2879), .A2(n_T_427[4]), .A3(n_T_427[516]), .A4(n2851), .Y(n2222) );
  NOR4X0_LVT U3344 ( .A1(n2219), .A2(n2220), .A3(n2221), .A4(n2222), .Y(n2223)
         );
  AO22X1_LVT U3345 ( .A1(n3917), .A2(n_T_427[1347]), .A3(n_T_427[1475]), .A4(
        n3923), .Y(n2224) );
  AO22X1_LVT U3346 ( .A1(n3927), .A2(n_T_427[1283]), .A3(n_T_427[1411]), .A4(
        n3933), .Y(n2225) );
  AO22X1_LVT U3347 ( .A1(n3937), .A2(n_T_427[1219]), .A3(n_T_427[1155]), .A4(
        n3943), .Y(n2226) );
  AO22X1_LVT U3348 ( .A1(n3947), .A2(n_T_427[963]), .A3(n_T_427[1091]), .A4(
        n3953), .Y(n2227) );
  NOR4X0_LVT U3349 ( .A1(n2224), .A2(n2225), .A3(n2226), .A4(n2227), .Y(n2228)
         );
  NAND2X0_LVT U3350 ( .A1(n4330), .A2(n3958), .Y(n2230) );
  NAND4X0_LVT U3351 ( .A1(n2223), .A2(n2228), .A3(n2229), .A4(n2230), .Y(
        id_rs_1[4]) );
  AOI22X1_LVT U3352 ( .A1(n_T_918[49]), .A2(n6855), .A3(io_fpu_toint_data[49]), 
        .A4(n6856), .Y(n2231) );
  NAND2X0_LVT U3353 ( .A1(n6857), .A2(n2231), .Y(N647) );
  INVX0_LVT U3354 ( .A(n_T_728[0]), .Y(n2232) );
  AOI21X1_LVT U3355 ( .A1(n_T_726[1]), .A2(n2232), .A3(n_T_728[1]), .Y(n2233)
         );
  AO221X1_LVT U3356 ( .A1(n9242), .A2(bpu_io_xcpt_if), .A3(n9242), .A4(n2233), 
        .A5(csr_io_interrupt), .Y(n74) );
  OAI22X1_LVT U3357 ( .A1(n589), .A2(n9163), .A3(n159), .A4(n9164), .Y(n2234)
         );
  NAND3X0_LVT U3358 ( .A1(n9157), .A2(n9155), .A3(n9156), .Y(n2235) );
  OA221X1_LVT U3359 ( .A1(n2235), .A2(io_fpu_dmem_resp_data[3]), .A3(n2235), 
        .A4(n9165), .A5(n9227), .Y(n2236) );
  AO222X1_LVT U3361 ( .A1(n4061), .A2(n9373), .A3(n4066), .A4(csr_io_evec[34]), 
        .A5(csr_io_pc[34]), .A6(n4062), .Y(io_imem_req_bits_pc[34]) );
  INVX0_LVT U3362 ( .A(n9230), .Y(n2238) );
  NAND2X0_LVT U3363 ( .A1(n3583), .A2(n5164), .Y(n2239) );
  OA221X1_LVT U3365 ( .A1(n2669), .A2(n5108), .A3(n2669), .A4(n2629), .A5(
        n2241), .Y(n5166) );
  AND2X1_LVT U3366 ( .A1(n_T_1187[24]), .A2(n2572), .Y(n2242) );
  NAND2X0_LVT U3367 ( .A1(n5379), .A2(n5307), .Y(n2243) );
  AO22X1_LVT U3368 ( .A1(n5366), .A2(n5305), .A3(n2242), .A4(n2243), .Y(N770)
         );
  AO222X1_LVT U3369 ( .A1(n_T_702[23]), .A2(n9301), .A3(n_T_702[7]), .A4(n2515), .A5(n4058), .A6(n_T_702[55]), .Y(N516) );
  AO22X1_LVT U3370 ( .A1(n3932), .A2(n_T_427[1445]), .A3(n_T_427[1381]), .A4(
        n3921), .Y(n2244) );
  AO22X1_LVT U3371 ( .A1(n3942), .A2(n_T_427[1189]), .A3(n_T_427[1317]), .A4(
        n3931), .Y(n2245) );
  AO22X1_LVT U3372 ( .A1(n3952), .A2(n_T_427[1125]), .A3(n_T_427[1253]), .A4(
        n3938), .Y(n2246) );
  AO22X1_LVT U3373 ( .A1(n3898), .A2(n_T_427[1061]), .A3(n_T_427[997]), .A4(
        n3948), .Y(n2247) );
  NOR4X0_LVT U3374 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .Y(n2248)
         );
  NOR4X0_LVT U3375 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .Y(n2250)
         );
  NAND3X0_LVT U3376 ( .A1(n2248), .A2(n2249), .A3(n2250), .Y(id_rs_1[38]) );
  AOI22X1_LVT U3377 ( .A1(n_T_918[50]), .A2(n6855), .A3(io_fpu_toint_data[50]), 
        .A4(n6856), .Y(n2251) );
  NAND2X0_LVT U3378 ( .A1(n6857), .A2(n2251), .Y(N648) );
  INVX0_LVT U3379 ( .A(n9448), .Y(n2252) );
  OR3X1_LVT U3380 ( .A1(bpu_io_xcpt_if), .A2(n_T_726[0]), .A3(n_T_728[0]), .Y(
        n2253) );
  OA221X1_LVT U3381 ( .A1(n9448), .A2(csr_io_interrupt_cause[0]), .A3(n2252), 
        .A4(n2253), .A5(n74), .Y(N303) );
  AO22X1_LVT U3382 ( .A1(io_fpu_dmem_resp_data[6]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[6]), .A4(n9065), .Y(n2254) );
  AO22X1_LVT U3383 ( .A1(n_T_628[6]), .A2(n2497), .A3(n_T_918[6]), .A4(n9066), 
        .Y(n2255) );
  OR2X1_LVT U3384 ( .A1(n2254), .A2(n2255), .Y(io_fpu_fromint_data[6]) );
  AO222X1_LVT U3385 ( .A1(n9302), .A2(n2515), .A3(n_T_702[63]), .A4(n4058), 
        .A5(n9301), .A6(n_T_702[31]), .Y(N524) );
  AO22X1_LVT U3386 ( .A1(n3919), .A2(n_T_427[1375]), .A3(n_T_427[1503]), .A4(
        n3924), .Y(n2256) );
  AO22X1_LVT U3387 ( .A1(n3928), .A2(n_T_427[1311]), .A3(n_T_427[1439]), .A4(
        n3934), .Y(n2257) );
  AO22X1_LVT U3388 ( .A1(n3939), .A2(n_T_427[1247]), .A3(n_T_427[1183]), .A4(
        n3944), .Y(n2258) );
  AO22X1_LVT U3389 ( .A1(n3949), .A2(n_T_427[991]), .A3(n_T_427[1119]), .A4(
        n3954), .Y(n2259) );
  NOR4X0_LVT U3390 ( .A1(n2256), .A2(n2257), .A3(n2258), .A4(n2259), .Y(n2260)
         );
  AOI22X1_LVT U3391 ( .A1(n6884), .A2(n_T_427[736]), .A3(n_T_427[96]), .A4(
        n2872), .Y(n2261) );
  AND4X1_LVT U3392 ( .A1(n2261), .A2(n2689), .A3(n2688), .A4(n2687), .Y(n2262)
         );
  AOI22X1_LVT U3393 ( .A1(n3888), .A2(n_T_427[1631]), .A3(n_T_427[1567]), .A4(
        n3894), .Y(n2263) );
  OA22X1_LVT U3394 ( .A1(n3081), .A2(n3143), .A3(n3082), .A4(n3496), .Y(n2264)
         );
  OA22X1_LVT U3395 ( .A1(n3878), .A2(n6110), .A3(n3276), .A4(n3881), .Y(n2265)
         );
  OA22X2_LVT U3396 ( .A1(n3803), .A2(n3144), .A3(n3495), .A4(n3800), .Y(n2266)
         );
  AND4X1_LVT U3397 ( .A1(n2263), .A2(n2264), .A3(n2265), .A4(n2266), .Y(n2267)
         );
  NAND2X0_LVT U3398 ( .A1(n4406), .A2(n3957), .Y(n2268) );
  NAND4X0_LVT U3399 ( .A1(n2260), .A2(n2262), .A3(n2267), .A4(n2268), .Y(
        id_rs_1[32]) );
  AOI22X1_LVT U3400 ( .A1(n_T_918[51]), .A2(n6855), .A3(io_fpu_toint_data[51]), 
        .A4(n6856), .Y(n2269) );
  NAND2X0_LVT U3401 ( .A1(n6857), .A2(n2269), .Y(N649) );
  AOI22X1_LVT U3402 ( .A1(n9500), .A2(ibuf_io_pc[13]), .A3(n9509), .A4(
        ibuf_io_pc[10]), .Y(n2270) );
  OA221X1_LVT U3403 ( .A1(n9500), .A2(ibuf_io_pc[13]), .A3(n9509), .A4(
        ibuf_io_pc[10]), .A5(n2270), .Y(n2271) );
  INVX0_LVT U3404 ( .A(ibuf_io_pc[15]), .Y(n2272) );
  AOI22X1_LVT U3405 ( .A1(n2272), .A2(n9355), .A3(n9490), .A4(ibuf_io_pc[11]), 
        .Y(n2273) );
  OA221X1_LVT U3406 ( .A1(n2272), .A2(n9355), .A3(n9490), .A4(ibuf_io_pc[11]), 
        .A5(n2273), .Y(n2274) );
  AOI22X1_LVT U3407 ( .A1(n9510), .A2(ibuf_io_pc[19]), .A3(n9504), .A4(
        ibuf_io_pc[29]), .Y(n2275) );
  OA221X1_LVT U3408 ( .A1(n9510), .A2(ibuf_io_pc[19]), .A3(n9504), .A4(
        ibuf_io_pc[29]), .A5(n2275), .Y(n2276) );
  INVX0_LVT U3409 ( .A(ibuf_io_pc[21]), .Y(n2277) );
  INVX0_LVT U3410 ( .A(n9361), .Y(n2278) );
  AO22X1_LVT U3411 ( .A1(ibuf_io_pc[21]), .A2(n9361), .A3(n2277), .A4(n2278), 
        .Y(n2279) );
  NAND4X0_LVT U3412 ( .A1(n2271), .A2(n2274), .A3(n2276), .A4(n2279), .Y(n4575) );
  INVX0_LVT U3413 ( .A(n5426), .Y(n2280) );
  AND2X1_LVT U3414 ( .A1(n2280), .A2(n5428), .Y(n5384) );
  AO22X1_LVT U3415 ( .A1(io_fpu_dmem_resp_data[8]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[8]), .A4(n9065), .Y(n2281) );
  AO22X1_LVT U3416 ( .A1(n_T_628[8]), .A2(n2493), .A3(n_T_918[8]), .A4(n9066), 
        .Y(n2282) );
  OR2X1_LVT U3417 ( .A1(n2281), .A2(n2282), .Y(io_fpu_fromint_data[8]) );
  AO22X1_LVT U3418 ( .A1(io_fpu_dmem_resp_data[16]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[16]), .A4(n9065), .Y(n2283) );
  AO22X1_LVT U3419 ( .A1(n_T_628[16]), .A2(n2497), .A3(n_T_918[16]), .A4(n9066), .Y(n2284) );
  OR2X1_LVT U3420 ( .A1(n2283), .A2(n2284), .Y(io_fpu_fromint_data[16]) );
  AO222X1_LVT U3421 ( .A1(n_T_702[22]), .A2(n9301), .A3(n_T_702[6]), .A4(n2515), .A5(n4058), .A6(n_T_702[54]), .Y(N515) );
  AO22X1_LVT U3422 ( .A1(n3932), .A2(n_T_427[1435]), .A3(n_T_427[1371]), .A4(
        n3921), .Y(n2285) );
  AO22X1_LVT U3423 ( .A1(n3942), .A2(n_T_427[1179]), .A3(n_T_427[1307]), .A4(
        n3931), .Y(n2286) );
  AO22X1_LVT U3424 ( .A1(n3952), .A2(n_T_427[1115]), .A3(n_T_427[1243]), .A4(
        n3941), .Y(n2287) );
  AO22X1_LVT U3425 ( .A1(n3898), .A2(n_T_427[1051]), .A3(n_T_427[987]), .A4(
        n3951), .Y(n2288) );
  NOR4X0_LVT U3426 ( .A1(n2285), .A2(n2286), .A3(n2287), .A4(n2288), .Y(n2289)
         );
  NOR4X0_LVT U3427 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .Y(n2291)
         );
  NAND3X0_LVT U3428 ( .A1(n2289), .A2(n2290), .A3(n2291), .Y(id_rs_1[28]) );
  AOI22X1_LVT U3429 ( .A1(n_T_918[52]), .A2(n6855), .A3(io_fpu_toint_data[52]), 
        .A4(n6856), .Y(n2292) );
  NAND2X0_LVT U3430 ( .A1(n6857), .A2(n2292), .Y(N650) );
  AO22X1_LVT U3431 ( .A1(n9510), .A2(n_T_698[19]), .A3(n9501), .A4(n_T_698[22]), .Y(n2293) );
  AO22X1_LVT U3432 ( .A1(n9488), .A2(n_T_698[23]), .A3(n9497), .A4(n_T_698[25]), .Y(n2294) );
  AO22X1_LVT U3433 ( .A1(n9499), .A2(n_T_698[7]), .A3(n9502), .A4(n_T_698[31]), 
        .Y(n2295) );
  AO22X1_LVT U3434 ( .A1(n9512), .A2(n_T_698[1]), .A3(n9495), .A4(n_T_698[4]), 
        .Y(n2296) );
  OR4X1_LVT U3435 ( .A1(n2293), .A2(n2294), .A3(n2295), .A4(n2296), .Y(n4599)
         );
  INVX0_LVT U3436 ( .A(n5423), .Y(n2297) );
  AND2X1_LVT U3437 ( .A1(n2297), .A2(n5306), .Y(n5335) );
  AO22X1_LVT U3438 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[11]), .A3(
        n_T_918[11]), .A4(n6899), .Y(n2298) );
  AO22X1_LVT U3439 ( .A1(n_T_635[11]), .A2(n6901), .A3(
        io_imem_sfence_bits_addr[11]), .A4(n6900), .Y(n2299) );
  OR2X1_LVT U3440 ( .A1(n2298), .A2(n2299), .Y(n_T_702[11]) );
  AO22X1_LVT U3441 ( .A1(io_fpu_dmem_resp_data[9]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[9]), .A4(n9065), .Y(n2300) );
  AO22X1_LVT U3442 ( .A1(n_T_628[9]), .A2(n2497), .A3(n_T_918[9]), .A4(n9066), 
        .Y(n2301) );
  OR2X1_LVT U3443 ( .A1(n2300), .A2(n2301), .Y(io_fpu_fromint_data[9]) );
  AO22X1_LVT U3444 ( .A1(io_fpu_dmem_resp_data[17]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[17]), .A4(n9065), .Y(n2302) );
  AO22X1_LVT U3445 ( .A1(n_T_628[17]), .A2(n2497), .A3(n_T_918[17]), .A4(n9066), .Y(n2303) );
  OR2X1_LVT U3446 ( .A1(n2302), .A2(n2303), .Y(io_fpu_fromint_data[17]) );
  NAND2X0_LVT U3447 ( .A1(n_T_427[1626]), .A2(n3648), .Y(n2304) );
  AND3X1_LVT U3448 ( .A1(n2304), .A2(n7761), .A3(n7762), .Y(n2305) );
  AND4X1_LVT U3449 ( .A1(n7759), .A2(n2305), .A3(n7758), .A4(n7757), .Y(n2306)
         );
  NAND4X0_LVT U3450 ( .A1(n3061), .A2(n2306), .A3(n3062), .A4(n3063), .Y(N707)
         );
  AO222X1_LVT U3451 ( .A1(n9300), .A2(n2515), .A3(n_T_702[30]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[62]), .Y(N523) );
  AO22X1_LVT U3452 ( .A1(n2862), .A2(n_T_427[144]), .A3(n_T_427[464]), .A4(
        n2824), .Y(n2307) );
  AO22X1_LVT U3453 ( .A1(n3810), .A2(n_T_427[272]), .A3(n3820), .A4(
        n_T_427[656]), .Y(n2308) );
  AO22X1_LVT U3454 ( .A1(n3835), .A2(n_T_427[400]), .A3(n3898), .A4(
        n_T_427[1039]), .Y(n2309) );
  AO22X1_LVT U3455 ( .A1(n3903), .A2(n_T_427[720]), .A3(n_T_427[783]), .A4(
        n2860), .Y(n2310) );
  NOR4X0_LVT U3456 ( .A1(n2307), .A2(n2308), .A3(n2309), .A4(n2310), .Y(n2311)
         );
  AO22X1_LVT U3457 ( .A1(n3918), .A2(n_T_427[1359]), .A3(n_T_427[1487]), .A4(
        n3923), .Y(n2312) );
  AO22X1_LVT U3458 ( .A1(n3928), .A2(n_T_427[1295]), .A3(n_T_427[1423]), .A4(
        n3933), .Y(n2313) );
  AO22X1_LVT U3459 ( .A1(n3938), .A2(n_T_427[1231]), .A3(n_T_427[1167]), .A4(
        n3943), .Y(n2314) );
  AO22X1_LVT U3460 ( .A1(n3948), .A2(n_T_427[975]), .A3(n_T_427[1103]), .A4(
        n3953), .Y(n2315) );
  NOR4X0_LVT U3461 ( .A1(n2312), .A2(n2313), .A3(n2314), .A4(n2315), .Y(n2316)
         );
  AOI22X1_LVT U3462 ( .A1(n3886), .A2(n_T_427[1615]), .A3(n_T_427[1551]), .A4(
        n3891), .Y(n2317) );
  AOI22X1_LVT U3463 ( .A1(n3826), .A2(n_T_427[1679]), .A3(n_T_427[1806]), .A4(
        n3830), .Y(n2318) );
  AND4X1_LVT U3464 ( .A1(n2317), .A2(n2755), .A3(n2756), .A4(n2318), .Y(n2319)
         );
  NAND2X0_LVT U3465 ( .A1(n4364), .A2(n3957), .Y(n2320) );
  NAND4X0_LVT U3466 ( .A1(n2311), .A2(n2316), .A3(n2319), .A4(n2320), .Y(
        id_rs_1[16]) );
  AOI22X1_LVT U3467 ( .A1(n_T_918[53]), .A2(n6855), .A3(io_fpu_toint_data[53]), 
        .A4(n6856), .Y(n2321) );
  NAND2X0_LVT U3468 ( .A1(n6857), .A2(n2321), .Y(N651) );
  AO22X1_LVT U3469 ( .A1(n_T_427[252]), .A2(n3986), .A3(n_T_427[636]), .A4(
        n4034), .Y(n2322) );
  AO22X1_LVT U3470 ( .A1(n4052), .A2(n_T_427[60]), .A3(n_T_427[188]), .A4(
        n2859), .Y(n2323) );
  AO22X1_LVT U3471 ( .A1(n_T_427[700]), .A2(n4021), .A3(n_T_427[955]), .A4(
        n4023), .Y(n2324) );
  OR3X1_LVT U3472 ( .A1(n2322), .A2(n2323), .A3(n2324), .Y(n8902) );
  AO22X1_LVT U3473 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[27]), .A3(
        n_T_918[27]), .A4(n6899), .Y(n2325) );
  AO22X1_LVT U3474 ( .A1(n_T_635[27]), .A2(n6901), .A3(
        io_imem_sfence_bits_addr[27]), .A4(n6900), .Y(n2326) );
  OR2X1_LVT U3475 ( .A1(n2325), .A2(n2326), .Y(n_T_702[27]) );
  AO22X1_LVT U3476 ( .A1(n4054), .A2(n_T_698[1]), .A3(n9103), .A4(
        io_fpu_fromint_data[1]), .Y(alu_io_in1[1]) );
  AO22X1_LVT U3477 ( .A1(io_fpu_dmem_resp_data[12]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[12]), .A4(n9065), .Y(n2327) );
  AO22X1_LVT U3478 ( .A1(n_T_628[12]), .A2(n2497), .A3(n_T_918[12]), .A4(n9066), .Y(n2328) );
  OR2X1_LVT U3479 ( .A1(n2327), .A2(n2328), .Y(io_fpu_fromint_data[12]) );
  NOR4X0_LVT U3480 ( .A1(n8197), .A2(n8196), .A3(n8206), .A4(n8205), .Y(n2329)
         );
  NAND2X0_LVT U3481 ( .A1(n3746), .A2(n2329), .Y(N720) );
  AND2X1_LVT U3482 ( .A1(n_T_1187[26]), .A2(n2572), .Y(n2330) );
  NAND2X0_LVT U3483 ( .A1(n5356), .A2(n5307), .Y(n2331) );
  AO22X1_LVT U3484 ( .A1(n5374), .A2(n5305), .A3(n2330), .A4(n2331), .Y(N772)
         );
  AO222X1_LVT U3485 ( .A1(n9299), .A2(n2515), .A3(n_T_702[29]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[61]), .Y(N522) );
  AO22X1_LVT U3486 ( .A1(n3923), .A2(n_T_427[1485]), .A3(n_T_427[1357]), .A4(
        n3918), .Y(n2332) );
  AO22X1_LVT U3487 ( .A1(n3933), .A2(n_T_427[1421]), .A3(n_T_427[1293]), .A4(
        n3928), .Y(n2333) );
  AO22X1_LVT U3488 ( .A1(n3943), .A2(n_T_427[1165]), .A3(n_T_427[1229]), .A4(
        n3938), .Y(n2334) );
  AO22X1_LVT U3489 ( .A1(n3953), .A2(n_T_427[1101]), .A3(n_T_427[973]), .A4(
        n3948), .Y(n2335) );
  NOR4X0_LVT U3490 ( .A1(n2332), .A2(n2333), .A3(n2334), .A4(n2335), .Y(n2336)
         );
  NOR4X0_LVT U3491 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .Y(n2338)
         );
  NAND4X0_LVT U3492 ( .A1(n2336), .A2(n2337), .A3(n2819), .A4(n2338), .Y(
        id_rs_1[14]) );
  AOI22X1_LVT U3493 ( .A1(n_T_918[54]), .A2(n6855), .A3(io_fpu_toint_data[54]), 
        .A4(n6856), .Y(n2339) );
  NAND2X0_LVT U3494 ( .A1(n6857), .A2(n2339), .Y(N652) );
  AO22X1_LVT U3495 ( .A1(n_T_427[48]), .A2(n4051), .A3(n_T_427[176]), .A4(
        n2859), .Y(n2340) );
  AO22X1_LVT U3496 ( .A1(n4027), .A2(n_T_427[879]), .A3(n_T_427[624]), .A4(
        n4035), .Y(n2341) );
  AO22X1_LVT U3497 ( .A1(n_T_427[240]), .A2(n3983), .A3(n_T_427[688]), .A4(
        n4022), .Y(n2342) );
  OR3X1_LVT U3498 ( .A1(n2340), .A2(n2341), .A3(n2342), .Y(n8470) );
  AO22X1_LVT U3499 ( .A1(io_fpu_dmem_resp_data[3]), .A2(n9064), .A3(n9065), 
        .A4(io_imem_sfence_bits_addr[3]), .Y(n2343) );
  AO22X1_LVT U3500 ( .A1(n9066), .A2(n_T_918[3]), .A3(n2497), .A4(n_T_628[3]), 
        .Y(n2344) );
  OR2X1_LVT U3501 ( .A1(n2343), .A2(n2344), .Y(io_fpu_fromint_data[3]) );
  INVX0_LVT U3502 ( .A(n9508), .Y(n2345) );
  AO222X1_LVT U3503 ( .A1(n2345), .A2(n4061), .A3(csr_io_evec[36]), .A4(n4067), 
        .A5(csr_io_pc[36]), .A6(n4062), .Y(io_imem_req_bits_pc[36]) );
  INVX0_LVT U3504 ( .A(N290), .Y(n2346) );
  NAND4X0_LVT U3505 ( .A1(n5090), .A2(io_dmem_req_bits_cmd[2]), .A3(n559), 
        .A4(io_dmem_req_bits_cmd[4]), .Y(n2347) );
  NAND3X0_LVT U3506 ( .A1(n9426), .A2(n5091), .A3(mem_reg_sfence), .Y(n2348)
         );
  OA21X1_LVT U3507 ( .A1(n2346), .A2(n2347), .A3(n2348), .Y(n2525) );
  AND2X1_LVT U3508 ( .A1(n_T_1187[25]), .A2(n2572), .Y(n2349) );
  NAND2X0_LVT U3509 ( .A1(n5339), .A2(n5307), .Y(n2350) );
  AO22X1_LVT U3510 ( .A1(n5383), .A2(n5305), .A3(n2349), .A4(n2350), .Y(N771)
         );
  AO22X1_LVT U3511 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[7]), .A3(n_T_918[7]), .A4(n6899), .Y(n2351) );
  AO22X1_LVT U3512 ( .A1(n_T_635[7]), .A2(n6901), .A3(
        io_imem_sfence_bits_addr[7]), .A4(n6900), .Y(n2352) );
  OR2X1_LVT U3513 ( .A1(n2351), .A2(n2352), .Y(n_T_702[7]) );
  AO222X1_LVT U3514 ( .A1(n9298), .A2(n2515), .A3(n_T_702[28]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[60]), .Y(N521) );
  AO222X1_LVT U3515 ( .A1(n6249), .A2(mem_br_target_11_), .A3(n_T_918[11]), 
        .A4(n6855), .A5(io_fpu_toint_data[11]), .A6(n6856), .Y(N609) );
  AOI22X1_LVT U3516 ( .A1(n_T_918[55]), .A2(n6855), .A3(io_fpu_toint_data[55]), 
        .A4(n6856), .Y(n2353) );
  NAND2X0_LVT U3517 ( .A1(n6857), .A2(n2353), .Y(N653) );
  AO22X1_LVT U3518 ( .A1(n_T_427[748]), .A2(n4048), .A3(n_T_427[812]), .A4(
        n3982), .Y(n2354) );
  NOR4X0_LVT U3519 ( .A1(n8387), .A2(n8386), .A3(n8385), .A4(n2354), .Y(n2355)
         );
  OR2X1_LVT U3520 ( .A1(n3656), .A2(n2355), .Y(n8388) );
  AO222X1_LVT U3521 ( .A1(n3852), .A2(io_dmem_resp_bits_data[22]), .A3(
        div_io_resp_bits_data[22]), .A4(n3855), .A5(n3849), .A6(
        io_imem_sfence_bits_addr[22]), .Y(n2356) );
  AOI21X1_LVT U3522 ( .A1(csr_io_rw_rdata[22]), .A2(n3844), .A3(n2356), .Y(
        n3094) );
  AOI22X1_LVT U3523 ( .A1(n3910), .A2(n_T_427[448]), .A3(n_T_427[320]), .A4(
        n1918), .Y(n2357) );
  AOI22X1_LVT U3524 ( .A1(n6830), .A2(n_T_427[384]), .A3(n_T_427[767]), .A4(
        n3906), .Y(n2358) );
  AND4X1_LVT U3525 ( .A1(n2357), .A2(n2358), .A3(n2881), .A4(n2880), .Y(n5464)
         );
  AO22X1_LVT U3526 ( .A1(io_fpu_dmem_resp_data[2]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[2]), .A4(n9065), .Y(n2359) );
  AO22X1_LVT U3527 ( .A1(n_T_628[2]), .A2(n2493), .A3(n_T_918[2]), .A4(n9066), 
        .Y(n2360) );
  OR2X1_LVT U3528 ( .A1(n2359), .A2(n2360), .Y(io_fpu_fromint_data[2]) );
  AO22X1_LVT U3529 ( .A1(io_fpu_dmem_resp_data[19]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[19]), .A4(n9065), .Y(n2361) );
  AO22X1_LVT U3530 ( .A1(n_T_628[19]), .A2(n2497), .A3(n_T_918[19]), .A4(n9066), .Y(n2362) );
  OR2X1_LVT U3531 ( .A1(n2361), .A2(n2362), .Y(io_fpu_fromint_data[19]) );
  AO22X1_LVT U3532 ( .A1(io_fpu_dmem_resp_data[29]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[29]), .A4(n9065), .Y(n2363) );
  AO22X1_LVT U3533 ( .A1(n_T_628[29]), .A2(n2497), .A3(n_T_918[29]), .A4(n9066), .Y(n2364) );
  OR2X1_LVT U3534 ( .A1(n2363), .A2(n2364), .Y(io_fpu_fromint_data[29]) );
  NAND2X0_LVT U3535 ( .A1(n3734), .A2(n2365), .Y(N737) );
  AO222X1_LVT U3536 ( .A1(n9297), .A2(n2515), .A3(n_T_702[27]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[59]), .Y(N520) );
  AO222X1_LVT U3537 ( .A1(n6249), .A2(mem_br_target_13_), .A3(n_T_918[13]), 
        .A4(n6855), .A5(io_fpu_toint_data[13]), .A6(n6856), .Y(N611) );
  AOI22X1_LVT U3538 ( .A1(n_T_918[56]), .A2(n6855), .A3(io_fpu_toint_data[56]), 
        .A4(n6856), .Y(n2366) );
  NAND2X0_LVT U3539 ( .A1(n6857), .A2(n2366), .Y(N654) );
  NAND3X0_LVT U3540 ( .A1(n5092), .A2(n5093), .A3(n5094), .Y(n2367) );
  AND2X1_LVT U3541 ( .A1(mem_ctrl_mem), .A2(n2367), .Y(n9424) );
  NOR4X0_LVT U3542 ( .A1(n7680), .A2(n7679), .A3(n7678), .A4(n7677), .Y(n2368)
         );
  NOR4X0_LVT U3543 ( .A1(n7676), .A2(n7675), .A3(n7674), .A4(n7673), .Y(n2369)
         );
  AO21X2_LVT U3544 ( .A1(n2368), .A2(n2369), .A3(n3631), .Y(n7681) );
  HADDX1_LVT U3545 ( .A0(n3104), .B0(n5405), .SO(n2370) );
  NAND2X0_LVT U3546 ( .A1(n2370), .A2(n3251), .Y(n5409) );
  INVX0_LVT U3547 ( .A(ibuf_io_pc[37]), .Y(n2371) );
  INVX0_LVT U3548 ( .A(n9494), .Y(n2372) );
  AO22X1_LVT U3549 ( .A1(ibuf_io_pc[37]), .A2(n9494), .A3(n2371), .A4(n2372), 
        .Y(n4577) );
  AO22X1_LVT U3550 ( .A1(io_fpu_dmem_resp_data[30]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[30]), .A4(n9065), .Y(n2373) );
  AO22X1_LVT U3551 ( .A1(n_T_628[30]), .A2(n2493), .A3(n_T_918[30]), .A4(n9066), .Y(n2374) );
  OR2X1_LVT U3552 ( .A1(n2373), .A2(n2374), .Y(io_fpu_fromint_data[30]) );
  AND2X1_LVT U3553 ( .A1(n_T_1187[28]), .A2(n2572), .Y(n2375) );
  NAND2X0_LVT U3554 ( .A1(n5367), .A2(n5314), .Y(n2376) );
  AO22X1_LVT U3555 ( .A1(n5366), .A2(n5317), .A3(n2375), .A4(n2376), .Y(N774)
         );
  AO222X1_LVT U3556 ( .A1(n_T_702[3]), .A2(n2515), .A3(n_T_702[19]), .A4(n9301), .A5(n4058), .A6(n_T_702[51]), .Y(N512) );
  AO222X1_LVT U3557 ( .A1(mem_br_target_12_), .A2(n6249), .A3(n_T_918[12]), 
        .A4(n6855), .A5(io_fpu_toint_data[12]), .A6(n6856), .Y(N610) );
  AOI22X1_LVT U3558 ( .A1(n_T_918[57]), .A2(n6855), .A3(io_fpu_toint_data[57]), 
        .A4(n6856), .Y(n2377) );
  NAND2X0_LVT U3559 ( .A1(n6857), .A2(n2377), .Y(N655) );
  INVX0_LVT U3560 ( .A(n5095), .Y(n2378) );
  AO221X1_LVT U3561 ( .A1(n5064), .A2(io_dmem_s2_nack), .A3(n5064), .A4(
        blocked), .A5(n2378), .Y(n2379) );
  AND2X1_LVT U3562 ( .A1(n5065), .A2(n2379), .Y(N811) );
  INVX0_LVT U3563 ( .A(n5191), .Y(n2380) );
  NAND3X0_LVT U3564 ( .A1(n5185), .A2(n5184), .A3(n2380), .Y(n5280) );
  INVX0_LVT U3565 ( .A(n5428), .Y(n2381) );
  AND2X1_LVT U3566 ( .A1(n2381), .A2(n5426), .Y(n5328) );
  AO22X1_LVT U3567 ( .A1(n3713), .A2(n_T_427[171]), .A3(n_T_427[555]), .A4(
        n3788), .Y(n8328) );
  AO22X1_LVT U3568 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[16]), .A3(n6899), 
        .A4(n_T_918[16]), .Y(n2382) );
  AO22X1_LVT U3569 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[16]), .A3(n6901), 
        .A4(n_T_635[16]), .Y(n2383) );
  OR2X1_LVT U3570 ( .A1(n2382), .A2(n2383), .Y(n_T_702[16]) );
  AO22X1_LVT U3571 ( .A1(io_fpu_dmem_resp_data[7]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[7]), .A4(n9065), .Y(n2384) );
  AO22X1_LVT U3572 ( .A1(n_T_628[7]), .A2(n2493), .A3(n_T_918[7]), .A4(n9066), 
        .Y(n2385) );
  OR2X1_LVT U3573 ( .A1(n2384), .A2(n2385), .Y(io_fpu_fromint_data[7]) );
  INVX0_LVT U3574 ( .A(io_dmem_s2_nack), .Y(n2386) );
  AND3X1_LVT U3575 ( .A1(wb_reg_valid), .A2(wb_ctrl_fence_i), .A3(n2386), .Y(
        io_imem_flush_icache) );
  NAND2X0_LVT U3576 ( .A1(n_T_427[1630]), .A2(n3652), .Y(n2387) );
  AND3X1_LVT U3577 ( .A1(n2387), .A2(n7881), .A3(n7882), .Y(n2388) );
  AND4X1_LVT U3578 ( .A1(n7879), .A2(n2388), .A3(n7878), .A4(n7877), .Y(n2389)
         );
  NAND4X0_LVT U3579 ( .A1(n3054), .A2(n2389), .A3(n3055), .A4(n3056), .Y(N711)
         );
  AO222X1_LVT U3580 ( .A1(n9296), .A2(n2515), .A3(n_T_702[26]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[58]), .Y(N519) );
  NAND2X0_LVT U3581 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[3]), .Y(n2390) );
  NAND4X0_LVT U3582 ( .A1(n9157), .A2(n9155), .A3(n9156), .A4(n2390), .Y(
        n_T_702[3]) );
  AO222X1_LVT U3583 ( .A1(n6249), .A2(mem_br_target_17_), .A3(n_T_918[17]), 
        .A4(n6855), .A5(io_fpu_toint_data[17]), .A6(n6856), .Y(N615) );
  AOI22X1_LVT U3584 ( .A1(n_T_918[63]), .A2(n6855), .A3(io_fpu_toint_data[63]), 
        .A4(n6856), .Y(n2391) );
  NAND2X0_LVT U3585 ( .A1(n6857), .A2(n2391), .Y(N661) );
  OA221X1_LVT U3586 ( .A1(n5396), .A2(io_fpu_inst[26]), .A3(n5396), .A4(n1847), 
        .A5(n2873), .Y(n2392) );
  INVX0_LVT U3587 ( .A(n5063), .Y(n2393) );
  OA221X1_LVT U3588 ( .A1(n2392), .A2(id_reg_fence), .A3(n2393), .A4(n2392), 
        .A5(n4498), .Y(n1821) );
  INVX0_LVT U3589 ( .A(ibuf_io_pc[30]), .Y(n2394) );
  INVX0_LVT U3590 ( .A(n9492), .Y(n2395) );
  AO22X1_LVT U3591 ( .A1(ibuf_io_pc[30]), .A2(n9492), .A3(n2394), .A4(n2395), 
        .Y(n4587) );
  AOI22X1_LVT U3592 ( .A1(n3745), .A2(n_T_427[246]), .A3(n3771), .A4(
        n_T_427[757]), .Y(n3719) );
  AO22X1_LVT U3593 ( .A1(io_fpu_dmem_resp_data[13]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[13]), .A4(n9065), .Y(n2396) );
  AO22X1_LVT U3594 ( .A1(n_T_628[13]), .A2(n2493), .A3(n_T_918[13]), .A4(n9066), .Y(n2397) );
  OR2X1_LVT U3595 ( .A1(n2396), .A2(n2397), .Y(io_fpu_fromint_data[13]) );
  INVX0_LVT U3596 ( .A(csr_io_interrupt_cause[3]), .Y(n2398) );
  OA21X1_LVT U3597 ( .A1(n9448), .A2(n2398), .A3(n74), .Y(n2507) );
  OA22X1_LVT U3598 ( .A1(n5237), .A2(n5292), .A3(n5295), .A4(n5238), .Y(n2399)
         );
  AO22X1_LVT U3599 ( .A1(n3793), .A2(n_T_1298[11]), .A3(n5298), .A4(n5239), 
        .Y(n2400) );
  AND2X1_LVT U3600 ( .A1(n2399), .A2(n2400), .Y(N790) );
  NAND2X0_LVT U3601 ( .A1(n_T_427[1627]), .A2(n3651), .Y(n2401) );
  AND3X1_LVT U3602 ( .A1(n2401), .A2(n7793), .A3(n7794), .Y(n2402) );
  AND4X1_LVT U3603 ( .A1(n7791), .A2(n2402), .A3(n7790), .A4(n7789), .Y(n2403)
         );
  NAND4X0_LVT U3604 ( .A1(n3051), .A2(n2403), .A3(n3052), .A4(n3053), .Y(N708)
         );
  AO222X1_LVT U3605 ( .A1(n_T_702[4]), .A2(n2515), .A3(n_T_702[20]), .A4(n9301), .A5(n4058), .A6(n_T_702[52]), .Y(N513) );
  AO22X1_LVT U3606 ( .A1(n6813), .A2(n_T_427[842]), .A3(n2826), .A4(
        n_T_427[11]), .Y(n2404) );
  OAI22X1_LVT U3607 ( .A1(n3879), .A2(n5681), .A3(n3186), .A4(n3596), .Y(n2405) );
  NOR4X0_LVT U3608 ( .A1(n5676), .A2(n5675), .A3(n2404), .A4(n2405), .Y(n2406)
         );
  AOI22X1_LVT U3609 ( .A1(n3827), .A2(n_T_427[1674]), .A3(n3890), .A4(
        n_T_427[1546]), .Y(n2407) );
  AOI22X1_LVT U3610 ( .A1(n3922), .A2(n_T_427[1482]), .A3(n_T_427[1610]), .A4(
        n3889), .Y(n2408) );
  AOI22X2_LVT U3611 ( .A1(n3828), .A2(n_T_427[1801]), .A3(n_T_427[1738]), .A4(
        n2866), .Y(n2409) );
  AND4X1_LVT U3612 ( .A1(n2407), .A2(n2750), .A3(n2409), .A4(n2408), .Y(n2410)
         );
  AO22X1_LVT U3613 ( .A1(n3932), .A2(n_T_427[1418]), .A3(n_T_427[1354]), .A4(
        n3921), .Y(n2411) );
  AO22X1_LVT U3614 ( .A1(n3942), .A2(n_T_427[1162]), .A3(n_T_427[1290]), .A4(
        n3931), .Y(n2412) );
  AO22X1_LVT U3615 ( .A1(n3952), .A2(n_T_427[1098]), .A3(n_T_427[1226]), .A4(
        n3941), .Y(n2413) );
  AO22X1_LVT U3616 ( .A1(n3898), .A2(n_T_427[1034]), .A3(n_T_427[970]), .A4(
        n3951), .Y(n2414) );
  NOR4X0_LVT U3617 ( .A1(n2411), .A2(n2412), .A3(n2413), .A4(n2414), .Y(n2415)
         );
  NAND2X0_LVT U3618 ( .A1(n3819), .A2(n_T_427[523]), .Y(n2416) );
  NAND4X0_LVT U3619 ( .A1(n2406), .A2(n2410), .A3(n2415), .A4(n2416), .Y(
        id_rs_1[11]) );
  AO222X1_LVT U3620 ( .A1(n6249), .A2(mem_br_target_19_), .A3(n_T_918[19]), 
        .A4(n6855), .A5(io_fpu_toint_data[19]), .A6(n6856), .Y(N617) );
  AOI22X1_LVT U3621 ( .A1(n_T_918[58]), .A2(n6855), .A3(io_fpu_toint_data[58]), 
        .A4(n6856), .Y(n2417) );
  NAND2X0_LVT U3622 ( .A1(n6857), .A2(n2417), .Y(N656) );
  INVX0_LVT U3623 ( .A(n4507), .Y(n2418) );
  OA22X1_LVT U3624 ( .A1(io_fpu_inst[5]), .A2(n9109), .A3(io_fpu_inst[13]), 
        .A4(n2418), .Y(n2419) );
  AOI22X1_LVT U3625 ( .A1(io_fpu_inst[5]), .A2(n3077), .A3(n2552), .A4(n5067), 
        .Y(n2420) );
  NAND2X0_LVT U3626 ( .A1(n2639), .A2(n5074), .Y(n2421) );
  NAND4X0_LVT U3627 ( .A1(n5174), .A2(n2419), .A3(n2420), .A4(n2421), .Y(
        id_ctrl_wxd) );
  OR4X1_LVT U3628 ( .A1(ex_ctrl_div), .A2(ex_ctrl_csr[0]), .A3(ex_ctrl_csr[2]), 
        .A4(io_dmem_req_bits_tag[0]), .Y(n2422) );
  NOR4X0_LVT U3629 ( .A1(ex_ctrl_mem), .A2(ex_ctrl_jalr), .A3(ex_ctrl_csr[1]), 
        .A4(n2422), .Y(n5051) );
  INVX0_LVT U3630 ( .A(n5191), .Y(n2423) );
  NAND3X0_LVT U3631 ( .A1(n5185), .A2(io_fpu_dmem_resp_tag[0]), .A3(n2423), 
        .Y(n5270) );
  AND3X1_LVT U3632 ( .A1(n5481), .A2(ex_reg_rs_bypass_1), .A3(n5483), .Y(n6899) );
  AO222X1_LVT U3633 ( .A1(n3851), .A2(io_dmem_resp_bits_data[11]), .A3(
        div_io_resp_bits_data[11]), .A4(n3854), .A5(n3850), .A6(
        io_imem_sfence_bits_addr[11]), .Y(n2424) );
  AOI21X1_LVT U3634 ( .A1(csr_io_rw_rdata[11]), .A2(n3842), .A3(n2424), .Y(
        n3186) );
  AO22X1_LVT U3635 ( .A1(io_fpu_dmem_resp_data[15]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[15]), .A4(n9065), .Y(n2425) );
  AO22X1_LVT U3636 ( .A1(n_T_628[15]), .A2(n2493), .A3(n_T_918[15]), .A4(n9066), .Y(n2426) );
  OR2X1_LVT U3637 ( .A1(n2425), .A2(n2426), .Y(io_fpu_fromint_data[15]) );
  AND4X1_LVT U3638 ( .A1(n2927), .A2(n3677), .A3(n2926), .A4(n3676), .Y(n2427)
         );
  NAND3X0_LVT U3639 ( .A1(n3779), .A2(n2427), .A3(n3690), .Y(N715) );
  AO222X1_LVT U3640 ( .A1(n_T_702[2]), .A2(n2515), .A3(n_T_702[18]), .A4(n9301), .A5(n4058), .A6(n_T_702[50]), .Y(N511) );
  AND4X1_LVT U3641 ( .A1(n2841), .A2(n2840), .A3(n2839), .A4(n2838), .Y(n2428)
         );
  AO22X1_LVT U3642 ( .A1(n3928), .A2(n_T_427[1298]), .A3(n_T_427[1426]), .A4(
        n3934), .Y(n2430) );
  AO22X1_LVT U3643 ( .A1(n3938), .A2(n_T_427[1234]), .A3(n_T_427[1170]), .A4(
        n3944), .Y(n2431) );
  AO22X1_LVT U3644 ( .A1(n3948), .A2(n_T_427[978]), .A3(n_T_427[1106]), .A4(
        n3954), .Y(n2432) );
  AO22X1_LVT U3645 ( .A1(n2830), .A2(n_T_427[211]), .A3(n_T_427[1042]), .A4(
        n3900), .Y(n2433) );
  NOR4X0_LVT U3646 ( .A1(n2430), .A2(n2431), .A3(n2432), .A4(n2433), .Y(n2434)
         );
  NAND3X0_LVT U3647 ( .A1(n2428), .A2(n2429), .A3(n2434), .Y(id_rs_1[19]) );
  AO222X1_LVT U3648 ( .A1(n6249), .A2(mem_br_target_14_), .A3(n_T_918[14]), 
        .A4(n6855), .A5(io_fpu_toint_data[14]), .A6(n6856), .Y(N612) );
  AO222X1_LVT U3649 ( .A1(n6249), .A2(mem_br_target_25_), .A3(n_T_918[25]), 
        .A4(n6855), .A5(io_fpu_toint_data[25]), .A6(n6856), .Y(N623) );
  AOI22X1_LVT U3650 ( .A1(n_T_918[59]), .A2(n6855), .A3(io_fpu_toint_data[59]), 
        .A4(n6856), .Y(n2435) );
  NAND2X0_LVT U3651 ( .A1(n6857), .A2(n2435), .Y(N657) );
  AOI21X1_LVT U3652 ( .A1(io_dmem_req_bits_cmd[1]), .A2(n560), .A3(n5078), .Y(
        n2436) );
  OA221X1_LVT U3653 ( .A1(io_dmem_req_bits_cmd[3]), .A2(
        io_dmem_req_bits_cmd[2]), .A3(io_dmem_req_bits_cmd[3]), .A4(n2436), 
        .A5(n3245), .Y(n997) );
  INVX0_LVT U3654 ( .A(n5169), .Y(n2437) );
  AO22X1_LVT U3655 ( .A1(io_imem_req_bits_speculative), .A2(mem_reg_replay), 
        .A3(io_imem_bht_update_valid), .A4(n2437), .Y(N530) );
  INVX0_LVT U3656 ( .A(io_fpu_sboard_clra[3]), .Y(n2438) );
  AND2X1_LVT U3657 ( .A1(n2438), .A2(io_fpu_sboard_clra[4]), .Y(n5258) );
  INVX0_LVT U3658 ( .A(io_fpu_sboard_clra[4]), .Y(n2439) );
  NAND2X0_LVT U3659 ( .A1(io_fpu_sboard_clra[3]), .A2(n2439), .Y(n5245) );
  AO22X1_LVT U3660 ( .A1(io_fpu_dmem_resp_data[10]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[10]), .A4(n9065), .Y(n2440) );
  AO22X1_LVT U3661 ( .A1(n_T_628[10]), .A2(n2497), .A3(n_T_918[10]), .A4(n9066), .Y(n2441) );
  OR2X1_LVT U3662 ( .A1(n2440), .A2(n2441), .Y(io_fpu_fromint_data[10]) );
  NAND2X0_LVT U3663 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[4]), .Y(n2442) );
  NAND4X0_LVT U3664 ( .A1(n9161), .A2(n9159), .A3(n9160), .A4(n2442), .Y(
        n_T_702[4]) );
  AO222X1_LVT U3665 ( .A1(n_T_702[0]), .A2(n2515), .A3(n_T_702[16]), .A4(n9301), .A5(n4058), .A6(n_T_702[48]), .Y(N509) );
  NAND2X0_LVT U3666 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[2]), .Y(n2443) );
  NAND4X0_LVT U3667 ( .A1(n9150), .A2(n9148), .A3(n9149), .A4(n2443), .Y(
        n_T_702[2]) );
  AO22X1_LVT U3668 ( .A1(n3932), .A2(n_T_427[1432]), .A3(n_T_427[1368]), .A4(
        n3921), .Y(n2444) );
  AO22X1_LVT U3669 ( .A1(n3942), .A2(n_T_427[1176]), .A3(n_T_427[1304]), .A4(
        n3931), .Y(n2445) );
  AO22X1_LVT U3670 ( .A1(n3952), .A2(n_T_427[1112]), .A3(n_T_427[1240]), .A4(
        n3941), .Y(n2446) );
  AO22X1_LVT U3671 ( .A1(n3898), .A2(n_T_427[1048]), .A3(n_T_427[984]), .A4(
        n3951), .Y(n2447) );
  NOR4X0_LVT U3672 ( .A1(n2444), .A2(n2445), .A3(n2446), .A4(n2447), .Y(n2448)
         );
  AO22X1_LVT U3673 ( .A1(n3922), .A2(n_T_427[1496]), .A3(n_T_427[1624]), .A4(
        n3889), .Y(n2449) );
  NOR4X0_LVT U3674 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n2449), .Y(n2450)
         );
  NOR4X0_LVT U3675 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .Y(n2451)
         );
  NAND3X0_LVT U3676 ( .A1(n2448), .A2(n2450), .A3(n2451), .Y(id_rs_1[25]) );
  AO222X1_LVT U3677 ( .A1(mem_br_target_8_), .A2(n6249), .A3(n_T_918[8]), .A4(
        n6855), .A5(io_fpu_toint_data[8]), .A6(n6856), .Y(N606) );
  AO222X1_LVT U3678 ( .A1(n6249), .A2(mem_br_target_15_), .A3(n_T_918[15]), 
        .A4(n6855), .A5(io_fpu_toint_data[15]), .A6(n6856), .Y(N613) );
  AO222X1_LVT U3679 ( .A1(mem_br_target_21_), .A2(n6249), .A3(n_T_918[21]), 
        .A4(n6855), .A5(io_fpu_toint_data[21]), .A6(n6856), .Y(N619) );
  AO222X1_LVT U3680 ( .A1(n6249), .A2(mem_br_target_27_), .A3(n_T_918[27]), 
        .A4(n6855), .A5(io_fpu_toint_data[27]), .A6(n6856), .Y(N625) );
  AOI22X1_LVT U3681 ( .A1(n_T_918[60]), .A2(n6855), .A3(io_fpu_toint_data[60]), 
        .A4(n6856), .Y(n2452) );
  NAND2X0_LVT U3682 ( .A1(n6857), .A2(n2452), .Y(N658) );
  OA221X1_LVT U3683 ( .A1(n1853), .A2(n3597), .A3(io_fpu_inst[3]), .A4(n9445), 
        .A5(n9109), .Y(n2453) );
  NOR2X0_LVT U3684 ( .A1(n1431), .A2(n2453), .Y(N275) );
  INVX0_LVT U3685 ( .A(io_imem_req_bits_speculative), .Y(n2454) );
  AOI221X1_LVT U3686 ( .A1(mem_reg_valid), .A2(mem_reg_sfence), .A3(
        mem_reg_valid), .A4(io_imem_bht_update_bits_mispredict), .A5(n2454), 
        .Y(n9418) );
  NAND2X0_LVT U3687 ( .A1(n118), .A2(n9361), .Y(n2455) );
  OA221X1_LVT U3688 ( .A1(n9501), .A2(n_T_698[22]), .A3(n118), .A4(n9361), 
        .A5(n2455), .Y(n4603) );
  INVX0_LVT U3689 ( .A(n5191), .Y(n2456) );
  NAND3X0_LVT U3690 ( .A1(io_fpu_dmem_resp_tag[1]), .A2(n5184), .A3(n2456), 
        .Y(n5261) );
  AO22X1_LVT U3691 ( .A1(io_fpu_dmem_resp_data[14]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[14]), .A4(n9065), .Y(n2457) );
  AO22X1_LVT U3692 ( .A1(n_T_628[14]), .A2(n2497), .A3(n_T_918[14]), .A4(n9066), .Y(n2458) );
  OR2X1_LVT U3693 ( .A1(n2457), .A2(n2458), .Y(io_fpu_fromint_data[14]) );
  AND2X1_LVT U3694 ( .A1(n_T_1187[29]), .A2(n2572), .Y(n2459) );
  NAND2X0_LVT U3695 ( .A1(n5385), .A2(n5314), .Y(n2460) );
  AO22X1_LVT U3696 ( .A1(n5383), .A2(n5317), .A3(n2459), .A4(n2460), .Y(N775)
         );
  OR4X1_LVT U3697 ( .A1(n8059), .A2(n8077), .A3(n8079), .A4(n8060), .Y(n2461)
         );
  AO222X1_LVT U3698 ( .A1(n_T_702[17]), .A2(n9301), .A3(n_T_702[1]), .A4(n2515), .A5(n4058), .A6(n_T_702[49]), .Y(N510) );
  AO222X1_LVT U3699 ( .A1(n6249), .A2(mem_br_target_9_), .A3(n_T_918[9]), .A4(
        n6855), .A5(io_fpu_toint_data[9]), .A6(n6856), .Y(N607) );
  AO222X1_LVT U3700 ( .A1(n6249), .A2(mem_br_target_16_), .A3(n_T_918[16]), 
        .A4(n6855), .A5(io_fpu_toint_data[16]), .A6(n6856), .Y(N614) );
  AO222X1_LVT U3701 ( .A1(n6249), .A2(mem_br_target_23_), .A3(n_T_918[23]), 
        .A4(n6855), .A5(io_fpu_toint_data[23]), .A6(n6856), .Y(N621) );
  AO222X1_LVT U3702 ( .A1(n6249), .A2(mem_br_target_29_), .A3(n_T_918[29]), 
        .A4(n6855), .A5(io_fpu_toint_data[29]), .A6(n6856), .Y(N627) );
  AO222X1_LVT U3703 ( .A1(n6249), .A2(mem_br_target_34_), .A3(n_T_918[34]), 
        .A4(n6855), .A5(io_fpu_toint_data[34]), .A6(n6856), .Y(N632) );
  AOI22X1_LVT U3704 ( .A1(n_T_918[61]), .A2(n6855), .A3(io_fpu_toint_data[61]), 
        .A4(n6856), .Y(n2462) );
  NAND2X0_LVT U3705 ( .A1(n6857), .A2(n2462), .Y(N659) );
  AOI22X1_LVT U3706 ( .A1(n5123), .A2(n5087), .A3(csr_io_decode_0_write_flush), 
        .A4(n5088), .Y(n2463) );
  INVX0_LVT U3707 ( .A(n1828), .Y(n2464) );
  NAND3X0_LVT U3708 ( .A1(n2463), .A2(n5122), .A3(n2464), .Y(n_T_731) );
  INVX0_LVT U3709 ( .A(div_io_req_ready), .Y(n2465) );
  NAND2X0_LVT U3710 ( .A1(n9422), .A2(n2465), .Y(n2466) );
  NAND3X0_LVT U3711 ( .A1(ex_reg_valid), .A2(n5175), .A3(ex_reg_load_use), .Y(
        n2467) );
  AND4X1_LVT U3712 ( .A1(n3233), .A2(n5095), .A3(n2466), .A4(n2467), .Y(n9421)
         );
  OA22X2_LVT U3713 ( .A1(n3803), .A2(n3170), .A3(n3488), .A4(n3800), .Y(n2468)
         );
  OA22X1_LVT U3714 ( .A1(n3082), .A2(n3489), .A3(n3081), .A4(n3171), .Y(n2469)
         );
  AOI22X1_LVT U3715 ( .A1(n3894), .A2(n_T_427[1598]), .A3(n_T_427[1662]), .A4(
        n3889), .Y(n2470) );
  AND4X1_LVT U3716 ( .A1(n2468), .A2(n6881), .A3(n2470), .A4(n2469), .Y(n2471)
         );
  AO22X1_LVT U3717 ( .A1(n3909), .A2(n_T_427[191]), .A3(n3911), .A4(
        n_T_427[511]), .Y(n2472) );
  AO22X1_LVT U3718 ( .A1(n3916), .A2(n_T_427[639]), .A3(n_T_427[63]), .A4(
        n3913), .Y(n2473) );
  AO22X1_LVT U3719 ( .A1(n3899), .A2(n_T_427[1086]), .A3(n_T_427[958]), .A4(
        n2831), .Y(n2474) );
  AO22X1_LVT U3720 ( .A1(n3905), .A2(n_T_427[766]), .A3(n_T_427[830]), .A4(
        n2861), .Y(n2475) );
  NOR4X0_LVT U3721 ( .A1(n2472), .A2(n2473), .A3(n2474), .A4(n2475), .Y(n2476)
         );
  AO22X1_LVT U3722 ( .A1(n3922), .A2(n_T_427[1534]), .A3(n_T_427[1406]), .A4(
        n3917), .Y(n2477) );
  AO22X1_LVT U3723 ( .A1(n3933), .A2(n_T_427[1470]), .A3(n_T_427[1342]), .A4(
        n3927), .Y(n2478) );
  AO22X1_LVT U3724 ( .A1(n3942), .A2(n_T_427[1214]), .A3(n_T_427[1278]), .A4(
        n3937), .Y(n2479) );
  AO22X1_LVT U3725 ( .A1(n3952), .A2(n_T_427[1150]), .A3(n_T_427[1022]), .A4(
        n3947), .Y(n2480) );
  NOR4X0_LVT U3726 ( .A1(n2477), .A2(n2478), .A3(n2479), .A4(n2480), .Y(n2481)
         );
  NAND2X0_LVT U3727 ( .A1(n4496), .A2(n3959), .Y(n2482) );
  NAND4X0_LVT U3728 ( .A1(n2471), .A2(n2476), .A3(n2481), .A4(n2482), .Y(
        id_rs_1[63]) );
  INVX0_LVT U3729 ( .A(io_fpu_sboard_clra[1]), .Y(n2483) );
  AND2X1_LVT U3730 ( .A1(n2483), .A2(io_fpu_sboard_clr), .Y(n5183) );
  NAND2X0_LVT U3731 ( .A1(n_T_427[59]), .A2(n8944), .Y(n2484) );
  NAND3X0_LVT U3732 ( .A1(n2484), .A2(n8887), .A3(n8886), .Y(n2582) );
  OAI21X1_LVT U3733 ( .A1(n2968), .A2(n1262), .A3(n9412), .Y(n9383) );
  INVX0_LVT U3734 ( .A(n5191), .Y(n2485) );
  NAND3X0_LVT U3735 ( .A1(io_fpu_dmem_resp_tag[0]), .A2(
        io_fpu_dmem_resp_tag[1]), .A3(n2485), .Y(n5292) );
  AO22X1_LVT U3736 ( .A1(io_fpu_dmem_resp_data[11]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[11]), .A4(n9065), .Y(n2486) );
  AO22X1_LVT U3737 ( .A1(n_T_628[11]), .A2(n2493), .A3(n_T_918[11]), .A4(n9066), .Y(n2487) );
  OR2X1_LVT U3738 ( .A1(n2486), .A2(n2487), .Y(io_fpu_fromint_data[11]) );
  AND3X1_LVT U3739 ( .A1(n9179), .A2(n9173), .A3(n9200), .Y(n9199) );
  AO222X1_LVT U3740 ( .A1(n_T_702[21]), .A2(n9301), .A3(n_T_702[5]), .A4(n2515), .A5(n4058), .A6(n_T_702[53]), .Y(N514) );
  INVX0_LVT U3741 ( .A(n5483), .Y(n2488) );
  NAND2X0_LVT U3742 ( .A1(io_fpu_dmem_resp_data[1]), .A2(n2488), .Y(n2489) );
  NAND4X0_LVT U3743 ( .A1(n9135), .A2(n9136), .A3(n9137), .A4(n2489), .Y(
        n_T_702[1]) );
  AO222X1_LVT U3744 ( .A1(n6249), .A2(mem_br_target_10_), .A3(n_T_918[10]), 
        .A4(n6855), .A5(io_fpu_toint_data[10]), .A6(n6856), .Y(N608) );
  AO222X1_LVT U3745 ( .A1(n6249), .A2(mem_br_target_18_), .A3(n_T_918[18]), 
        .A4(n6855), .A5(io_fpu_toint_data[18]), .A6(n6856), .Y(N616) );
  AO222X1_LVT U3746 ( .A1(n6249), .A2(mem_br_target_20_), .A3(n_T_918[20]), 
        .A4(n6855), .A5(io_fpu_toint_data[20]), .A6(n6856), .Y(N618) );
  AO222X1_LVT U3747 ( .A1(mem_br_target_22_), .A2(n6249), .A3(n_T_918[22]), 
        .A4(n6855), .A5(io_fpu_toint_data[22]), .A6(n6856), .Y(N620) );
  AO222X1_LVT U3748 ( .A1(n6249), .A2(mem_br_target_24_), .A3(n_T_918[24]), 
        .A4(n6855), .A5(io_fpu_toint_data[24]), .A6(n6856), .Y(N622) );
  AO222X1_LVT U3749 ( .A1(n6249), .A2(mem_br_target_26_), .A3(n_T_918[26]), 
        .A4(n6855), .A5(io_fpu_toint_data[26]), .A6(n6856), .Y(N624) );
  AO222X1_LVT U3750 ( .A1(n6249), .A2(mem_br_target_28_), .A3(n_T_918[28]), 
        .A4(n6855), .A5(io_fpu_toint_data[28]), .A6(n6856), .Y(N626) );
  AO222X1_LVT U3751 ( .A1(n6249), .A2(mem_br_target_30_), .A3(n_T_918[30]), 
        .A4(n6855), .A5(io_fpu_toint_data[30]), .A6(n6856), .Y(N628) );
  AO222X1_LVT U3752 ( .A1(n6249), .A2(mem_br_target_36_), .A3(n_T_918[36]), 
        .A4(n6855), .A5(io_fpu_toint_data[36]), .A6(n6856), .Y(N634) );
  AO222X1_LVT U3753 ( .A1(n6249), .A2(mem_br_target_37_), .A3(n_T_918[37]), 
        .A4(n6855), .A5(io_fpu_toint_data[37]), .A6(n6856), .Y(N635) );
  AOI22X1_LVT U3754 ( .A1(n_T_918[62]), .A2(n6855), .A3(io_fpu_toint_data[62]), 
        .A4(n6856), .Y(n2490) );
  NAND2X0_LVT U3755 ( .A1(n6857), .A2(n2490), .Y(N660) );
  AO221X1_LVT U3756 ( .A1(n1853), .A2(io_fpu_inst[31]), .A3(n1853), .A4(n5099), 
        .A5(io_fpu_inst[6]), .Y(id_ctrl_mem_cmd_2_) );
  IBUFFX2_LVT U3757 ( .A(n3081), .Y(n2765) );
  IBUFFX2_LVT U3758 ( .A(n3081), .Y(n3830) );
  IBUFFX2_LVT U3759 ( .A(n3081), .Y(n3828) );
  IBUFFX2_LVT U3760 ( .A(n3081), .Y(n3829) );
  IBUFFX2_LVT U3761 ( .A(n6765), .Y(n3805) );
  AND2X4_LVT U3762 ( .A1(n5453), .A2(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(
        n6765) );
  IBUFFX2_LVT U3763 ( .A(n3805), .Y(n3804) );
  IBUFFX2_LVT U3764 ( .A(n3012), .Y(n9008) );
  DELLN1X2_LVT U3765 ( .A(n3803), .Y(n2875) );
  IBUFFX2_LVT U3766 ( .A(n3186), .Y(n4351) );
  AOI21X2_LVT U3767 ( .A1(n3841), .A2(csr_io_rw_rdata[4]), .A3(n5529), .Y(
        n3190) );
  IBUFFX2_LVT U3768 ( .A(n3190), .Y(n4330) );
  IBUFFX2_LVT U3769 ( .A(n3692), .Y(n3989) );
  IBUFFX2_LVT U3770 ( .A(n3692), .Y(n2969) );
  IBUFFX2_LVT U3771 ( .A(n3692), .Y(n3988) );
  IBUFFX2_LVT U3772 ( .A(n6871), .Y(n3876) );
  AND2X4_LVT U3773 ( .A1(n5449), .A2(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(
        n6871) );
  IBUFFX2_LVT U3774 ( .A(n3876), .Y(n3875) );
  IBUFFX2_LVT U3775 ( .A(n3876), .Y(n3874) );
  IBUFFX2_LVT U3776 ( .A(n3783), .Y(n2552) );
  IBUFFX2_LVT U3777 ( .A(n9524), .Y(n9446) );
  NBUFFX2_LVT U3778 ( .A(n9036), .Y(n3060) );
  NBUFFX2_LVT U3779 ( .A(n9036), .Y(n2982) );
  IBUFFX2_LVT U3780 ( .A(n3184), .Y(n4023) );
  IBUFFX2_LVT U3781 ( .A(n3184), .Y(n4025) );
  IBUFFX2_LVT U3782 ( .A(n3184), .Y(n4024) );
  IBUFFX2_LVT U3783 ( .A(n6422), .Y(n6866) );
  DELLN1X2_LVT U3784 ( .A(n6866), .Y(n3864) );
  IBUFFX2_LVT U3785 ( .A(n6767), .Y(n6867) );
  DELLN1X2_LVT U3786 ( .A(n6867), .Y(n3865) );
  IBUFFX2_LVT U3787 ( .A(io_fpu_inst[12]), .Y(n3583) );
  IBUFFX2_LVT U3788 ( .A(clock), .Y(n3784) );
  DELLN1X2_LVT U3789 ( .A(n4499), .Y(n3594) );
  DELLN1X2_LVT U3790 ( .A(n4499), .Y(n3595) );
  INVX1_LVT U3791 ( .A(n3101), .Y(n2497) );
  INVX1_LVT U3792 ( .A(n3246), .Y(n2498) );
  AOI21X2_LVT U3793 ( .A1(io_fpu_inst[25]), .A2(n1847), .A3(n1828), .Y(n4855)
         );
  NAND3X2_LVT U3794 ( .A1(n9075), .A2(n9522), .A3(n9435), .Y(n4856) );
  NAND3X2_LVT U3795 ( .A1(io_fpu_inst[24]), .A2(n9522), .A3(io_fpu_inst[21]), 
        .Y(n5151) );
  AND2X1_LVT U3806 ( .A1(n1699), .A2(n3039), .Y(n2512) );
  AND2X1_LVT U3813 ( .A1(div_io_req_ready), .A2(n9422), .Y(n2524) );
  NBUFFX2_LVT U3814 ( .A(n2527), .Y(n2526) );
  NAND2X0_LVT U3815 ( .A1(n2527), .A2(n_T_427[424]), .Y(n8219) );
  NAND2X0_LVT U3816 ( .A1(n2527), .A2(n_T_427[436]), .Y(n2598) );
  NAND2X0_LVT U3817 ( .A1(n2527), .A2(n_T_427[429]), .Y(n8395) );
  NAND2X0_LVT U3818 ( .A1(n2527), .A2(n_T_427[446]), .Y(n8998) );
  NAND2X0_LVT U3819 ( .A1(n2527), .A2(n_T_427[441]), .Y(n8811) );
  NAND2X0_LVT U3820 ( .A1(n2527), .A2(n_T_427[423]), .Y(n8157) );
  NAND2X0_LVT U3821 ( .A1(n2527), .A2(n_T_427[417]), .Y(n7963) );
  NAND2X0_LVT U3822 ( .A1(n2527), .A2(n_T_427[437]), .Y(n8641) );
  NAND2X0_LVT U3823 ( .A1(n2526), .A2(n_T_427[432]), .Y(n8486) );
  NAND2X0_LVT U3824 ( .A1(n2526), .A2(n_T_427[419]), .Y(n8025) );
  NAND2X0_LVT U3825 ( .A1(n2526), .A2(n_T_427[421]), .Y(n8106) );
  NAND2X0_LVT U3826 ( .A1(n2526), .A2(n_T_427[438]), .Y(n8679) );
  AND2X4_LVT U3827 ( .A1(n8105), .A2(n3968), .Y(n2527) );
  NAND3X0_LVT U3828 ( .A1(n5142), .A2(n9437), .A3(n9443), .Y(n2528) );
  NAND2X0_LVT U3829 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[24]), .Y(n7683)
         );
  NAND2X0_LVT U3830 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[16]), .Y(n7442)
         );
  NAND2X0_LVT U3831 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[21]), .Y(n7591)
         );
  NAND2X0_LVT U3832 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[18]), .Y(n7499)
         );
  NAND2X0_LVT U3833 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[19]), .Y(n7532)
         );
  NAND2X0_LVT U3834 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[20]), .Y(n7559)
         );
  NAND2X0_LVT U3835 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[22]), .Y(n7622)
         );
  NAND2X0_LVT U3836 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[23]), .Y(n7655)
         );
  NAND2X0_LVT U3837 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[25]), .Y(n7718)
         );
  NAND2X0_LVT U3838 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[26]), .Y(n7751)
         );
  NAND2X0_LVT U3839 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[27]), .Y(n7783)
         );
  NAND2X0_LVT U3840 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[28]), .Y(n7815)
         );
  NAND2X0_LVT U3841 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[29]), .Y(n7848)
         );
  NAND2X0_LVT U3842 ( .A1(n2529), .A2(n1859), .Y(n7875) );
  NAND2X0_LVT U3843 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_inst_rs3_4_), .Y(
        n7903) );
  AND3X1_LVT U3844 ( .A1(n8943), .A2(n8945), .A3(n2531), .Y(n2530) );
  NAND2X0_LVT U3845 ( .A1(n3707), .A2(n_T_427[125]), .Y(n2531) );
  NAND4X0_LVT U3846 ( .A1(n2630), .A2(n2670), .A3(n9446), .A4(n9104), .Y(n2629) );
  AND2X4_LVT U3847 ( .A1(n3590), .A2(io_fpu_inst[6]), .Y(n5163) );
  AND3X1_LVT U3848 ( .A1(n6908), .A2(n6909), .A3(n6907), .Y(n2532) );
  OA21X1_LVT U3849 ( .A1(n9395), .A2(n9386), .A3(n9397), .Y(n9388) );
  AND3X1_LVT U3850 ( .A1(n3073), .A2(n6913), .A3(n6935), .Y(n6914) );
  NOR2X0_LVT U3851 ( .A1(n6910), .A2(n6911), .Y(n2533) );
  AND3X1_LVT U3852 ( .A1(n2534), .A2(n2535), .A3(n2536), .Y(n3737) );
  AND3X1_LVT U3853 ( .A1(n8627), .A2(n8626), .A3(n8625), .Y(n2534) );
  AND2X1_LVT U3854 ( .A1(n8632), .A2(n2617), .Y(n2535) );
  AND2X1_LVT U3855 ( .A1(n8629), .A2(n8628), .Y(n2536) );
  NAND2X0_LVT U3856 ( .A1(n4844), .A2(n4845), .Y(n2538) );
  NAND4X1_LVT U3857 ( .A1(n5162), .A2(n5161), .A3(n2624), .A4(n2623), .Y(n2539) );
  OR2X2_LVT U3858 ( .A1(n9524), .A2(n3078), .Y(n9079) );
  NAND3X1_LVT U3859 ( .A1(n5067), .A2(n9524), .A3(n9528), .Y(n1531) );
  OR2X2_LVT U3860 ( .A1(io_fpu_inst[12]), .A2(n9524), .Y(n5075) );
  NBUFFX2_LVT U3861 ( .A(n9521), .Y(io_fpu_inst[27]) );
  OR2X4_LVT U3862 ( .A1(n9520), .A2(n9521), .Y(n5099) );
  OA22X2_LVT U3863 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .Y(n5160)
         );
  NAND3X0_LVT U3864 ( .A1(n2541), .A2(n2542), .A3(n2543), .Y(N724) );
  AND4X1_LVT U3865 ( .A1(n2956), .A2(n2957), .A3(n8350), .A4(n2590), .Y(n2541)
         );
  AND3X1_LVT U3866 ( .A1(n8357), .A2(n8356), .A3(n8355), .Y(n2542) );
  AND3X2_LVT U3867 ( .A1(n6991), .A2(n9288), .A3(n6992), .Y(n2544) );
  OR2X2_LVT U3868 ( .A1(n9111), .A2(n5073), .Y(n5077) );
  AND2X4_LVT U3869 ( .A1(n6238), .A2(n5437), .Y(n5446) );
  AND2X4_LVT U3870 ( .A1(n6238), .A2(n5448), .Y(n5457) );
  NAND4X1_LVT U3871 ( .A1(n5433), .A2(n5430), .A3(n5432), .A4(n5431), .Y(n6238) );
  NAND3X0_LVT U3872 ( .A1(n6991), .A2(n9288), .A3(n6992), .Y(n1262) );
  NBUFFX2_LVT U3873 ( .A(n9527), .Y(io_fpu_inst[4]) );
  NAND2X0_LVT U3874 ( .A1(n_T_427[1899]), .A2(n3992), .Y(n7483) );
  AOI21X2_LVT U3875 ( .A1(n3039), .A2(n5069), .A3(n5068), .Y(n5123) );
  OR2X2_LVT U3876 ( .A1(n5099), .A2(n2568), .Y(n2669) );
  OA21X2_LVT U3877 ( .A1(n3276), .A2(n3993), .A3(n7934), .Y(n7937) );
  OR2X4_LVT U3878 ( .A1(n3531), .A2(n3993), .Y(n7077) );
  OR2X4_LVT U3879 ( .A1(n2496), .A2(n3993), .Y(n8352) );
  OR2X4_LVT U3880 ( .A1(n3277), .A2(n3993), .Y(n2593) );
  NAND2X0_LVT U3881 ( .A1(n3782), .A2(n3588), .Y(n9288) );
  NOR3X4_LVT U3882 ( .A1(io_fpu_inst[29]), .A2(n5130), .A3(io_fpu_inst[7]), 
        .Y(n5131) );
  AND4X2_LVT U3883 ( .A1(n9230), .A2(io_fpu_inst[6]), .A3(io_fpu_inst[29]), 
        .A4(n5136), .Y(n5137) );
  AND2X1_LVT U3884 ( .A1(n2544), .A2(n6906), .Y(n2548) );
  IBUFFX2_LVT U3885 ( .A(n9519), .Y(n9436) );
  NAND3X2_LVT U3886 ( .A1(n5138), .A2(n9445), .A3(io_fpu_inst[29]), .Y(n2641)
         );
  NAND3X2_LVT U3887 ( .A1(io_fpu_inst[29]), .A2(n3078), .A3(n9445), .Y(n5152)
         );
  NAND3X0_LVT U3888 ( .A1(n2549), .A2(n2550), .A3(n2551), .Y(N734) );
  AND3X1_LVT U3889 ( .A1(n8681), .A2(n8680), .A3(n8679), .Y(n2549) );
  AND3X1_LVT U3890 ( .A1(n3718), .A2(n3719), .A3(n3720), .Y(n2550) );
  NOR2X0_LVT U3891 ( .A1(n8705), .A2(n8706), .Y(n2551) );
  DELLN2X2_LVT U3892 ( .A(n9529), .Y(io_fpu_inst[2]) );
  AND2X4_LVT U3893 ( .A1(n9105), .A2(n9529), .Y(n9097) );
  AO21X2_LVT U3894 ( .A1(io_fpu_inst[13]), .A2(n9105), .A3(n9529), .Y(n5100)
         );
  NAND3X2_LVT U3895 ( .A1(io_dmem_resp_bits_replay), .A2(n2029), .A3(n2626), 
        .Y(n5403) );
  NAND2X0_LVT U3896 ( .A1(n4351), .A2(n3060), .Y(n2595) );
  DELLN3X2_LVT U3897 ( .A(n9036), .Y(n3665) );
  AND2X1_LVT U3898 ( .A1(n3765), .A2(n6923), .Y(n3773) );
  IBUFFX2_LVT U3899 ( .A(n5134), .Y(n5132) );
  NAND4X1_LVT U3900 ( .A1(n5166), .A2(n3049), .A3(n2130), .A4(io_fpu_inst[26]), 
        .Y(n6964) );
  NOR3X4_LVT U3901 ( .A1(n9438), .A2(n9110), .A3(n5129), .Y(n5070) );
  OR3X2_LVT U3902 ( .A1(io_fpu_inst[31]), .A2(io_fpu_inst[14]), .A3(n5129), 
        .Y(n5134) );
  AND2X1_LVT U3903 ( .A1(n6923), .A2(n6922), .Y(n6975) );
  IBUFFX2_LVT U3904 ( .A(n9518), .Y(n9435) );
  NBUFFX2_LVT U3905 ( .A(n9520), .Y(io_fpu_inst[28]) );
  OR2X2_LVT U3906 ( .A1(n8424), .A2(n3632), .Y(n8425) );
  NAND3X0_LVT U3907 ( .A1(n2555), .A2(n2556), .A3(n2557), .Y(N717) );
  AND3X1_LVT U3908 ( .A1(n2952), .A2(n2951), .A3(n2950), .Y(n2555) );
  AND3X1_LVT U3909 ( .A1(n8108), .A2(n8107), .A3(n8106), .Y(n2556) );
  NAND3X0_LVT U3910 ( .A1(n2558), .A2(n2559), .A3(n2560), .Y(N712) );
  AND3X1_LVT U3911 ( .A1(n7909), .A2(n7908), .A3(n7907), .Y(n2558) );
  AND3X1_LVT U3912 ( .A1(n7924), .A2(n7923), .A3(n7922), .Y(n2559) );
  AND3X1_LVT U3913 ( .A1(n2919), .A2(n2918), .A3(n2585), .Y(n2560) );
  AND2X1_LVT U3914 ( .A1(n6964), .A2(n2548), .Y(n6923) );
  NAND3X0_LVT U3915 ( .A1(n2562), .A2(n2563), .A3(n2564), .Y(N731) );
  AND3X1_LVT U3916 ( .A1(n8575), .A2(n8574), .A3(n8573), .Y(n2562) );
  AND3X1_LVT U3917 ( .A1(n3725), .A2(n3726), .A3(n3727), .Y(n2563) );
  NOR2X0_LVT U3918 ( .A1(n8600), .A2(n8599), .Y(n2564) );
  AND4X2_LVT U3919 ( .A1(n9442), .A2(n9438), .A3(n9441), .A4(n5148), .Y(n2565)
         );
  AO21X1_LVT U3920 ( .A1(n2629), .A2(n5108), .A3(n2669), .Y(n5165) );
  NAND3X1_LVT U3921 ( .A1(n9445), .A2(n3078), .A3(n2618), .Y(n3580) );
  NAND3X2_LVT U3922 ( .A1(n6995), .A2(n9288), .A3(n6992), .Y(n6944) );
  NAND3X1_LVT U3923 ( .A1(n6993), .A2(n572), .A3(n6992), .Y(n6994) );
  OR2X4_LVT U3924 ( .A1(n5051), .A2(n6992), .Y(n9281) );
  NAND4X1_LVT U3925 ( .A1(n4758), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .A3(
        n4757), .A4(n6963), .Y(n4759) );
  OA21X2_LVT U3926 ( .A1(n4996), .A2(n4995), .A3(n2825), .Y(n4997) );
  OR3X2_LVT U3927 ( .A1(n2878), .A2(ibuf_io_inst_0_bits_inst_rs2[4]), .A3(
        n5435), .Y(n5421) );
  AND2X1_LVT U3928 ( .A1(ibuf_io_inst_0_bits_inst_rs2[3]), .A2(
        ibuf_io_inst_0_bits_inst_rs2[4]), .Y(n5437) );
  XOR2X1_LVT U3929 ( .A1(n3782), .A2(n2566), .Y(n3581) );
  AND3X2_LVT U3930 ( .A1(n2068), .A2(n6957), .A3(n6975), .Y(n3769) );
  AND3X2_LVT U3931 ( .A1(n6975), .A2(n6954), .A3(n6973), .Y(n9015) );
  IBUFFX2_LVT U3932 ( .A(n9527), .Y(n3577) );
  AND4X1_LVT U3933 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n2625), .Y(n2567)
         );
  NAND4X1_LVT U3934 ( .A1(n9442), .A2(n9438), .A3(n9441), .A4(n5148), .Y(n5143) );
  AND3X2_LVT U3935 ( .A1(n9107), .A2(io_fpu_inst[5]), .A3(n9108), .Y(n1823) );
  AND3X2_LVT U3936 ( .A1(n2671), .A2(n2561), .A3(n6922), .Y(n3715) );
  NAND3X2_LVT U3937 ( .A1(n4857), .A2(io_fpu_inst[5]), .A3(n9104), .Y(n1532)
         );
  OR2X2_LVT U3938 ( .A1(io_fpu_inst[5]), .A2(io_fpu_inst[12]), .Y(n5133) );
  NAND3X2_LVT U3939 ( .A1(n9440), .A2(io_fpu_inst[4]), .A3(n9443), .Y(n5130)
         );
  NOR3X2_LVT U3940 ( .A1(n1262), .A2(n6935), .A3(n2968), .Y(n6937) );
  IBUFFX2_LVT U3941 ( .A(io_fpu_inst[26]), .Y(n9439) );
  AND2X4_LVT U3942 ( .A1(n2981), .A2(n6796), .Y(n6886) );
  AND2X4_LVT U3943 ( .A1(n6877), .A2(n3836), .Y(n6887) );
  AND2X4_LVT U3944 ( .A1(n6877), .A2(n3812), .Y(n6885) );
  AND2X4_LVT U3945 ( .A1(n2981), .A2(n3863), .Y(n6812) );
  AND2X4_LVT U3946 ( .A1(n2981), .A2(n3871), .Y(n6774) );
  AND2X4_LVT U3947 ( .A1(n6877), .A2(n3865), .Y(n6830) );
  AND2X4_LVT U3948 ( .A1(n6877), .A2(n3811), .Y(n6882) );
  AND2X4_LVT U3949 ( .A1(n6877), .A2(n6765), .Y(n6884) );
  AND2X4_LVT U3950 ( .A1(n2981), .A2(n3840), .Y(n6888) );
  AND2X4_LVT U3951 ( .A1(n2981), .A2(n3859), .Y(n6773) );
  AND2X4_LVT U3952 ( .A1(n6877), .A2(n6868), .Y(n6810) );
  AND2X4_LVT U3953 ( .A1(n6877), .A2(n6871), .Y(n6813) );
  NAND3X2_LVT U3954 ( .A1(n3773), .A2(n6973), .A3(n6972), .Y(n3663) );
  AND3X2_LVT U3955 ( .A1(n6973), .A2(n6948), .A3(n3709), .Y(n3666) );
  AND3X2_LVT U3956 ( .A1(n6975), .A2(n6948), .A3(n6973), .Y(n9030) );
  AND3X2_LVT U3957 ( .A1(n6973), .A2(n6972), .A3(n2983), .Y(n3768) );
  NAND4X1_LVT U3958 ( .A1(n5148), .A2(io_fpu_inst[28]), .A3(n9445), .A4(n9440), 
        .Y(n5150) );
  OR2X2_LVT U3959 ( .A1(n3079), .A2(n9520), .Y(n5129) );
  NAND3X2_LVT U3960 ( .A1(n2650), .A2(n6923), .A3(n6922), .Y(n3012) );
  AND3X2_LVT U3961 ( .A1(n6941), .A2(n6974), .A3(n6940), .Y(n9021) );
  AND3X2_LVT U3962 ( .A1(n6940), .A2(n6972), .A3(n3772), .Y(n9012) );
  AND2X4_LVT U3963 ( .A1(n2143), .A2(n6917), .Y(n6940) );
  INVX1_LVT U3964 ( .A(n9418), .Y(io_imem_req_valid) );
  IBUFFX2_LVT U3965 ( .A(n3683), .Y(n2645) );
  INVX1_LVT U3966 ( .A(n9383), .Y(n6995) );
  NOR4X1_LVT U3967 ( .A1(n1917), .A2(n9284), .A3(n9283), .A4(n9285), .Y(n1822)
         );
  AND2X1_LVT U3968 ( .A1(n6962), .A2(n6965), .Y(n6922) );
  INVX1_LVT U3969 ( .A(io_dmem_req_bits_addr[38]), .Y(n9328) );
  INVX1_LVT U3970 ( .A(n9280), .Y(n2834) );
  INVX1_LVT U3971 ( .A(n5021), .Y(n4934) );
  INVX1_LVT U3972 ( .A(n9099), .Y(n2675) );
  INVX1_LVT U3973 ( .A(n4040), .Y(n4038) );
  NOR2X1_LVT U3974 ( .A1(n9243), .A2(bpu_io_xcpt_if), .Y(n9099) );
  INVX1_LVT U3975 ( .A(n9413), .Y(n4931) );
  INVX1_LVT U3976 ( .A(n4040), .Y(n4039) );
  NOR2X0_LVT U3977 ( .A1(n6991), .A2(n2569), .Y(n2673) );
  INVX1_LVT U3978 ( .A(n6954), .Y(n4772) );
  INVX1_LVT U3979 ( .A(n6957), .Y(n4771) );
  INVX1_LVT U3980 ( .A(n4040), .Y(n9040) );
  INVX1_LVT U3981 ( .A(bpu_io_xcpt_if), .Y(n9244) );
  INVX1_LVT U3982 ( .A(n4729), .Y(n4707) );
  INVX1_LVT U3983 ( .A(n6948), .Y(n4773) );
  INVX1_LVT U3984 ( .A(n4364), .Y(n3710) );
  INVX1_LVT U3985 ( .A(n6972), .Y(n4774) );
  INVX1_LVT U3986 ( .A(n4318), .Y(n3686) );
  AND3X1_LVT U3987 ( .A1(n2570), .A2(n3077), .A3(n9446), .Y(n5396) );
  INVX1_LVT U3988 ( .A(n9288), .Y(n2569) );
  INVX1_LVT U3989 ( .A(n9109), .Y(n9073) );
  INVX1_LVT U3990 ( .A(n4691), .Y(n4692) );
  INVX1_LVT U3991 ( .A(n4401), .Y(n3645) );
  INVX1_LVT U3992 ( .A(n4445), .Y(n3660) );
  AND2X1_LVT U3993 ( .A1(n4642), .A2(ibuf_io_inst_0_bits_inst_rd[1]), .Y(n4729) );
  INVX1_LVT U3994 ( .A(n3097), .Y(n4388) );
  NOR2X0_LVT U3995 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(
        ibuf_io_inst_0_bits_inst_rd[1]), .Y(n4731) );
  INVX1_LVT U3996 ( .A(n4321), .Y(n3679) );
  AND2X1_LVT U3997 ( .A1(n4971), .A2(n2038), .Y(n6946) );
  INVX1_LVT U3998 ( .A(n5144), .Y(n5139) );
  INVX1_LVT U3999 ( .A(ibuf_io_inst_0_bits_inst_rd[0]), .Y(n4642) );
  INVX1_LVT U4000 ( .A(n9089), .Y(n9091) );
  INVX1_LVT U4001 ( .A(n5086), .Y(n9108) );
  INVX1_LVT U4002 ( .A(n3099), .Y(n4403) );
  INVX1_LVT U4003 ( .A(ibuf_io_inst_0_bits_inst_rd[4]), .Y(n4719) );
  INVX1_LVT U4004 ( .A(ibuf_io_inst_0_bits_inst_rd[1]), .Y(n4641) );
  INVX1_LVT U4005 ( .A(n3090), .Y(n4395) );
  INVX1_LVT U4006 ( .A(n4398), .Y(n3711) );
  INVX1_LVT U4007 ( .A(n4436), .Y(n3688) );
  INVX1_LVT U4008 ( .A(n9511), .Y(n9346) );
  INVX1_LVT U4009 ( .A(n3091), .Y(n4408) );
  INVX1_LVT U4010 ( .A(n9507), .Y(n9348) );
  INVX1_LVT U4011 ( .A(io_fpu_inst[20]), .Y(n9444) );
  INVX1_LVT U4012 ( .A(n3183), .Y(n4413) );
  INVX1_LVT U4013 ( .A(io_fpu_inst[9]), .Y(n3587) );
  INVX1_LVT U4014 ( .A(n4475), .Y(n3644) );
  INVX1_LVT U4015 ( .A(n2981), .Y(n3586) );
  NOR2X1_LVT U4016 ( .A1(io_fpu_inst[23]), .A2(io_fpu_inst[7]), .Y(n2616) );
  INVX1_LVT U4017 ( .A(n3092), .Y(n4356) );
  INVX1_LVT U4018 ( .A(ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4662) );
  INVX1_LVT U4019 ( .A(n4858), .Y(n4634) );
  INVX1_LVT U4020 ( .A(n3094), .Y(n4380) );
  INVX1_LVT U4021 ( .A(n3093), .Y(n4361) );
  INVX1_LVT U4022 ( .A(n9485), .Y(n9342) );
  INVX1_LVT U4023 ( .A(ibuf_io_inst_0_bits_inst_rs1[0]), .Y(n4747) );
  INVX1_LVT U4024 ( .A(n3096), .Y(n4390) );
  INVX0_LVT U4025 ( .A(ibuf_io_inst_0_bits_inst_rs1[1]), .Y(n2790) );
  INVX1_LVT U4026 ( .A(n4442), .Y(n3659) );
  INVX1_LVT U4027 ( .A(n9499), .Y(n9344) );
  INVX1_LVT U4028 ( .A(n9484), .Y(n9340) );
  INVX1_LVT U4029 ( .A(n9495), .Y(n9338) );
  INVX1_LVT U4030 ( .A(ibuf_io_inst_0_bits_replay), .Y(n9433) );
  INVX1_LVT U4031 ( .A(n4416), .Y(n3687) );
  INVX1_LVT U4032 ( .A(n5456), .Y(n4905) );
  INVX1_LVT U4033 ( .A(n5451), .Y(n4894) );
  INVX1_LVT U4034 ( .A(n3083), .Y(n3861) );
  NOR2X0_LVT U4035 ( .A1(n5436), .A2(n5435), .Y(n6837) );
  INVX1_LVT U4036 ( .A(n3083), .Y(n3862) );
  INVX1_LVT U4037 ( .A(n3095), .Y(n4378) );
  INVX1_LVT U4038 ( .A(n9425), .Y(n1281) );
  INVX1_LVT U4039 ( .A(n3098), .Y(n4421) );
  INVX1_LVT U4040 ( .A(n9503), .Y(n9336) );
  INVX1_LVT U4041 ( .A(n5454), .Y(n4873) );
  INVX1_LVT U4042 ( .A(n5449), .Y(n4874) );
  INVX1_LVT U4043 ( .A(n5450), .Y(n5438) );
  AND2X1_LVT U4044 ( .A1(n4890), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5451) );
  OR2X1_LVT U4045 ( .A1(n5434), .A2(n2878), .Y(n5447) );
  INVX1_LVT U4046 ( .A(n5452), .Y(n4906) );
  INVX1_LVT U4047 ( .A(n4890), .Y(n4898) );
  AND2X1_LVT U4048 ( .A1(n4889), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5450) );
  AND2X1_LVT U4049 ( .A1(n4900), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5449) );
  INVX1_LVT U4050 ( .A(n4889), .Y(n4899) );
  INVX1_LVT U4051 ( .A(n4860), .Y(n4633) );
  INVX0_LVT U4052 ( .A(ibuf_io_inst_0_bits_rvc), .Y(n4497) );
  INVX0_LVT U4053 ( .A(n9332), .Y(n9378) );
  INVX1_LVT U4054 ( .A(n3185), .Y(n2572) );
  INVX1_LVT U4055 ( .A(ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n4815) );
  OR2X1_LVT U4056 ( .A1(n9399), .A2(n9398), .Y(n9402) );
  INVX1_LVT U4057 ( .A(n5358), .Y(n5304) );
  AND2X1_LVT U4058 ( .A1(n5358), .A2(n5302), .Y(n3185) );
  AOI21X1_LVT U4059 ( .A1(n9256), .A2(n9255), .A3(n9254), .Y(n9276) );
  INVX1_LVT U4060 ( .A(n5254), .Y(n5256) );
  INVX1_LVT U4061 ( .A(io_fpu_fromint_data[62]), .Y(n9307) );
  INVX1_LVT U4062 ( .A(io_fpu_fromint_data[63]), .Y(n9308) );
  INVX1_LVT U4063 ( .A(io_fpu_fromint_data[61]), .Y(n9309) );
  INVX1_LVT U4064 ( .A(io_fpu_fromint_data[59]), .Y(n9310) );
  INVX1_LVT U4065 ( .A(io_fpu_fromint_data[60]), .Y(n9303) );
  INVX1_LVT U4066 ( .A(io_fpu_fromint_data[58]), .Y(n9304) );
  INVX1_LVT U4067 ( .A(io_fpu_fromint_data[56]), .Y(n9305) );
  INVX1_LVT U4068 ( .A(io_fpu_fromint_data[57]), .Y(n9306) );
  AND3X1_LVT U4069 ( .A1(n9392), .A2(n2574), .A3(n2061), .Y(n9405) );
  INVX1_LVT U4070 ( .A(n9397), .Y(n9399) );
  INVX1_LVT U4071 ( .A(n9386), .Y(n9387) );
  INVX1_LVT U4072 ( .A(n9403), .Y(n9400) );
  AND3X1_LVT U4073 ( .A1(n5314), .A2(n3046), .A3(n2575), .Y(n5307) );
  AND3X1_LVT U4074 ( .A1(n3046), .A2(n5351), .A3(n2575), .Y(n5357) );
  AND2X1_LVT U4075 ( .A1(n9120), .A2(ex_reg_rs_bypass_1), .Y(n9165) );
  AND2X1_LVT U4076 ( .A1(n9201), .A2(ex_ctrl_sel_alu2[1]), .Y(n9227) );
  NOR2X1_LVT U4077 ( .A1(n9201), .A2(n9200), .Y(n9222) );
  INVX1_LVT U4078 ( .A(wb_cause[0]), .Y(n9256) );
  INVX1_LVT U4079 ( .A(n5408), .Y(n5406) );
  INVX1_LVT U4080 ( .A(n5051), .Y(n5052) );
  INVX1_LVT U4081 ( .A(n5084), .Y(n5082) );
  INVX1_LVT U4082 ( .A(n5009), .Y(n4866) );
  INVX1_LVT U4083 ( .A(ibuf_io_inst_0_bits_raw[27]), .Y(n4781) );
  INVX1_LVT U4084 ( .A(n5301), .Y(n4944) );
  INVX0_LVT U4085 ( .A(n9179), .Y(n9201) );
  INVX1_LVT U4086 ( .A(n9172), .Y(n9174) );
  INVX1_LVT U4087 ( .A(n9178), .Y(n9180) );
  AND2X1_LVT U4088 ( .A1(n7017), .A2(n7019), .Y(n9064) );
  INVX1_LVT U4089 ( .A(n5326), .Y(n5327) );
  INVX1_LVT U4090 ( .A(n5412), .Y(n5414) );
  INVX1_LVT U4091 ( .A(n5303), .Y(n5392) );
  INVX1_LVT U4092 ( .A(n5306), .Y(n5427) );
  INVX1_LVT U4093 ( .A(n5313), .Y(n2575) );
  INVX1_LVT U4094 ( .A(n4948), .Y(n4859) );
  INVX1_LVT U4095 ( .A(csr_io_status_isa[2]), .Y(n6912) );
  INVX1_LVT U4096 ( .A(div_io_req_ready), .Y(n4917) );
  INVX1_LVT U4097 ( .A(n9330), .Y(n9331) );
  INVX1_LVT U4098 ( .A(n5413), .Y(n6860) );
  INVX0_LVT U4099 ( .A(reset), .Y(n4498) );
  INVX1_LVT U4100 ( .A(io_fpu_dec_ren2), .Y(n4837) );
  INVX1_LVT U4101 ( .A(io_fpu_sboard_clra[0]), .Y(n5182) );
  INVX0_LVT U4102 ( .A(io_dmem_s2_xcpt_pf_ld), .Y(n9246) );
  INVX1_LVT U4103 ( .A(io_fpu_dmem_resp_tag[0]), .Y(n5184) );
  INVX0_LVT U4104 ( .A(io_dmem_s2_xcpt_ma_ld), .Y(n9247) );
  INVX1_LVT U4105 ( .A(io_fpu_dec_ren3), .Y(n4838) );
  INVX0_LVT U4106 ( .A(n2030), .Y(n4943) );
  INVX1_LVT U4107 ( .A(io_fpu_sboard_clra[2]), .Y(n5257) );
  INVX1_LVT U4108 ( .A(io_fpu_dec_ren1), .Y(n4945) );
  INVX1_LVT U4109 ( .A(io_fpu_sboard_clr), .Y(n5177) );
  INVX1_LVT U4110 ( .A(io_fpu_dmem_resp_tag[2]), .Y(n5259) );
  NAND4X0_LVT U4111 ( .A1(n3023), .A2(n2655), .A3(n3705), .A4(n3022), .Y(N701)
         );
  NOR2X1_LVT U4112 ( .A1(n8835), .A2(n8836), .Y(n3732) );
  NOR2X1_LVT U4113 ( .A1(n8872), .A2(n8871), .Y(n3729) );
  NAND4X0_LVT U4114 ( .A1(n3021), .A2(n2651), .A3(n3020), .A4(n3696), .Y(N697)
         );
  NOR2X1_LVT U4115 ( .A1(n9033), .A2(n9034), .Y(n3749) );
  OA21X1_LVT U4116 ( .A1(n3476), .A2(n3994), .A3(n8553), .Y(n8556) );
  AND3X1_LVT U4117 ( .A1(n7545), .A2(n2664), .A3(n2663), .Y(n2662) );
  AO21X1_LVT U4118 ( .A1(n7350), .A2(n7351), .A3(n2645), .Y(n7352) );
  OR2X1_LVT U4119 ( .A1(n8842), .A2(n2645), .Y(n8843) );
  OR2X1_LVT U4120 ( .A1(n3371), .A2(n3988), .Y(n2661) );
  OR2X1_LVT U4121 ( .A1(n3309), .A2(n4012), .Y(n2607) );
  AOI22X1_LVT U4122 ( .A1(n_T_427[1162]), .A2(n2611), .A3(n3639), .A4(
        n_T_427[1226]), .Y(n7301) );
  AOI21X1_LVT U4123 ( .A1(n3717), .A2(n_T_427[1078]), .A3(n3776), .Y(n8740) );
  AOI21X1_LVT U4124 ( .A1(n3717), .A2(n_T_427[1064]), .A3(n3777), .Y(n8256) );
  OA21X1_LVT U4125 ( .A1(n2081), .A2(n3306), .A3(n8975), .Y(n8978) );
  OA21X1_LVT U4126 ( .A1(n4008), .A2(n3336), .A3(n8113), .Y(n8116) );
  OR2X1_LVT U4127 ( .A1(n3341), .A2(n4011), .Y(n2608) );
  OR2X1_LVT U4128 ( .A1(n8319), .A2(n2154), .Y(n8320) );
  OA21X1_LVT U4129 ( .A1(n3664), .A2(n3298), .A3(n7970), .Y(n7973) );
  OA21X1_LVT U4130 ( .A1(n2081), .A2(n3342), .A3(n8362), .Y(n8365) );
  OA21X1_LVT U4131 ( .A1(n4009), .A2(n3354), .A3(n8595), .Y(n8598) );
  OR2X1_LVT U4132 ( .A1(n9088), .A2(n1431), .Y(n9233) );
  NAND4X0_LVT U4133 ( .A1(n2677), .A2(n9231), .A3(io_fpu_inst[30]), .A4(n9230), 
        .Y(n9232) );
  OR2X1_LVT U4134 ( .A1(n9077), .A2(n1431), .Y(n9228) );
  INVX0_LVT U4135 ( .A(n2984), .Y(n4011) );
  NBUFFX2_LVT U4136 ( .A(n3658), .Y(n2897) );
  XOR2X1_LVT U4137 ( .A1(n9377), .A2(ibuf_io_pc[39]), .Y(n4574) );
  AO21X1_LVT U4138 ( .A1(n9439), .A2(n2539), .A3(n3075), .Y(n6936) );
  XOR2X1_LVT U4139 ( .A1(n9508), .A2(ibuf_io_pc[36]), .Y(n4565) );
  XOR2X1_LVT U4140 ( .A1(n9498), .A2(ibuf_io_pc[38]), .Y(n4521) );
  XOR2X1_LVT U4141 ( .A1(n9505), .A2(ibuf_io_pc[32]), .Y(n4593) );
  NOR2X1_LVT U4142 ( .A1(n5845), .A2(n5844), .Y(n5855) );
  NOR2X1_LVT U4143 ( .A1(n5566), .A2(n5565), .Y(n5576) );
  NOR2X1_LVT U4144 ( .A1(n5935), .A2(n5934), .Y(n5945) );
  XOR2X1_LVT U4145 ( .A1(n9493), .A2(ibuf_io_pc[33]), .Y(n4583) );
  NOR2X1_LVT U4146 ( .A1(n5658), .A2(n5657), .Y(n5668) );
  XOR2X1_LVT U4147 ( .A1(n9374), .A2(ibuf_io_pc[35]), .Y(n4576) );
  XOR2X1_LVT U4148 ( .A1(n9502), .A2(ibuf_io_pc[31]), .Y(n4563) );
  XOR2X1_LVT U4149 ( .A1(n9373), .A2(n4557), .Y(n4558) );
  NOR2X1_LVT U4150 ( .A1(n6330), .A2(n6329), .Y(n6340) );
  NOR2X1_LVT U4151 ( .A1(n6495), .A2(n6494), .Y(n6505) );
  NOR2X1_LVT U4152 ( .A1(n6172), .A2(n6171), .Y(n6182) );
  NOR2X1_LVT U4153 ( .A1(n5979), .A2(n5978), .Y(n5989) );
  NOR2X1_LVT U4154 ( .A1(n5515), .A2(n5514), .Y(n5525) );
  OA22X1_LVT U4155 ( .A1(n3559), .A2(n3882), .A3(n3877), .A4(n6549), .Y(n6552)
         );
  OA22X1_LVT U4156 ( .A1(n3539), .A2(n3880), .A3(n3879), .A4(n5751), .Y(n5753)
         );
  OA22X1_LVT U4157 ( .A1(n3542), .A2(n3881), .A3(n3879), .A4(n5813), .Y(n5814)
         );
  AOI22X1_LVT U4158 ( .A1(n3834), .A2(n_T_427[405]), .A3(n_T_427[469]), .A4(
        n2824), .Y(n2845) );
  OA22X1_LVT U4159 ( .A1(n3564), .A2(n3882), .A3(n1993), .A4(n6674), .Y(n6677)
         );
  OA22X1_LVT U4160 ( .A1(n3533), .A2(n3880), .A3(n3879), .A4(n5595), .Y(n5598)
         );
  OA22X1_LVT U4161 ( .A1(n3560), .A2(n3882), .A3(n1993), .A4(n6577), .Y(n6580)
         );
  AOI22X1_LVT U4162 ( .A1(n5776), .A2(n1992), .A3(n_T_427[1897]), .A4(n3884), 
        .Y(n2756) );
  OA22X1_LVT U4163 ( .A1(n3540), .A2(n3880), .A3(n3879), .A4(n5784), .Y(n5788)
         );
  OA22X1_LVT U4164 ( .A1(n3558), .A2(n3882), .A3(n1993), .A4(n6500), .Y(n6502)
         );
  AOI22X1_LVT U4165 ( .A1(n2856), .A2(n_T_427[342]), .A3(n_T_427[86]), .A4(
        n2872), .Y(n2683) );
  AOI22X1_LVT U4166 ( .A1(n2872), .A2(n_T_427[71]), .A3(n_T_427[902]), .A4(
        n3897), .Y(n2729) );
  OA22X1_LVT U4167 ( .A1(n3562), .A2(n3882), .A3(n3877), .A4(n6622), .Y(n6625)
         );
  OA22X1_LVT U4168 ( .A1(n3277), .A2(n3882), .A3(n1993), .A4(n6525), .Y(n6527)
         );
  AOI22X1_LVT U4169 ( .A1(n5495), .A2(n6877), .A3(n_T_427[1884]), .A4(n3884), 
        .Y(n2789) );
  OA22X1_LVT U4170 ( .A1(n3536), .A2(n3880), .A3(n3879), .A4(n5663), .Y(n5666)
         );
  AOI22X1_LVT U4171 ( .A1(n5545), .A2(n6877), .A3(n_T_427[1886]), .A4(n3884), 
        .Y(n2785) );
  AND4X1_LVT U4172 ( .A1(n9096), .A2(n9095), .A3(n9109), .A4(n9094), .Y(n2676)
         );
  NOR2X1_LVT U4173 ( .A1(n6280), .A2(n6279), .Y(n6290) );
  OA22X1_LVT U4174 ( .A1(n3538), .A2(n3880), .A3(n3879), .A4(n5712), .Y(n5714)
         );
  OA22X1_LVT U4175 ( .A1(n3531), .A2(n3880), .A3(n3879), .A4(n5520), .Y(n5523)
         );
  AOI22X1_LVT U4176 ( .A1(n6258), .A2(n6877), .A3(n_T_427[1919]), .A4(n3884), 
        .Y(n2760) );
  AOI22X1_LVT U4177 ( .A1(n3798), .A2(n_T_427[1762]), .A3(n_T_427[1823]), .A4(
        n3830), .Y(n2746) );
  AOI22X1_LVT U4178 ( .A1(n6772), .A2(n1992), .A3(n_T_427[1939]), .A4(n3884), 
        .Y(n2823) );
  AOI22X1_LVT U4179 ( .A1(n3901), .A2(n_T_427[1070]), .A3(n_T_427[239]), .A4(
        n6773), .Y(n2736) );
  AOI22X1_LVT U4180 ( .A1(n3835), .A2(n_T_427[431]), .A3(n_T_427[750]), .A4(
        n3905), .Y(n2737) );
  AOI22X1_LVT U4181 ( .A1(n3902), .A2(n_T_427[1081]), .A3(n_T_427[250]), .A4(
        n3807), .Y(n2732) );
  OR3X1_LVT U4182 ( .A1(n5133), .A2(n9109), .A3(n9096), .Y(n1612) );
  AOI22X1_LVT U4183 ( .A1(n2864), .A2(n_T_427[429]), .A3(n_T_427[109]), .A4(
        n3833), .Y(n2709) );
  OA22X1_LVT U4184 ( .A1(n3555), .A2(n3882), .A3(n3877), .A4(n6402), .Y(n6405)
         );
  OA22X1_LVT U4185 ( .A1(n3532), .A2(n3880), .A3(n3879), .A4(n5571), .Y(n5574)
         );
  OA22X1_LVT U4186 ( .A1(n3537), .A2(n3880), .A3(n3879), .A4(n5694), .Y(n5697)
         );
  AOI22X1_LVT U4187 ( .A1(n6376), .A2(n1992), .A3(n_T_427[1924]), .A4(n3884), 
        .Y(n2764) );
  NOR2X1_LVT U4188 ( .A1(n5689), .A2(n5688), .Y(n5699) );
  AOI22X1_LVT U4189 ( .A1(n2867), .A2(n_T_427[1756]), .A3(n_T_427[1818]), .A4(
        n3829), .Y(n2766) );
  XOR2X1_LVT U4190 ( .A1(n9486), .A2(ibuf_io_pc[20]), .Y(n4585) );
  XOR2X1_LVT U4191 ( .A1(n9501), .A2(ibuf_io_pc[22]), .Y(n4584) );
  OA22X1_LVT U4192 ( .A1(n3535), .A2(n3880), .A3(n3879), .A4(n5639), .Y(n5642)
         );
  XOR2X1_LVT U4193 ( .A1(n9364), .A2(ibuf_io_pc[24]), .Y(n4590) );
  XOR2X1_LVT U4194 ( .A1(n9368), .A2(ibuf_io_pc[28]), .Y(n4589) );
  XOR2X1_LVT U4195 ( .A1(n9488), .A2(ibuf_io_pc[23]), .Y(n4560) );
  XOR2X1_LVT U4196 ( .A1(n9483), .A2(ibuf_io_pc[26]), .Y(n4520) );
  XOR2X1_LVT U4197 ( .A1(n9489), .A2(ibuf_io_pc[27]), .Y(n4561) );
  OA22X1_LVT U4198 ( .A1(n3534), .A2(n3880), .A3(n3879), .A4(n5615), .Y(n5618)
         );
  AOI22X1_LVT U4199 ( .A1(n3893), .A2(n_T_427[1579]), .A3(n_T_427[1643]), .A4(
        n3887), .Y(n2763) );
  AOI22X1_LVT U4200 ( .A1(n3945), .A2(n_T_427[1194]), .A3(n_T_427[1258]), .A4(
        n3940), .Y(n2694) );
  XOR2X1_LVT U4201 ( .A1(n9506), .A2(ibuf_io_pc[14]), .Y(n4555) );
  AOI22X1_LVT U4202 ( .A1(n3945), .A2(n_T_427[1198]), .A3(n_T_427[1262]), .A4(
        n3939), .Y(n2734) );
  XOR2X1_LVT U4203 ( .A1(n9491), .A2(ibuf_io_pc[12]), .Y(n4554) );
  AOI22X1_LVT U4204 ( .A1(n3955), .A2(n_T_427[1130]), .A3(n_T_427[1002]), .A4(
        n3950), .Y(n2695) );
  AOI22X1_LVT U4205 ( .A1(n3955), .A2(n_T_427[1134]), .A3(n_T_427[1006]), .A4(
        n3949), .Y(n2735) );
  OR2X1_LVT U4206 ( .A1(n2644), .A2(n5143), .Y(n2643) );
  NOR2X1_LVT U4207 ( .A1(csr_io_interrupt), .A2(bpu_io_debug_if), .Y(n5167) );
  XOR2X1_LVT U4208 ( .A1(n9496), .A2(ibuf_io_pc[18]), .Y(n4556) );
  AOI22X1_LVT U4209 ( .A1(n3955), .A2(n_T_427[1132]), .A3(n_T_427[1004]), .A4(
        n3949), .Y(n2707) );
  AOI22X1_LVT U4210 ( .A1(n3945), .A2(n_T_427[1196]), .A3(n_T_427[1260]), .A4(
        n3939), .Y(n2706) );
  AOI22X1_LVT U4211 ( .A1(n3901), .A2(n_T_427[1059]), .A3(n_T_427[931]), .A4(
        n3895), .Y(n2740) );
  AOI22X1_LVT U4212 ( .A1(n2824), .A2(n_T_427[484]), .A3(n_T_427[739]), .A4(
        n3904), .Y(n2741) );
  AOI22X1_LVT U4213 ( .A1(n3955), .A2(n_T_427[1135]), .A3(n_T_427[1007]), .A4(
        n3950), .Y(n2723) );
  INVX1_LVT U4214 ( .A(n4040), .Y(n4037) );
  AOI22X1_LVT U4215 ( .A1(n3945), .A2(n_T_427[1191]), .A3(n_T_427[1255]), .A4(
        n3939), .Y(n2718) );
  AOI22X1_LVT U4216 ( .A1(n3955), .A2(n_T_427[1127]), .A3(n_T_427[999]), .A4(
        n3949), .Y(n2719) );
  NAND3X0_LVT U4217 ( .A1(n2565), .A2(n3078), .A3(n9436), .Y(n5146) );
  AOI22X1_LVT U4218 ( .A1(n2861), .A2(n_T_427[810]), .A3(n_T_427[746]), .A4(
        n3904), .Y(n2697) );
  XOR2X1_LVT U4219 ( .A1(n9497), .A2(ibuf_io_pc[25]), .Y(n4582) );
  AOI22X1_LVT U4220 ( .A1(n2866), .A2(n_T_427[1760]), .A3(n_T_427[1821]), .A4(
        n3829), .Y(n2751) );
  XOR2X1_LVT U4221 ( .A1(n9356), .A2(n4518), .Y(n4519) );
  AOI22X1_LVT U4222 ( .A1(n3945), .A2(n_T_427[1200]), .A3(n_T_427[1264]), .A4(
        n3939), .Y(n2698) );
  AOI22X1_LVT U4223 ( .A1(n3955), .A2(n_T_427[1136]), .A3(n_T_427[1008]), .A4(
        n3949), .Y(n2699) );
  AOI22X1_LVT U4224 ( .A1(n3890), .A2(n_T_427[1537]), .A3(n_T_427[1601]), .A4(
        n3885), .Y(n2788) );
  AOI22X1_LVT U4225 ( .A1(n3893), .A2(n_T_427[1581]), .A3(n_T_427[1645]), .A4(
        n3888), .Y(n2780) );
  AOI22X1_LVT U4226 ( .A1(n6428), .A2(n1992), .A3(n_T_427[1926]), .A4(n3884), 
        .Y(n2781) );
  AOI22X1_LVT U4227 ( .A1(n3924), .A2(n_T_427[1498]), .A3(n_T_427[1370]), .A4(
        n3918), .Y(n2773) );
  AOI22X1_LVT U4228 ( .A1(n3901), .A2(n_T_427[1068]), .A3(n_T_427[940]), .A4(
        n2831), .Y(n2708) );
  AOI22X1_LVT U4229 ( .A1(n3945), .A2(n_T_427[1199]), .A3(n_T_427[1263]), .A4(
        n3940), .Y(n2722) );
  AOI22X1_LVT U4230 ( .A1(n2861), .A2(n_T_427[788]), .A3(n_T_427[341]), .A4(
        n2857), .Y(n2843) );
  INVX1_LVT U4231 ( .A(n6949), .Y(n8982) );
  AOI22X1_LVT U4232 ( .A1(n2824), .A2(n_T_427[470]), .A3(n_T_427[917]), .A4(
        n2831), .Y(n2682) );
  NOR2X1_LVT U4233 ( .A1(n6956), .A2(n6947), .Y(n9038) );
  AOI22X1_LVT U4234 ( .A1(n3923), .A2(n_T_427[1491]), .A3(n_T_427[1363]), .A4(
        n3918), .Y(n2802) );
  AOI22X1_LVT U4235 ( .A1(n3956), .A2(n_T_427[1144]), .A3(n_T_427[1016]), .A4(
        n3951), .Y(n2743) );
  AOI22X1_LVT U4236 ( .A1(n3946), .A2(n_T_427[1208]), .A3(n_T_427[1272]), .A4(
        n3941), .Y(n2742) );
  AOI22X1_LVT U4237 ( .A1(n3927), .A2(n_T_427[1280]), .A3(n_T_427[1216]), .A4(
        n3937), .Y(n2855) );
  AOI22X1_LVT U4238 ( .A1(n2860), .A2(n_T_427[825]), .A3(n_T_427[761]), .A4(
        n3905), .Y(n2733) );
  AOI22X1_LVT U4239 ( .A1(n3956), .A2(n_T_427[1145]), .A3(n_T_427[1017]), .A4(
        n3951), .Y(n2731) );
  AOI22X1_LVT U4240 ( .A1(n3946), .A2(n_T_427[1209]), .A3(n_T_427[1273]), .A4(
        n3941), .Y(n2730) );
  INVX0_LVT U4241 ( .A(n6991), .Y(n6993) );
  AOI22X1_LVT U4242 ( .A1(n3923), .A2(n_T_427[1481]), .A3(n_T_427[1353]), .A4(
        n3917), .Y(n2794) );
  NOR2X1_LVT U4243 ( .A1(n1531), .A2(io_fpu_inst[14]), .Y(n5116) );
  AOI22X1_LVT U4244 ( .A1(n3924), .A2(n_T_427[1489]), .A3(n_T_427[1361]), .A4(
        n3918), .Y(n2818) );
  NAND2X0_LVT U4245 ( .A1(n5067), .A2(n3578), .Y(n2635) );
  AOI22X1_LVT U4246 ( .A1(n1919), .A2(n_T_427[337]), .A3(n_T_427[529]), .A4(
        n3819), .Y(n2679) );
  AOI22X1_LVT U4247 ( .A1(n3823), .A2(n_T_427[848]), .A3(n_T_427[657]), .A4(
        n3821), .Y(n2681) );
  AOI22X1_LVT U4248 ( .A1(n3894), .A2(n_T_427[1595]), .A3(n_T_427[1659]), .A4(
        n3888), .Y(n2822) );
  AOI22X1_LVT U4249 ( .A1(n3829), .A2(n_T_427[1846]), .A3(n_T_427[1723]), .A4(
        n3824), .Y(n2821) );
  AOI22X1_LVT U4250 ( .A1(n3907), .A2(n_T_427[786]), .A3(n_T_427[467]), .A4(
        n3910), .Y(n2839) );
  AOI22X1_LVT U4251 ( .A1(n3924), .A2(n_T_427[1480]), .A3(n_T_427[1352]), .A4(
        n3917), .Y(n2814) );
  AOI22X1_LVT U4252 ( .A1(n3955), .A2(n_T_427[1138]), .A3(n_T_427[1010]), .A4(
        n3950), .Y(n2711) );
  AOI22X1_LVT U4253 ( .A1(n3945), .A2(n_T_427[1202]), .A3(n_T_427[1266]), .A4(
        n3940), .Y(n2710) );
  AOI22X1_LVT U4254 ( .A1(n3956), .A2(n_T_427[1141]), .A3(n_T_427[1013]), .A4(
        n3951), .Y(n2691) );
  AOI22X1_LVT U4255 ( .A1(n3946), .A2(n_T_427[1205]), .A3(n_T_427[1269]), .A4(
        n3941), .Y(n2690) );
  AOI22X1_LVT U4256 ( .A1(n3818), .A2(n_T_427[512]), .A3(n_T_427[576]), .A4(
        n3916), .Y(n2880) );
  AOI22X1_LVT U4257 ( .A1(n3956), .A2(n_T_427[1143]), .A3(n_T_427[1015]), .A4(
        n3950), .Y(n2703) );
  AOI22X1_LVT U4258 ( .A1(n3946), .A2(n_T_427[1207]), .A3(n_T_427[1271]), .A4(
        n3940), .Y(n2702) );
  NAND3X0_LVT U4259 ( .A1(n3566), .A2(n5136), .A3(n3567), .Y(n2644) );
  INVX1_LVT U4260 ( .A(n3097), .Y(n4387) );
  NAND3X0_LVT U4261 ( .A1(n9076), .A2(n9075), .A3(io_fpu_inst[30]), .Y(n9077)
         );
  AND2X1_LVT U4262 ( .A1(n4749), .A2(n2038), .Y(n6954) );
  OR2X1_LVT U4263 ( .A1(n2825), .A2(n6955), .Y(n6949) );
  NOR2X1_LVT U4264 ( .A1(n6956), .A2(n6955), .Y(n3182) );
  INVX1_LVT U4265 ( .A(n6955), .Y(n6926) );
  INVX1_LVT U4266 ( .A(n4730), .Y(n4708) );
  INVX0_LVT U4267 ( .A(n4847), .Y(n4618) );
  NAND4X0_LVT U4268 ( .A1(n4690), .A2(n3046), .A3(n4689), .A4(n4688), .Y(n4695) );
  XOR2X1_LVT U4269 ( .A1(n9487), .A2(ibuf_io_pc[17]), .Y(n4551) );
  NAND4X0_LVT U4270 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n2625), .Y(n5036) );
  XOR2X1_LVT U4271 ( .A1(n9507), .A2(ibuf_io_pc[9]), .Y(n4547) );
  XOR2X1_LVT U4272 ( .A1(n9511), .A2(ibuf_io_pc[8]), .Y(n4549) );
  AND2X1_LVT U4273 ( .A1(n4641), .A2(ibuf_io_inst_0_bits_inst_rd[0]), .Y(n4732) );
  INVX1_LVT U4274 ( .A(n3195), .Y(n4358) );
  OR2X1_LVT U4275 ( .A1(io_fpu_inst[6]), .A2(io_fpu_inst[2]), .Y(n9109) );
  AOI21X1_LVT U4276 ( .A1(n3843), .A2(csr_io_rw_rdata[25]), .A3(n5953), .Y(
        n3097) );
  NAND4X0_LVT U4277 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n3046), .Y(n5003) );
  INVX1_LVT U4278 ( .A(n3195), .Y(n4357) );
  XOR2X1_LVT U4279 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n3202), .Y(n4946) );
  NAND4X0_LVT U4280 ( .A1(n9445), .A2(n1867), .A3(io_fpu_inst[6]), .A4(n3577), 
        .Y(n9081) );
  AO21X1_LVT U4281 ( .A1(io_fpu_inst[5]), .A2(io_fpu_inst[14]), .A3(
        io_fpu_inst[2]), .Y(n9094) );
  AND3X1_LVT U4282 ( .A1(n3044), .A2(io_fpu_inst[14]), .A3(n9435), .Y(n5107)
         );
  NAND2X0_LVT U4283 ( .A1(n5100), .A2(n2552), .Y(n2636) );
  NAND2X0_LVT U4284 ( .A1(n5446), .A2(n5452), .Y(n3082) );
  INVX1_LVT U4285 ( .A(n3189), .Y(n4345) );
  AO21X1_LVT U4286 ( .A1(io_fpu_inst[14]), .A2(n9105), .A3(n9435), .Y(n5097)
         );
  INVX1_LVT U4287 ( .A(n3192), .Y(n4342) );
  OR2X1_LVT U4288 ( .A1(io_fpu_inst[21]), .A2(io_fpu_inst[20]), .Y(n5394) );
  INVX1_LVT U4289 ( .A(n3193), .Y(n4354) );
  XOR2X1_LVT U4290 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n588), .Y(n5031)
         );
  XOR2X1_LVT U4291 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n590), .Y(n5033)
         );
  NOR4X0_LVT U4292 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n2877), .A3(
        ibuf_io_inst_0_bits_inst_rs1[0]), .A4(ibuf_io_inst_0_bits_inst_rs1[2]), 
        .Y(n3588) );
  NOR2X1_LVT U4293 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(
        ibuf_io_inst_0_bits_inst_rd[4]), .Y(n4700) );
  INVX1_LVT U4294 ( .A(n3192), .Y(n4340) );
  INVX1_LVT U4295 ( .A(ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4733) );
  INVX1_LVT U4296 ( .A(n3190), .Y(n4329) );
  INVX1_LVT U4297 ( .A(n3092), .Y(n4355) );
  INVX1_LVT U4298 ( .A(n3193), .Y(n4352) );
  AND2X1_LVT U4299 ( .A1(n5434), .A2(n6238), .Y(n6877) );
  INVX1_LVT U4300 ( .A(n3189), .Y(n4343) );
  INVX1_LVT U4301 ( .A(n3099), .Y(n4402) );
  INVX1_LVT U4302 ( .A(n3091), .Y(n4407) );
  IBUFFX2_LVT U4303 ( .A(n6238), .Y(n6898) );
  INVX1_LVT U4304 ( .A(n3090), .Y(n4394) );
  INVX1_LVT U4305 ( .A(n3193), .Y(n4353) );
  INVX1_LVT U4306 ( .A(n3183), .Y(n4412) );
  XOR2X1_LVT U4307 ( .A1(n9485), .A2(ibuf_io_pc[6]), .Y(n4546) );
  INVX1_LVT U4308 ( .A(n3192), .Y(n4341) );
  INVX1_LVT U4309 ( .A(n3190), .Y(n4328) );
  INVX1_LVT U4310 ( .A(n3189), .Y(n4344) );
  INVX1_LVT U4311 ( .A(n3186), .Y(n4350) );
  INVX1_LVT U4312 ( .A(n3196), .Y(n4323) );
  AOI21X1_LVT U4313 ( .A1(n3842), .A2(csr_io_rw_rdata[13]), .A3(n5707), .Y(
        n3092) );
  INVX1_LVT U4314 ( .A(n3187), .Y(n4326) );
  INVX1_LVT U4315 ( .A(n3197), .Y(n4332) );
  INVX1_LVT U4316 ( .A(n3194), .Y(n4335) );
  INVX1_LVT U4317 ( .A(n3191), .Y(n4338) );
  NOR2X1_LVT U4318 ( .A1(csr_io_interrupt), .A2(ibuf_io_inst_0_bits_replay), 
        .Y(n9385) );
  AOI21X1_LVT U4319 ( .A1(n3842), .A2(csr_io_rw_rdata[12]), .A3(n5683), .Y(
        n3193) );
  AOI21X1_LVT U4320 ( .A1(n3843), .A2(csr_io_rw_rdata[28]), .A3(n6014), .Y(
        n3090) );
  INVX1_LVT U4321 ( .A(n3187), .Y(n4327) );
  INVX1_LVT U4322 ( .A(n3196), .Y(n4322) );
  INVX1_LVT U4323 ( .A(ibuf_io_inst_0_bits_inst_rs1[4]), .Y(n6963) );
  INVX1_LVT U4324 ( .A(n3197), .Y(n4331) );
  INVX1_LVT U4325 ( .A(n3094), .Y(n4379) );
  INVX1_LVT U4326 ( .A(n3191), .Y(n4339) );
  INVX1_LVT U4327 ( .A(n3096), .Y(n4389) );
  AOI21X1_LVT U4328 ( .A1(n3843), .A2(csr_io_rw_rdata[31]), .A3(n6083), .Y(
        n3099) );
  AOI21X1_LVT U4329 ( .A1(n3842), .A2(csr_io_rw_rdata[9]), .A3(n5628), .Y(
        n3189) );
  INVX1_LVT U4330 ( .A(n3196), .Y(n4324) );
  AOI21X1_LVT U4331 ( .A1(n3842), .A2(csr_io_rw_rdata[8]), .A3(n5604), .Y(
        n3192) );
  INVX1_LVT U4332 ( .A(n3197), .Y(n4333) );
  INVX1_LVT U4333 ( .A(n3187), .Y(n4325) );
  INVX1_LVT U4334 ( .A(n3194), .Y(n4334) );
  INVX1_LVT U4335 ( .A(csr_io_interrupt), .Y(n9448) );
  INVX1_LVT U4336 ( .A(n3191), .Y(n4337) );
  INVX1_LVT U4337 ( .A(n3194), .Y(n4336) );
  INVX1_LVT U4338 ( .A(n3093), .Y(n4360) );
  INVX1_LVT U4339 ( .A(n3186), .Y(n4349) );
  OR2X1_LVT U4340 ( .A1(csr_io_status_isa[3]), .A2(n3583), .Y(n3570) );
  AOI21X1_LVT U4341 ( .A1(n3841), .A2(csr_io_rw_rdata[7]), .A3(n5584), .Y(
        n3191) );
  AOI21X1_LVT U4342 ( .A1(n3841), .A2(csr_io_rw_rdata[3]), .A3(n5505), .Y(
        n3187) );
  INVX1_LVT U4343 ( .A(n3188), .Y(n4348) );
  INVX0_LVT U4344 ( .A(n9525), .Y(n5067) );
  AOI21X1_LVT U4345 ( .A1(n3841), .A2(csr_io_rw_rdata[6]), .A3(n5560), .Y(
        n3194) );
  IBUFFX2_LVT U4346 ( .A(n5075), .Y(n2571) );
  INVX1_LVT U4347 ( .A(n3083), .Y(n3863) );
  NBUFFX2_LVT U4348 ( .A(n6794), .Y(n3811) );
  AOI21X1_LVT U4349 ( .A1(n3843), .A2(csr_io_rw_rdata[15]), .A3(n5746), .Y(
        n3093) );
  AOI21X1_LVT U4350 ( .A1(n3843), .A2(csr_io_rw_rdata[26]), .A3(n5973), .Y(
        n3096) );
  INVX1_LVT U4351 ( .A(n3188), .Y(n4346) );
  INVX1_LVT U4352 ( .A(n3188), .Y(n4347) );
  AOI21X1_LVT U4353 ( .A1(n3841), .A2(csr_io_rw_rdata[2]), .A3(n5486), .Y(
        n3196) );
  AOI21X1_LVT U4354 ( .A1(n3841), .A2(csr_io_rw_rdata[5]), .A3(n5536), .Y(
        n3197) );
  INVX1_LVT U4355 ( .A(n3095), .Y(n4377) );
  INVX1_LVT U4356 ( .A(n3098), .Y(n4420) );
  AND2X1_LVT U4357 ( .A1(n4890), .A2(n4816), .Y(n5456) );
  INVX1_LVT U4358 ( .A(n5435), .Y(n5455) );
  AOI21X1_LVT U4359 ( .A1(n3844), .A2(csr_io_rw_rdata[21]), .A3(n5863), .Y(
        n3095) );
  AOI21X1_LVT U4360 ( .A1(n3842), .A2(csr_io_rw_rdata[10]), .A3(n5652), .Y(
        n3188) );
  NBUFFX2_LVT U4361 ( .A(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(n3781) );
  OR2X1_LVT U4362 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n4814), .Y(n5435) );
  AOI21X1_LVT U4363 ( .A1(n3842), .A2(csr_io_rw_rdata[38]), .A3(n6232), .Y(
        n3098) );
  AND2X1_LVT U4364 ( .A1(n4889), .A2(n4816), .Y(n5452) );
  AND2X1_LVT U4365 ( .A1(n4900), .A2(n4816), .Y(n5454) );
  NOR2X0_LVT U4366 ( .A1(wb_reg_flush_pipe), .A2(n9332), .Y(
        io_imem_req_bits_speculative) );
  NOR2X1_LVT U4367 ( .A1(n_T_726[1]), .A2(n_T_726[0]), .Y(n9430) );
  NAND4X0_LVT U4368 ( .A1(n4870), .A2(n4869), .A3(n3046), .A4(n4868), .Y(n4888) );
  AND2X1_LVT U4369 ( .A1(n9387), .A2(n9388), .Y(n9394) );
  NOR2X1_LVT U4370 ( .A1(n9400), .A2(n9402), .Y(n9401) );
  NOR2X1_LVT U4371 ( .A1(n9331), .A2(n4065), .Y(n9414) );
  NOR2X0_LVT U4372 ( .A1(n9403), .A2(n9402), .Y(n9410) );
  OR2X1_LVT U4373 ( .A1(n5359), .A2(n5358), .Y(n5393) );
  NOR2X1_LVT U4374 ( .A1(n5362), .A2(n5358), .Y(n5378) );
  OR2X1_LVT U4375 ( .A1(n5327), .A2(n5358), .Y(n5334) );
  NOR2X1_LVT U4376 ( .A1(n5381), .A2(n5358), .Y(n5366) );
  NOR2X1_LVT U4377 ( .A1(n5365), .A2(n5358), .Y(n5383) );
  NAND2X0_LVT U4378 ( .A1(n9380), .A2(n4498), .Y(n5358) );
  AO21X1_LVT U4379 ( .A1(n9103), .A2(io_fpu_fromint_data[43]), .A3(n9102), .Y(
        alu_io_in1[43]) );
  AO21X1_LVT U4380 ( .A1(n9103), .A2(io_fpu_fromint_data[41]), .A3(n9102), .Y(
        alu_io_in1[41]) );
  NOR2X1_LVT U4381 ( .A1(n5365), .A2(n5254), .Y(n5275) );
  AO22X1_LVT U4382 ( .A1(n_T_698[27]), .A2(n9101), .A3(io_fpu_fromint_data[27]), .A4(n9103), .Y(alu_io_in1[27]) );
  AO22X1_LVT U4383 ( .A1(n_T_698[28]), .A2(n9101), .A3(io_fpu_fromint_data[28]), .A4(n9103), .Y(alu_io_in1[28]) );
  AO21X1_LVT U4384 ( .A1(n9103), .A2(io_fpu_fromint_data[55]), .A3(n9102), .Y(
        alu_io_in1[55]) );
  NOR2X1_LVT U4385 ( .A1(n5381), .A2(n5254), .Y(n5265) );
  AO22X1_LVT U4386 ( .A1(n_T_698[25]), .A2(n9101), .A3(io_fpu_fromint_data[25]), .A4(n9103), .Y(alu_io_in1[25]) );
  AO21X1_LVT U4387 ( .A1(n9103), .A2(io_fpu_fromint_data[51]), .A3(n9102), .Y(
        alu_io_in1[51]) );
  AO22X1_LVT U4388 ( .A1(n4054), .A2(n_T_698[26]), .A3(io_fpu_fromint_data[26]), .A4(n9103), .Y(alu_io_in1[26]) );
  AO21X1_LVT U4389 ( .A1(n9103), .A2(io_fpu_fromint_data[49]), .A3(n9102), .Y(
        alu_io_in1[49]) );
  AO22X1_LVT U4390 ( .A1(n9101), .A2(n_T_698[11]), .A3(io_fpu_fromint_data[11]), .A4(n9103), .Y(alu_io_in1[11]) );
  AO21X1_LVT U4391 ( .A1(n9103), .A2(io_fpu_fromint_data[39]), .A3(n9102), .Y(
        alu_io_in1[39]) );
  AO22X1_LVT U4392 ( .A1(n_T_698[8]), .A2(n4054), .A3(io_fpu_fromint_data[8]), 
        .A4(n9103), .Y(alu_io_in1[8]) );
  AO22X1_LVT U4393 ( .A1(n_T_698[9]), .A2(n4054), .A3(io_fpu_fromint_data[9]), 
        .A4(n9103), .Y(alu_io_in1[9]) );
  AO22X1_LVT U4394 ( .A1(n9101), .A2(n_T_698[5]), .A3(io_fpu_fromint_data[5]), 
        .A4(n9103), .Y(alu_io_in1[5]) );
  NOR2X1_LVT U4395 ( .A1(n5362), .A2(n5254), .Y(n5285) );
  AO21X1_LVT U4396 ( .A1(n9103), .A2(io_fpu_fromint_data[63]), .A3(n9102), .Y(
        alu_io_in1[63]) );
  AND3X1_LVT U4397 ( .A1(n9400), .A2(n9398), .A3(n9397), .Y(n9396) );
  AO22X1_LVT U4398 ( .A1(n_T_698[31]), .A2(n9101), .A3(io_fpu_fromint_data[31]), .A4(n9103), .Y(alu_io_in1[31]) );
  NOR2X1_LVT U4399 ( .A1(n5392), .A2(n5254), .Y(n5248) );
  OR2X1_LVT U4400 ( .A1(n7905), .A2(n7904), .Y(io_fpu_fromint_data[31]) );
  NAND2X0_LVT U4401 ( .A1(csr_io_retire), .A2(n5176), .Y(n5254) );
  INVX0_LVT U4402 ( .A(ibuf_io_inst_0_bits_raw[1]), .Y(n3646) );
  IBUFFX2_LVT U4403 ( .A(n3042), .Y(n2573) );
  NOR3X1_LVT U4404 ( .A1(n3203), .A2(n9330), .A3(csr_io_exception), .Y(
        csr_io_retire) );
  IBUFFX2_LVT U4405 ( .A(n3040), .Y(n2574) );
  MUX21X1_LVT U4406 ( .A1(wb_reg_cause[1]), .A2(n9251), .S0(n576), .Y(
        wb_cause[1]) );
  NOR2X1_LVT U4407 ( .A1(n_T_728[1]), .A2(n_T_728[0]), .Y(n9118) );
  OR2X1_LVT U4408 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(
        ibuf_io_inst_0_bits_raw[28]), .Y(n4804) );
  NOR2X0_LVT U4409 ( .A1(n6860), .A2(n5415), .Y(n6861) );
  NOR2X1_LVT U4410 ( .A1(mem_ctrl_jalr), .A2(mem_reg_sfence), .Y(n4591) );
  NOR2X1_LVT U4411 ( .A1(n5426), .A2(n5428), .Y(n5314) );
  INVX0_LVT U4412 ( .A(ibuf_io_inst_0_bits_raw[28]), .Y(n4782) );
  AND3X1_LVT U4413 ( .A1(n7019), .A2(n3101), .A3(n3255), .Y(n9066) );
  OR2X1_LVT U4414 ( .A1(io_dmem_s2_nack), .A2(wb_reg_replay), .Y(n9330) );
  NBUFFX2_LVT U4415 ( .A(net34480), .Y(n4285) );
  INVX1_LVT U4416 ( .A(n3784), .Y(n3785) );
  INVX1_LVT U4417 ( .A(io_fpu_dmem_resp_tag[4]), .Y(n5228) );
  AND2X1_LVT U4418 ( .A1(io_dmem_resp_valid), .A2(io_dmem_resp_bits_has_data), 
        .Y(n2626) );
  INVX1_LVT U4419 ( .A(io_fpu_dmem_resp_tag[1]), .Y(n5185) );
  INVX0_LVT U4420 ( .A(io_dmem_perf_grant), .Y(n5065) );
  INVX1_LVT U4421 ( .A(io_fpu_dmem_resp_tag[3]), .Y(n5249) );
  INVX0_LVT U4422 ( .A(io_fpu_fcsr_rdy), .Y(n4918) );
  INVX0_LVT U4423 ( .A(io_dmem_req_ready), .Y(n5064) );
  OR2X1_LVT U4424 ( .A1(io_fpu_dmem_resp_tag[3]), .A2(io_fpu_dmem_resp_tag[4]), 
        .Y(n5192) );
  NAND3X0_LVT U4425 ( .A1(n8870), .A2(n8868), .A3(n2577), .Y(n8871) );
  OA21X1_LVT U4426 ( .A1(n4011), .A2(n3368), .A3(n8869), .Y(n2577) );
  OA21X1_LVT U4427 ( .A1(n4012), .A2(n3356), .A3(n8618), .Y(n2578) );
  OA21X1_LVT U4428 ( .A1(n4012), .A2(n3347), .A3(n8451), .Y(n2579) );
  OA21X1_LVT U4429 ( .A1(n4013), .A2(n3350), .A3(n8515), .Y(n2580) );
  NAND2X0_LVT U4430 ( .A1(n_T_427[490]), .A2(n3614), .Y(n8264) );
  IBUFFX2_LVT U4431 ( .A(n3663), .Y(n2611) );
  NAND4X0_LVT U4432 ( .A1(n3662), .A2(n3780), .A3(n2910), .A4(n2581), .Y(N735)
         );
  NOR3X0_LVT U4433 ( .A1(n2582), .A2(n8888), .A3(n8889), .Y(n3730) );
  AND3X1_LVT U4434 ( .A1(n7355), .A2(n7356), .A3(n2583), .Y(n2958) );
  OA21X1_LVT U4435 ( .A1(n3439), .A2(n4008), .A3(n7357), .Y(n2583) );
  AND3X1_LVT U4436 ( .A1(n2935), .A2(n7271), .A3(n7272), .Y(n2584) );
  AND3X1_LVT U4437 ( .A1(n7937), .A2(n7936), .A3(n7938), .Y(n2585) );
  NAND2X0_LVT U4438 ( .A1(n_T_427[486]), .A2(n3614), .Y(n8125) );
  IBUFFX2_LVT U4439 ( .A(n2984), .Y(n4012) );
  OR2X1_LVT U4440 ( .A1(n3427), .A2(n3653), .Y(n2586) );
  NAND2X0_LVT U4441 ( .A1(n2611), .A2(n_T_427[1155]), .Y(n2587) );
  NAND2X0_LVT U4442 ( .A1(n_T_427[1219]), .A2(n3638), .Y(n2588) );
  OR3X2_LVT U4443 ( .A1(io_fpu_inst[4]), .A2(n3593), .A3(n9528), .Y(n9113) );
  NAND2X0_LVT U4444 ( .A1(n_T_427[303]), .A2(n3790), .Y(n2589) );
  AND2X1_LVT U4445 ( .A1(n8218), .A2(n8219), .Y(n2602) );
  NAND2X0_LVT U4446 ( .A1(n_T_427[498]), .A2(n3614), .Y(n8550) );
  AND4X1_LVT U4447 ( .A1(n8099), .A2(n8100), .A3(n8098), .A4(n8097), .Y(n2950)
         );
  NAND2X0_LVT U4448 ( .A1(n_T_427[480]), .A2(n3614), .Y(n7923) );
  AND2X1_LVT U4449 ( .A1(n8349), .A2(n8348), .Y(n2590) );
  AND4X1_LVT U4450 ( .A1(n7958), .A2(n7957), .A3(n7956), .A4(n7955), .Y(n2963)
         );
  NAND2X0_LVT U4451 ( .A1(n_T_427[312]), .A2(n3790), .Y(n2591) );
  NAND2X0_LVT U4452 ( .A1(n_T_427[1431]), .A2(n3629), .Y(n2592) );
  AND3X1_LVT U4453 ( .A1(n2594), .A2(n8961), .A3(n3050), .Y(n2987) );
  AND2X1_LVT U4454 ( .A1(n8962), .A2(n8960), .Y(n2594) );
  AOI21X1_LVT U4455 ( .A1(n9429), .A2(n9107), .A3(n9445), .Y(n2657) );
  NAND2X0_LVT U4456 ( .A1(n2596), .A2(n2646), .Y(n4513) );
  NOR4X1_LVT U4457 ( .A1(n4501), .A2(n9437), .A3(n2606), .A4(n4500), .Y(n2596)
         );
  OR2X1_LVT U4458 ( .A1(n3191), .A2(n2089), .Y(n2597) );
  AND2X1_LVT U4459 ( .A1(n3960), .A2(n8105), .Y(n9052) );
  AND2X1_LVT U4460 ( .A1(n8631), .A2(n2598), .Y(n2617) );
  DELLN1X2_LVT U4461 ( .A(n9052), .Y(n3614) );
  AND2X1_LVT U4462 ( .A1(n3678), .A2(n2599), .Y(n2910) );
  AND3X1_LVT U4463 ( .A1(n8739), .A2(n8738), .A3(n8740), .Y(n2599) );
  NOR3X0_LVT U4464 ( .A1(n2601), .A2(n8222), .A3(n8221), .Y(n3746) );
  OA21X1_LVT U4465 ( .A1(n4011), .A2(n3344), .A3(n8383), .Y(n2604) );
  OA21X1_LVT U4466 ( .A1(n4012), .A2(n3300), .A3(n8418), .Y(n2605) );
  OR2X1_LVT U4467 ( .A1(io_fpu_inst[7]), .A2(io_fpu_inst[26]), .Y(n2606) );
  NAND4X0_LVT U4468 ( .A1(n9032), .A2(n9027), .A3(n9031), .A4(n2607), .Y(n9033) );
  NAND4X0_LVT U4469 ( .A1(n8204), .A2(n8202), .A3(n8203), .A4(n2609), .Y(n8205) );
  OR2X1_LVT U4470 ( .A1(n3338), .A2(n4013), .Y(n2609) );
  NAND2X0_LVT U4471 ( .A1(n_T_427[1457]), .A2(n3627), .Y(n8562) );
  OA21X1_LVT U4472 ( .A1(n3752), .A2(n3282), .A3(n7426), .Y(n2610) );
  IBUFFX2_LVT U4473 ( .A(n3768), .Y(n3664) );
  IBUFFX2_LVT U4474 ( .A(n3768), .Y(n4008) );
  IBUFFX2_LVT U4475 ( .A(n3768), .Y(n4009) );
  AOI22X1_LVT U4476 ( .A1(n4330), .A2(n2982), .A3(n2966), .A4(n_T_427[1411]), 
        .Y(n7105) );
  OR2X1_LVT U4477 ( .A1(n3459), .A2(n3658), .Y(n2612) );
  NAND4X0_LVT U4478 ( .A1(n8074), .A2(n8076), .A3(n8075), .A4(n2613), .Y(n8077) );
  OR2X1_LVT U4479 ( .A1(n3455), .A2(n3658), .Y(n2613) );
  OR2X1_LVT U4480 ( .A1(n3403), .A2(n3658), .Y(n2614) );
  AND2X1_LVT U4481 ( .A1(n9446), .A2(n2616), .Y(n2615) );
  NBUFFX2_LVT U4482 ( .A(io_fpu_inst[12]), .Y(n2618) );
  IBUFFX2_LVT U4483 ( .A(n3683), .Y(n3631) );
  IBUFFX2_LVT U4484 ( .A(n9527), .Y(n3783) );
  NAND2X0_LVT U4485 ( .A1(n9438), .A2(n5144), .Y(n2620) );
  AND2X1_LVT U4486 ( .A1(n2544), .A2(n6906), .Y(n2621) );
  OA21X1_LVT U4487 ( .A1(n4010), .A2(n3428), .A3(n7190), .Y(n2622) );
  OA21X1_LVT U4488 ( .A1(n2643), .A2(n2639), .A3(n2640), .Y(n2624) );
  XNOR2X1_LVT U4489 ( .A1(n3782), .A2(n589), .Y(n2625) );
  OR2X2_LVT U4490 ( .A1(n5036), .A2(n5013), .Y(n6992) );
  INVX1_LVT U4491 ( .A(n6931), .Y(n6947) );
  NAND2X0_LVT U4492 ( .A1(n6956), .A2(n6931), .Y(n4040) );
  AND2X1_LVT U4493 ( .A1(n2038), .A2(n4970), .Y(n6931) );
  MUX21X1_LVT U4494 ( .A1(n3043), .A2(n5313), .S0(n9381), .Y(n3042) );
  MUX21X1_LVT U4495 ( .A1(io_fpu_dmem_resp_tag[2]), .A2(
        div_io_resp_bits_tag[2]), .S0(n5403), .Y(n5313) );
  NAND2X0_LVT U4496 ( .A1(n2153), .A2(n4685), .Y(n5413) );
  AND3X1_LVT U4497 ( .A1(n5124), .A2(n2628), .A3(n2627), .Y(n6939) );
  NAND2X0_LVT U4498 ( .A1(n5122), .A2(n3049), .Y(n6916) );
  OA21X1_LVT U4499 ( .A1(n3072), .A2(n5123), .A3(
        csr_io_decode_0_system_illegal), .Y(n6915) );
  OR2X1_LVT U4500 ( .A1(csr_io_status_isa[2]), .A2(n4497), .Y(n2628) );
  AND2X1_LVT U4501 ( .A1(n5106), .A2(n5105), .Y(n2630) );
  AND2X1_LVT U4502 ( .A1(n2631), .A2(n2658), .Y(n2633) );
  OA22X1_LVT U4503 ( .A1(n2635), .A2(n2636), .A3(n5098), .A4(n2634), .Y(n2631)
         );
  AND4X1_LVT U4504 ( .A1(n5104), .A2(n5103), .A3(n9445), .A4(n2632), .Y(n2637)
         );
  NAND2X0_LVT U4505 ( .A1(n3635), .A2(n_T_427[1271]), .Y(n2638) );
  OA21X1_LVT U4506 ( .A1(n5135), .A2(n5134), .A3(n5140), .Y(n2640) );
  OR2X1_LVT U4507 ( .A1(n3656), .A2(n8521), .Y(n8522) );
  AO21X1_LVT U4508 ( .A1(n7321), .A2(n7322), .A3(n2154), .Y(n7323) );
  AO21X1_LVT U4509 ( .A1(n7377), .A2(n7378), .A3(n3632), .Y(n7379) );
  AO21X1_LVT U4510 ( .A1(n7779), .A2(n7780), .A3(n2645), .Y(n7781) );
  AO21X1_LVT U4511 ( .A1(n7811), .A2(n7812), .A3(n2154), .Y(n7813) );
  AO21X1_LVT U4512 ( .A1(n7747), .A2(n7748), .A3(n2155), .Y(n7749) );
  AO21X1_LVT U4513 ( .A1(n7871), .A2(n7872), .A3(n3656), .Y(n7873) );
  AND2X1_LVT U4514 ( .A1(n4503), .A2(n4502), .Y(n2646) );
  AND2X1_LVT U4515 ( .A1(n3577), .A2(n9439), .Y(n2647) );
  AND2X1_LVT U4516 ( .A1(n3077), .A2(n3577), .Y(n2648) );
  AND2X1_LVT U4517 ( .A1(io_fpu_inst[3]), .A2(n5163), .Y(n9428) );
  NAND2X0_LVT U4518 ( .A1(n3577), .A2(n5067), .Y(n9095) );
  AND3X1_LVT U4519 ( .A1(n6966), .A2(n6917), .A3(n6946), .Y(n2650) );
  AND4X1_LVT U4520 ( .A1(n2652), .A2(n7455), .A3(n2653), .A4(n3697), .Y(n2651)
         );
  AND2X1_LVT U4521 ( .A1(n7456), .A2(n7457), .Y(n2652) );
  OR2X1_LVT U4522 ( .A1(n3139), .A2(n3987), .Y(n2653) );
  AND4X1_LVT U4523 ( .A1(n3706), .A2(n2656), .A3(n7576), .A4(n2654), .Y(n2655)
         );
  AND2X1_LVT U4524 ( .A1(n7577), .A2(n7578), .Y(n2654) );
  AND2X1_LVT U4525 ( .A1(n5102), .A2(n9104), .Y(n9429) );
  NAND2X0_LVT U4526 ( .A1(n3991), .A2(n_T_427[1903]), .Y(n2660) );
  AND3X1_LVT U4527 ( .A1(n3701), .A2(n3702), .A3(n2659), .Y(n3028) );
  AND4X1_LVT U4528 ( .A1(n7609), .A2(n7608), .A3(n2661), .A4(n2660), .Y(n2659)
         );
  NAND2X0_LVT U4529 ( .A1(n2882), .A2(n_T_427[1901]), .Y(n2663) );
  AND4X1_LVT U4530 ( .A1(n3703), .A2(n3704), .A3(n7546), .A4(n2662), .Y(n3017)
         );
  NAND3X0_LVT U4531 ( .A1(n3006), .A2(n2666), .A3(n2665), .Y(N710) );
  AND4X1_LVT U4532 ( .A1(n3005), .A2(n3065), .A3(n3064), .A4(n2668), .Y(n2665)
         );
  AND2X1_LVT U4533 ( .A1(n2667), .A2(n7860), .Y(n2666) );
  AND2X1_LVT U4534 ( .A1(n7861), .A2(n7862), .Y(n2667) );
  AND2X1_LVT U4535 ( .A1(n3180), .A2(n3580), .Y(n2670) );
  AND2X1_LVT U4536 ( .A1(n3765), .A2(n2561), .Y(n6941) );
  AND2X1_LVT U4537 ( .A1(n2143), .A2(n2672), .Y(n2671) );
  AND2X1_LVT U4538 ( .A1(n6917), .A2(n6954), .Y(n2672) );
  XOR2X1_LVT U4539 ( .A1(n2876), .A2(n591), .Y(n5037) );
  NAND2X0_LVT U4540 ( .A1(n2673), .A2(n2538), .Y(n5094) );
  AOI21X1_LVT U4541 ( .A1(n2676), .A2(n9116), .A3(n2675), .Y(N279) );
  INVX1_LVT U4542 ( .A(n4732), .Y(n4675) );
  AND2X1_LVT U4543 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(
        ibuf_io_inst_0_bits_inst_rd[0]), .Y(n4730) );
  AOI21X1_LVT U4544 ( .A1(n9281), .A2(n3048), .A3(n9280), .Y(n9283) );
  AOI22X1_LVT U4545 ( .A1(n3903), .A2(n_T_427[721]), .A3(n_T_427[17]), .A4(
        n3914), .Y(n2680) );
  AOI22X1_LVT U4546 ( .A1(n3908), .A2(n_T_427[149]), .A3(n_T_427[277]), .A4(
        n2828), .Y(n2844) );
  AOI22X1_LVT U4547 ( .A1(n2864), .A2(n_T_427[401]), .A3(n_T_427[1040]), .A4(
        n3898), .Y(n2678) );
  AND4X1_LVT U4548 ( .A1(n2678), .A2(n2679), .A3(n2680), .A4(n2681), .Y(n5794)
         );
  AND2X1_LVT U4549 ( .A1(n2682), .A2(n2683), .Y(n5895) );
  AOI22X1_LVT U4550 ( .A1(n3902), .A2(n_T_427[1080]), .A3(n_T_427[249]), .A4(
        n3808), .Y(n2744) );
  OA22X1_LVT U4551 ( .A1(n3371), .A2(n3080), .A3(n3881), .A4(n2684), .Y(n2775)
         );
  AND2X1_LVT U4552 ( .A1(n2685), .A2(n2686), .Y(n6132) );
  AOI22X1_LVT U4553 ( .A1(n3833), .A2(n_T_427[97]), .A3(n_T_427[225]), .A4(
        n3806), .Y(n2685) );
  AOI22X1_LVT U4554 ( .A1(n2831), .A2(n_T_427[928]), .A3(n_T_427[161]), .A4(
        n2862), .Y(n2686) );
  AOI22X1_LVT U4555 ( .A1(n3900), .A2(n_T_427[1055]), .A3(n_T_427[224]), .A4(
        n3808), .Y(n2687) );
  AOI22X1_LVT U4556 ( .A1(n2870), .A2(n_T_427[608]), .A3(n_T_427[32]), .A4(
        n2879), .Y(n2688) );
  AOI22X1_LVT U4557 ( .A1(n3819), .A2(n_T_427[544]), .A3(n_T_427[863]), .A4(
        n3823), .Y(n2689) );
  AND4X1_LVT U4558 ( .A1(n2690), .A2(n2691), .A3(n2692), .A4(n2693), .Y(n6628)
         );
  AOI22X1_LVT U4559 ( .A1(n3902), .A2(n_T_427[1077]), .A3(n_T_427[949]), .A4(
        n3895), .Y(n2692) );
  AOI22X1_LVT U4560 ( .A1(n3906), .A2(n_T_427[821]), .A3(n_T_427[438]), .A4(
        n2865), .Y(n2693) );
  AND4X1_LVT U4561 ( .A1(n2694), .A2(n2695), .A3(n2696), .A4(n2697), .Y(n6362)
         );
  AOI22X1_LVT U4562 ( .A1(n3901), .A2(n_T_427[1066]), .A3(n_T_427[938]), .A4(
        n3896), .Y(n2696) );
  AND4X1_LVT U4563 ( .A1(n2698), .A2(n2699), .A3(n2700), .A4(n2701), .Y(n6506)
         );
  AOI22X1_LVT U4564 ( .A1(n3901), .A2(n_T_427[1072]), .A3(n_T_427[113]), .A4(
        n3833), .Y(n2700) );
  AOI22X1_LVT U4565 ( .A1(n3910), .A2(n_T_427[497]), .A3(n_T_427[752]), .A4(
        n2827), .Y(n2701) );
  AND4X1_LVT U4566 ( .A1(n2702), .A2(n2703), .A3(n2704), .A4(n2705), .Y(n6680)
         );
  AOI22X1_LVT U4567 ( .A1(n3902), .A2(n_T_427[1079]), .A3(n_T_427[951]), .A4(
        n3897), .Y(n2704) );
  AOI22X1_LVT U4568 ( .A1(n3835), .A2(n_T_427[440]), .A3(n_T_427[184]), .A4(
        n2863), .Y(n2705) );
  AOI22X1_LVT U4569 ( .A1(n2856), .A2(n_T_427[351]), .A3(n_T_427[95]), .A4(
        n3831), .Y(n2847) );
  AND4X1_LVT U4570 ( .A1(n2706), .A2(n2707), .A3(n2708), .A4(n2709), .Y(n6408)
         );
  AND4X1_LVT U4571 ( .A1(n2710), .A2(n2711), .A3(n2712), .A4(n2713), .Y(n6555)
         );
  AOI22X1_LVT U4572 ( .A1(n3902), .A2(n_T_427[1074]), .A3(n_T_427[243]), .A4(
        n2830), .Y(n2712) );
  AOI22X1_LVT U4573 ( .A1(n2832), .A2(n_T_427[946]), .A3(n_T_427[754]), .A4(
        n2827), .Y(n2713) );
  AND4X1_LVT U4574 ( .A1(n2714), .A2(n2715), .A3(n2716), .A4(n2717), .Y(n6224)
         );
  AOI22X1_LVT U4575 ( .A1(n3944), .A2(n_T_427[1188]), .A3(n_T_427[1252]), .A4(
        n3939), .Y(n2714) );
  AOI22X1_LVT U4576 ( .A1(n3954), .A2(n_T_427[1124]), .A3(n_T_427[996]), .A4(
        n3949), .Y(n2715) );
  AOI22X1_LVT U4577 ( .A1(n3901), .A2(n_T_427[1060]), .A3(n_T_427[229]), .A4(
        n3807), .Y(n2716) );
  AOI22X1_LVT U4578 ( .A1(n3832), .A2(n_T_427[101]), .A3(n_T_427[740]), .A4(
        n6884), .Y(n2717) );
  AND4X1_LVT U4579 ( .A1(n2718), .A2(n2719), .A3(n2720), .A4(n2721), .Y(n6291)
         );
  AOI22X1_LVT U4580 ( .A1(n3901), .A2(n_T_427[1063]), .A3(n_T_427[232]), .A4(
        n3808), .Y(n2720) );
  AOI22X1_LVT U4581 ( .A1(n3833), .A2(n_T_427[104]), .A3(n_T_427[935]), .A4(
        n3896), .Y(n2721) );
  AND4X1_LVT U4582 ( .A1(n2722), .A2(n2723), .A3(n2724), .A4(n2725), .Y(n6482)
         );
  AOI22X1_LVT U4583 ( .A1(n3901), .A2(n_T_427[1071]), .A3(n_T_427[240]), .A4(
        n3807), .Y(n2724) );
  AOI22X1_LVT U4584 ( .A1(n3834), .A2(n_T_427[432]), .A3(n_T_427[943]), .A4(
        n2832), .Y(n2725) );
  AND4X1_LVT U4585 ( .A1(n2726), .A2(n2727), .A3(n2728), .A4(n2729), .Y(n5601)
         );
  AOI22X1_LVT U4586 ( .A1(n3943), .A2(n_T_427[1158]), .A3(n_T_427[1222]), .A4(
        n3937), .Y(n2726) );
  AOI22X1_LVT U4587 ( .A1(n3953), .A2(n_T_427[1094]), .A3(n_T_427[966]), .A4(
        n3947), .Y(n2727) );
  AOI22X1_LVT U4588 ( .A1(n3899), .A2(n_T_427[1030]), .A3(n_T_427[199]), .A4(
        n3808), .Y(n2728) );
  AND4X1_LVT U4589 ( .A1(n2730), .A2(n2731), .A3(n2732), .A4(n2733), .Y(n6726)
         );
  AND4X1_LVT U4590 ( .A1(n2734), .A2(n2735), .A3(n2736), .A4(n2737), .Y(n6457)
         );
  AND4X1_LVT U4591 ( .A1(n2738), .A2(n2739), .A3(n2740), .A4(n2741), .Y(n6203)
         );
  AOI22X1_LVT U4592 ( .A1(n3944), .A2(n_T_427[1187]), .A3(n_T_427[1251]), .A4(
        n3939), .Y(n2738) );
  AOI22X1_LVT U4593 ( .A1(n3954), .A2(n_T_427[1123]), .A3(n_T_427[995]), .A4(
        n3949), .Y(n2739) );
  AND4X1_LVT U4594 ( .A1(n2742), .A2(n2743), .A3(n2744), .A4(n2745), .Y(n6701)
         );
  AOI22X1_LVT U4595 ( .A1(n3831), .A2(n_T_427[121]), .A3(n_T_427[760]), .A4(
        n3905), .Y(n2745) );
  IBUFFX2_LVT U4596 ( .A(n6878), .Y(n3884) );
  AND4X1_LVT U4597 ( .A1(n2746), .A2(n2747), .A3(n2748), .A4(n2749), .Y(n6184)
         );
  AOI22X1_LVT U4598 ( .A1(n2028), .A2(n_T_427[1876]), .A3(n3884), .A4(
        n_T_427[1915]), .Y(n2747) );
  AOI22X1_LVT U4599 ( .A1(n3827), .A2(n_T_427[1698]), .A3(n_T_427[1570]), .A4(
        n3890), .Y(n2748) );
  AOI22X1_LVT U4600 ( .A1(n3889), .A2(n_T_427[1634]), .A3(n_T_427[1506]), .A4(
        n3922), .Y(n2749) );
  AOI22X1_LVT U4601 ( .A1(n2028), .A2(n_T_427[1857]), .A3(n3884), .A4(
        n_T_427[1892]), .Y(n2750) );
  AND4X1_LVT U4602 ( .A1(n2751), .A2(n2752), .A3(n2753), .A4(n2754), .Y(n6134)
         );
  AOI22X1_LVT U4603 ( .A1(n3801), .A2(n_T_427[1874]), .A3(n3884), .A4(
        n_T_427[1913]), .Y(n2752) );
  AOI22X1_LVT U4604 ( .A1(n3827), .A2(n_T_427[1696]), .A3(n_T_427[1568]), .A4(
        n3890), .Y(n2753) );
  AOI22X1_LVT U4605 ( .A1(n3889), .A2(n_T_427[1632]), .A3(n_T_427[1504]), .A4(
        n3922), .Y(n2754) );
  AOI22X1_LVT U4606 ( .A1(n6764), .A2(n_T_427[1862]), .A3(n_T_427[1743]), .A4(
        n3798), .Y(n2755) );
  AND4X1_LVT U4607 ( .A1(n2757), .A2(n2758), .A3(n2759), .A4(n2760), .Y(n6270)
         );
  AOI22X1_LVT U4608 ( .A1(n3801), .A2(n_T_427[1878]), .A3(n_T_427[1766]), .A4(
        n2867), .Y(n2757) );
  AOI22X1_LVT U4609 ( .A1(n2765), .A2(n_T_427[1827]), .A3(n_T_427[1702]), .A4(
        n3825), .Y(n2758) );
  AOI22X1_LVT U4610 ( .A1(n3892), .A2(n_T_427[1574]), .A3(n_T_427[1638]), .A4(
        n3887), .Y(n2759) );
  AND4X1_LVT U4611 ( .A1(n2761), .A2(n2762), .A3(n2763), .A4(n2764), .Y(n6388)
         );
  AOI22X1_LVT U4612 ( .A1(n6764), .A2(n_T_427[1879]), .A3(n_T_427[1771]), .A4(
        n2866), .Y(n2761) );
  AOI22X1_LVT U4613 ( .A1(n3828), .A2(n_T_427[1832]), .A3(n_T_427[1707]), .A4(
        n3825), .Y(n2762) );
  AND4X1_LVT U4614 ( .A1(n2766), .A2(n2767), .A3(n2768), .A4(n2769), .Y(n6047)
         );
  AOI22X1_LVT U4615 ( .A1(n3801), .A2(n_T_427[1872]), .A3(n3884), .A4(
        n_T_427[1910]), .Y(n2767) );
  AOI22X1_LVT U4616 ( .A1(n3826), .A2(n_T_427[1692]), .A3(n_T_427[1564]), .A4(
        n3890), .Y(n2768) );
  AOI22X1_LVT U4617 ( .A1(n3889), .A2(n_T_427[1628]), .A3(n_T_427[1500]), .A4(
        n3922), .Y(n2769) );
  AND4X1_LVT U4618 ( .A1(n2770), .A2(n2771), .A3(n2772), .A4(n2773), .Y(n6011)
         );
  AOI22X1_LVT U4619 ( .A1(n6764), .A2(n_T_427[1870]), .A3(n_T_427[1754]), .A4(
        n2867), .Y(n2770) );
  AOI22X1_LVT U4620 ( .A1(n3830), .A2(n_T_427[1816]), .A3(n_T_427[1690]), .A4(
        n3826), .Y(n2771) );
  AOI22X1_LVT U4621 ( .A1(n3892), .A2(n_T_427[1562]), .A3(n_T_427[1626]), .A4(
        n3886), .Y(n2772) );
  AND4X1_LVT U4622 ( .A1(n2774), .A2(n2775), .A3(n2776), .A4(n2777), .Y(n5897)
         );
  AOI22X1_LVT U4623 ( .A1(n3798), .A2(n_T_427[1749]), .A3(n_T_427[1811]), .A4(
        n2765), .Y(n2774) );
  AOI22X1_LVT U4624 ( .A1(n3827), .A2(n_T_427[1685]), .A3(n_T_427[1557]), .A4(
        n3890), .Y(n2776) );
  AOI22X1_LVT U4625 ( .A1(n3889), .A2(n_T_427[1621]), .A3(n_T_427[1493]), .A4(
        n3922), .Y(n2777) );
  AND4X1_LVT U4626 ( .A1(n2778), .A2(n2779), .A3(n2780), .A4(n2781), .Y(n6435)
         );
  AOI22X1_LVT U4627 ( .A1(n3802), .A2(n_T_427[1880]), .A3(n_T_427[1773]), .A4(
        n2867), .Y(n2778) );
  AOI22X1_LVT U4628 ( .A1(n3828), .A2(n_T_427[1834]), .A3(n_T_427[1709]), .A4(
        n3825), .Y(n2779) );
  AND4X1_LVT U4629 ( .A1(n2782), .A2(n2783), .A3(n2784), .A4(n2785), .Y(n5552)
         );
  AOI22X1_LVT U4630 ( .A1(n6764), .A2(n_T_427[1851]), .A3(n_T_427[1732]), .A4(
        n2866), .Y(n2782) );
  AOI22X1_LVT U4631 ( .A1(n3828), .A2(n_T_427[1795]), .A3(n_T_427[1668]), .A4(
        n3826), .Y(n2783) );
  AOI22X1_LVT U4632 ( .A1(n3892), .A2(n_T_427[1540]), .A3(n_T_427[1604]), .A4(
        n3885), .Y(n2784) );
  AND4X1_LVT U4633 ( .A1(n2786), .A2(n2787), .A3(n2788), .A4(n2789), .Y(n5501)
         );
  AOI22X1_LVT U4634 ( .A1(n3802), .A2(n_T_427[1848]), .A3(n_T_427[1729]), .A4(
        n2867), .Y(n2786) );
  AOI22X1_LVT U4635 ( .A1(n3829), .A2(n_T_427[1792]), .A3(n_T_427[1665]), .A4(
        n3826), .Y(n2787) );
  AND4X1_LVT U4636 ( .A1(n2791), .A2(n2792), .A3(n2793), .A4(n2794), .Y(n5670)
         );
  AOI22X1_LVT U4637 ( .A1(n3801), .A2(n_T_427[1856]), .A3(n_T_427[1737]), .A4(
        n2868), .Y(n2791) );
  AOI22X1_LVT U4638 ( .A1(n3830), .A2(n_T_427[1800]), .A3(n_T_427[1673]), .A4(
        n3826), .Y(n2792) );
  AOI22X1_LVT U4639 ( .A1(n3891), .A2(n_T_427[1545]), .A3(n_T_427[1609]), .A4(
        n3885), .Y(n2793) );
  AND4X1_LVT U4640 ( .A1(n2795), .A2(n2796), .A3(n2797), .A4(n2798), .Y(n5622)
         );
  AOI22X1_LVT U4641 ( .A1(n3802), .A2(n_T_427[1854]), .A3(n_T_427[1735]), .A4(
        n2867), .Y(n2795) );
  AOI22X1_LVT U4642 ( .A1(n2765), .A2(n_T_427[1798]), .A3(n_T_427[1671]), .A4(
        n3826), .Y(n2796) );
  AOI22X1_LVT U4643 ( .A1(n3891), .A2(n_T_427[1543]), .A3(n_T_427[1607]), .A4(
        n3885), .Y(n2797) );
  AOI22X1_LVT U4644 ( .A1(n3923), .A2(n_T_427[1479]), .A3(n_T_427[1351]), .A4(
        n3917), .Y(n2798) );
  AND4X1_LVT U4645 ( .A1(n2799), .A2(n2800), .A3(n2801), .A4(n2802), .Y(n5857)
         );
  AOI22X1_LVT U4646 ( .A1(n3802), .A2(n_T_427[1865]), .A3(n_T_427[1747]), .A4(
        n2866), .Y(n2799) );
  AOI22X1_LVT U4647 ( .A1(n3892), .A2(n_T_427[1555]), .A3(n_T_427[1619]), .A4(
        n3886), .Y(n2801) );
  AND4X1_LVT U4648 ( .A1(n2803), .A2(n2804), .A3(n2805), .A4(n2806), .Y(n5701)
         );
  AOI22X1_LVT U4649 ( .A1(n3801), .A2(n_T_427[1858]), .A3(n_T_427[1739]), .A4(
        n2868), .Y(n2803) );
  AOI22X1_LVT U4650 ( .A1(n3828), .A2(n_T_427[1802]), .A3(n_T_427[1675]), .A4(
        n3826), .Y(n2804) );
  AOI22X1_LVT U4651 ( .A1(n3891), .A2(n_T_427[1547]), .A3(n_T_427[1611]), .A4(
        n3885), .Y(n2805) );
  AOI22X1_LVT U4652 ( .A1(n3923), .A2(n_T_427[1483]), .A3(n_T_427[1355]), .A4(
        n3917), .Y(n2806) );
  AND4X1_LVT U4653 ( .A1(n2807), .A2(n2808), .A3(n2809), .A4(n2810), .Y(n5578)
         );
  AOI22X1_LVT U4654 ( .A1(n3802), .A2(n_T_427[1852]), .A3(n_T_427[1733]), .A4(
        n2868), .Y(n2807) );
  AOI22X1_LVT U4655 ( .A1(n3829), .A2(n_T_427[1796]), .A3(n_T_427[1669]), .A4(
        n3826), .Y(n2808) );
  AOI22X1_LVT U4656 ( .A1(n3891), .A2(n_T_427[1541]), .A3(n_T_427[1605]), .A4(
        n3885), .Y(n2809) );
  AOI22X1_LVT U4657 ( .A1(n3923), .A2(n_T_427[1477]), .A3(n_T_427[1349]), .A4(
        n3917), .Y(n2810) );
  AND4X1_LVT U4658 ( .A1(n2811), .A2(n2812), .A3(n2813), .A4(n2814), .Y(n5646)
         );
  AOI22X1_LVT U4659 ( .A1(n3801), .A2(n_T_427[1855]), .A3(n_T_427[1736]), .A4(
        n2866), .Y(n2811) );
  AOI22X1_LVT U4660 ( .A1(n3830), .A2(n_T_427[1799]), .A3(n_T_427[1672]), .A4(
        n3826), .Y(n2812) );
  AOI22X1_LVT U4661 ( .A1(n3891), .A2(n_T_427[1544]), .A3(n_T_427[1608]), .A4(
        n3885), .Y(n2813) );
  AND4X1_LVT U4662 ( .A1(n2815), .A2(n2816), .A3(n2817), .A4(n2818), .Y(n5820)
         );
  AOI22X1_LVT U4663 ( .A1(n6764), .A2(n_T_427[1863]), .A3(n_T_427[1745]), .A4(
        n2867), .Y(n2815) );
  AOI22X1_LVT U4664 ( .A1(n3830), .A2(n_T_427[1807]), .A3(n_T_427[1681]), .A4(
        n3825), .Y(n2816) );
  AOI22X1_LVT U4665 ( .A1(n3892), .A2(n_T_427[1553]), .A3(n_T_427[1617]), .A4(
        n3886), .Y(n2817) );
  AOI22X1_LVT U4666 ( .A1(n2028), .A2(n_T_427[1860]), .A3(n_T_427[1741]), .A4(
        n3798), .Y(n2819) );
  AND4X1_LVT U4667 ( .A1(n2820), .A2(n2821), .A3(n2822), .A4(n2823), .Y(n6786)
         );
  AOI22X1_LVT U4668 ( .A1(n6764), .A2(n_T_427[1881]), .A3(n_T_427[1787]), .A4(
        n3798), .Y(n2820) );
  NBUFFX2_LVT U4669 ( .A(n6887), .Y(n2824) );
  NBUFFX2_LVT U4670 ( .A(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(n2825) );
  NBUFFX2_LVT U4671 ( .A(n6888), .Y(n2826) );
  NBUFFX2_LVT U4672 ( .A(n6884), .Y(n2827) );
  NBUFFX2_LVT U4673 ( .A(n6774), .Y(n2828) );
  NBUFFX2_LVT U4674 ( .A(n6812), .Y(n2829) );
  NBUFFX2_LVT U4675 ( .A(n6773), .Y(n2830) );
  IBUFFX2_LVT U4676 ( .A(n3781), .Y(n5436) );
  INVX1_LVT U4677 ( .A(n5906), .Y(n6796) );
  NBUFFX2_LVT U4678 ( .A(n6882), .Y(n2831) );
  NBUFFX2_LVT U4679 ( .A(n6882), .Y(n2832) );
  AOI22X1_LVT U4680 ( .A1(n3895), .A2(n_T_427[926]), .A3(n_T_427[735]), .A4(
        n3904), .Y(n2846) );
  AOI22X1_LVT U4681 ( .A1(n3834), .A2(n_T_427[385]), .A3(n_T_427[65]), .A4(
        n3832), .Y(n2852) );
  NBUFFX2_LVT U4682 ( .A(n6813), .Y(n2833) );
  NAND2X0_LVT U4683 ( .A1(n2834), .A2(n2835), .Y(n5060) );
  AND3X1_LVT U4684 ( .A1(n5008), .A2(n5007), .A3(n5006), .Y(n2835) );
  NBUFFX2_LVT U4685 ( .A(n9041), .Y(n2836) );
  NBUFFX2_LVT U4686 ( .A(n9041), .Y(n2837) );
  XOR2X1_LVT U4687 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n3202), .Y(
        n4846) );
  AOI22X1_LVT U4688 ( .A1(n3835), .A2(n_T_427[403]), .A3(n_T_427[83]), .A4(
        n2871), .Y(n2838) );
  AOI22X1_LVT U4689 ( .A1(n3817), .A2(n_T_427[339]), .A3(n6774), .A4(
        n_T_427[275]), .Y(n2840) );
  AND2X1_LVT U4690 ( .A1(n5833), .A2(n5832), .Y(n2841) );
  AND4X1_LVT U4691 ( .A1(n2842), .A2(n2843), .A3(n2844), .A4(n2845), .Y(n5877)
         );
  AND2X1_LVT U4692 ( .A1(n5870), .A2(n5869), .Y(n2842) );
  AND4X1_LVT U4693 ( .A1(n2846), .A2(n2847), .A3(n2848), .A4(n2849), .Y(n6097)
         );
  AOI22X1_LVT U4694 ( .A1(n3823), .A2(n_T_427[862]), .A3(n_T_427[159]), .A4(
        n2863), .Y(n2848) );
  AND2X1_LVT U4695 ( .A1(n6089), .A2(n6090), .Y(n2849) );
  NBUFFX2_LVT U4696 ( .A(n6811), .Y(n2850) );
  NBUFFX2_LVT U4697 ( .A(n6811), .Y(n2851) );
  INVX1_LVT U4698 ( .A(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(n4816) );
  AOI22X1_LVT U4699 ( .A1(n3943), .A2(n_T_427[1152]), .A3(n_T_427[1024]), .A4(
        n3898), .Y(n2853) );
  AOI22X1_LVT U4700 ( .A1(n3953), .A2(n_T_427[1088]), .A3(n_T_427[960]), .A4(
        n3947), .Y(n2854) );
  IBUFFX2_LVT U4701 ( .A(n6423), .Y(n6865) );
  NBUFFX2_LVT U4702 ( .A(n6810), .Y(n2856) );
  NBUFFX2_LVT U4703 ( .A(n6810), .Y(n2857) );
  NBUFFX2_LVT U4704 ( .A(n8932), .Y(n2858) );
  NBUFFX2_LVT U4705 ( .A(n6885), .Y(n2860) );
  NBUFFX2_LVT U4706 ( .A(n6885), .Y(n2861) );
  NBUFFX2_LVT U4707 ( .A(n6886), .Y(n2862) );
  NBUFFX2_LVT U4708 ( .A(n6886), .Y(n2863) );
  NBUFFX2_LVT U4709 ( .A(n6830), .Y(n2864) );
  NBUFFX2_LVT U4710 ( .A(n6830), .Y(n2865) );
  NBUFFX2_LVT U4711 ( .A(n6763), .Y(n2866) );
  IBUFFX2_LVT U4712 ( .A(n3799), .Y(n2867) );
  IBUFFX2_LVT U4713 ( .A(n3799), .Y(n2868) );
  AND2X1_LVT U4714 ( .A1(n5446), .A2(n2034), .Y(n6763) );
  IBUFFX2_LVT U4715 ( .A(n6763), .Y(n3800) );
  NBUFFX2_LVT U4716 ( .A(n6889), .Y(n2869) );
  NBUFFX2_LVT U4717 ( .A(n6889), .Y(n2870) );
  NBUFFX2_LVT U4718 ( .A(n6829), .Y(n2871) );
  NBUFFX2_LVT U4719 ( .A(n6829), .Y(n2872) );
  AND2X1_LVT U4720 ( .A1(n9417), .A2(n5062), .Y(n2873) );
  AND3X1_LVT U4721 ( .A1(n5395), .A2(n5396), .A3(n406), .Y(n5401) );
  NAND2X0_LVT U4722 ( .A1(n9417), .A2(n5062), .Y(n2874) );
  AND2X1_LVT U4723 ( .A1(n406), .A2(n9383), .Y(N744) );
  AND2X1_LVT U4724 ( .A1(n2873), .A2(n9382), .Y(N745) );
  AND2X1_LVT U4725 ( .A1(n9286), .A2(n2873), .Y(io_fpu_valid) );
  AND2X1_LVT U4726 ( .A1(n9417), .A2(n5062), .Y(n406) );
  NBUFFX2_LVT U4727 ( .A(ibuf_io_inst_0_bits_inst_rs1[1]), .Y(n2876) );
  NBUFFX2_LVT U4728 ( .A(ibuf_io_inst_0_bits_inst_rs1[1]), .Y(n2877) );
  NBUFFX2_LVT U4729 ( .A(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(n2878) );
  NBUFFX2_LVT U4730 ( .A(n6888), .Y(n2879) );
  AND2X1_LVT U4731 ( .A1(n5444), .A2(n5445), .Y(n2881) );
  IBUFFX2_LVT U4732 ( .A(n3012), .Y(n2882) );
  AND3X1_LVT U4733 ( .A1(n6986), .A2(n6985), .A3(n6984), .Y(n2883) );
  AND3X1_LVT U4734 ( .A1(n6982), .A2(n6981), .A3(n6980), .Y(n2884) );
  INVX1_LVT U4735 ( .A(n6766), .Y(n6868) );
  AND3X1_LVT U4736 ( .A1(n7118), .A2(n7117), .A3(n7116), .Y(n2885) );
  AND3X1_LVT U4737 ( .A1(n7114), .A2(n7113), .A3(n7112), .Y(n2886) );
  AND3X1_LVT U4738 ( .A1(n7397), .A2(n7396), .A3(n7395), .Y(n2887) );
  AND3X1_LVT U4739 ( .A1(n7393), .A2(n7392), .A3(n7391), .Y(n2888) );
  AND3X1_LVT U4740 ( .A1(n7312), .A2(n7311), .A3(n7310), .Y(n2889) );
  AND3X1_LVT U4741 ( .A1(n7308), .A2(n7307), .A3(n7306), .Y(n2890) );
  AND3X1_LVT U4742 ( .A1(n7256), .A2(n7255), .A3(n7254), .Y(n2891) );
  AND3X1_LVT U4743 ( .A1(n7252), .A2(n7251), .A3(n7250), .Y(n2892) );
  AND3X1_LVT U4744 ( .A1(n7230), .A2(n7229), .A3(n7228), .Y(n2893) );
  AND3X1_LVT U4745 ( .A1(n7226), .A2(n7225), .A3(n7224), .Y(n2894) );
  AND3X1_LVT U4746 ( .A1(n7058), .A2(n7057), .A3(n7056), .Y(n2895) );
  AND3X1_LVT U4747 ( .A1(n7054), .A2(n7053), .A3(n7052), .Y(n2896) );
  AND3X1_LVT U4748 ( .A1(n6988), .A2(n6989), .A3(n6990), .Y(n2898) );
  AND3X1_LVT U4749 ( .A1(n7014), .A2(n7013), .A3(n7012), .Y(n2899) );
  AND3X1_LVT U4750 ( .A1(n6998), .A2(n6997), .A3(n6996), .Y(n2900) );
  NAND3X0_LVT U4751 ( .A1(n2901), .A2(n2902), .A3(n2903), .Y(N673) );
  AND3X1_LVT U4752 ( .A1(n2953), .A2(n2954), .A3(n2955), .Y(n2901) );
  AND3X1_LVT U4753 ( .A1(n6929), .A2(n6928), .A3(n6927), .Y(n2902) );
  AND3X1_LVT U4754 ( .A1(n6921), .A2(n6920), .A3(n6919), .Y(n2903) );
  AND3X1_LVT U4755 ( .A1(n7368), .A2(n7367), .A3(n7366), .Y(n2904) );
  AND3X1_LVT U4756 ( .A1(n7364), .A2(n7363), .A3(n7362), .Y(n2905) );
  AND3X1_LVT U4757 ( .A1(n7146), .A2(n7145), .A3(n7144), .Y(n2906) );
  AND3X1_LVT U4758 ( .A1(n7142), .A2(n7141), .A3(n7140), .Y(n2907) );
  AND3X1_LVT U4759 ( .A1(n7030), .A2(n7029), .A3(n7028), .Y(n2908) );
  AND3X1_LVT U4760 ( .A1(n7026), .A2(n7025), .A3(n7024), .Y(n2909) );
  AND3X1_LVT U4761 ( .A1(n8733), .A2(n8732), .A3(n8731), .Y(n2911) );
  AND4X1_LVT U4762 ( .A1(n2912), .A2(n2913), .A3(n2914), .A4(n2915), .Y(n5463)
         );
  OA22X1_LVT U4763 ( .A1(n1994), .A2(n3633), .A3(n3256), .A4(n3799), .Y(n2912)
         );
  AOI22X1_LVT U4764 ( .A1(n3828), .A2(n_T_427[1791]), .A3(n_T_427[1663]), .A4(
        n3824), .Y(n2913) );
  AOI22X1_LVT U4765 ( .A1(n3892), .A2(n_T_427[1535]), .A3(n_T_427[1599]), .A4(
        n3886), .Y(n2914) );
  AOI22X1_LVT U4766 ( .A1(n3924), .A2(n_T_427[1471]), .A3(n_T_427[1343]), .A4(
        n3919), .Y(n2915) );
  AND3X1_LVT U4767 ( .A1(n7341), .A2(n7340), .A3(n7339), .Y(n2916) );
  AND3X1_LVT U4768 ( .A1(n7337), .A2(n7336), .A3(n7335), .Y(n2917) );
  AND3X1_LVT U4769 ( .A1(n7932), .A2(n7931), .A3(n7930), .Y(n2918) );
  AND3X1_LVT U4770 ( .A1(n7928), .A2(n7927), .A3(n7926), .Y(n2919) );
  AND2X1_LVT U4771 ( .A1(n2920), .A2(n2921), .Y(n3741) );
  AND3X1_LVT U4772 ( .A1(n8441), .A2(n8440), .A3(n8439), .Y(n2920) );
  AND3X1_LVT U4773 ( .A1(n8445), .A2(n8444), .A3(n8443), .Y(n2921) );
  NBUFFX2_LVT U4774 ( .A(n9012), .Y(n2922) );
  AND3X1_LVT U4775 ( .A1(n7997), .A2(n7996), .A3(n7995), .Y(n2923) );
  AND3X1_LVT U4776 ( .A1(n8001), .A2(n8000), .A3(n7999), .Y(n2924) );
  AND2X1_LVT U4777 ( .A1(n3623), .A2(n3622), .Y(n2925) );
  AND3X1_LVT U4778 ( .A1(n8030), .A2(n8029), .A3(n8028), .Y(n2926) );
  AND3X1_LVT U4779 ( .A1(n8034), .A2(n8033), .A3(n8032), .Y(n2927) );
  OA22X1_LVT U4780 ( .A1(n2875), .A2(n3654), .A3(n3257), .A4(n3799), .Y(n2928)
         );
  AOI22X1_LVT U4781 ( .A1(n3827), .A2(n_T_427[1664]), .A3(n_T_427[1600]), .A4(
        n3885), .Y(n2929) );
  AOI22X1_LVT U4782 ( .A1(n3891), .A2(n_T_427[1536]), .A3(n_T_427[1408]), .A4(
        n3932), .Y(n2930) );
  AOI22X1_LVT U4783 ( .A1(n3923), .A2(n_T_427[1472]), .A3(n_T_427[1344]), .A4(
        n3917), .Y(n2931) );
  AND3X1_LVT U4784 ( .A1(n8293), .A2(n8292), .A3(n8291), .Y(n2932) );
  AND3X1_LVT U4785 ( .A1(n8289), .A2(n8288), .A3(n8287), .Y(n2933) );
  AND2X1_LVT U4786 ( .A1(n8278), .A2(n8277), .Y(n2934) );
  AND3X1_LVT U4787 ( .A1(n7277), .A2(n7276), .A3(n7275), .Y(n2935) );
  AND3X1_LVT U4788 ( .A1(n7269), .A2(n7268), .A3(n7267), .Y(n2936) );
  AND3X1_LVT U4789 ( .A1(n7243), .A2(n7242), .A3(n7241), .Y(n2937) );
  AND3X1_LVT U4790 ( .A1(n7410), .A2(n7409), .A3(n7408), .Y(n2938) );
  AND3X1_LVT U4791 ( .A1(n7329), .A2(n7328), .A3(n7327), .Y(n2939) );
  AND3X1_LVT U4792 ( .A1(n7333), .A2(n7332), .A3(n7331), .Y(n2940) );
  AND3X1_LVT U4793 ( .A1(n7325), .A2(n7324), .A3(n7323), .Y(n2941) );
  AND3X1_LVT U4794 ( .A1(n7075), .A2(n7074), .A3(n7073), .Y(n2942) );
  AND3X1_LVT U4795 ( .A1(n7079), .A2(n7078), .A3(n7077), .Y(n2943) );
  AND3X1_LVT U4796 ( .A1(n7071), .A2(n7070), .A3(n7069), .Y(n2944) );
  NAND3X0_LVT U4797 ( .A1(n2945), .A2(n2946), .A3(n2947), .Y(N728) );
  AND3X1_LVT U4798 ( .A1(n8487), .A2(n8486), .A3(n8485), .Y(n2946) );
  NOR2X0_LVT U4799 ( .A1(n8497), .A2(n8496), .Y(n2947) );
  AND3X1_LVT U4800 ( .A1(n8249), .A2(n8248), .A3(n8247), .Y(n2948) );
  AND3X1_LVT U4801 ( .A1(n8245), .A2(n8244), .A3(n8243), .Y(n2949) );
  AND2X1_LVT U4802 ( .A1(n8096), .A2(n8095), .Y(n2951) );
  AND3X1_LVT U4803 ( .A1(n8094), .A2(n8092), .A3(n8093), .Y(n2952) );
  AND3X1_LVT U4804 ( .A1(n6944), .A2(n6943), .A3(n6942), .Y(n2953) );
  AND3X1_LVT U4805 ( .A1(n6934), .A2(n6933), .A3(n6932), .Y(n2954) );
  AND3X1_LVT U4806 ( .A1(n6978), .A2(n6977), .A3(n6976), .Y(n2955) );
  AND2X1_LVT U4807 ( .A1(n8345), .A2(n8344), .Y(n2956) );
  AND3X1_LVT U4808 ( .A1(n8343), .A2(n8341), .A3(n8342), .Y(n2957) );
  AND3X1_LVT U4809 ( .A1(n7358), .A2(n7359), .A3(n7360), .Y(n2959) );
  AND3X1_LVT U4810 ( .A1(n7354), .A2(n7353), .A3(n7352), .Y(n2960) );
  AND2X1_LVT U4811 ( .A1(n8478), .A2(n8477), .Y(n2961) );
  AND3X1_LVT U4812 ( .A1(n8476), .A2(n8474), .A3(n8475), .Y(n2962) );
  AND2X1_LVT U4813 ( .A1(n7954), .A2(n7953), .Y(n2964) );
  AND3X1_LVT U4814 ( .A1(n7952), .A2(n7951), .A3(n7950), .Y(n2965) );
  AND3X2_LVT U4815 ( .A1(n3773), .A2(n6946), .A3(n6973), .Y(n2966) );
  NBUFFX2_LVT U4816 ( .A(n9007), .Y(n2967) );
  AND2X1_LVT U4817 ( .A1(n4027), .A2(n8105), .Y(n8991) );
  AND2X1_LVT U4818 ( .A1(n4051), .A2(n8105), .Y(n8944) );
  AND2X1_LVT U4819 ( .A1(n4041), .A2(n8105), .Y(n8994) );
  AND2X1_LVT U4820 ( .A1(n3973), .A2(n8105), .Y(n9059) );
  AND2X4_LVT U4821 ( .A1(n8105), .A2(n3979), .Y(n9056) );
  AND2X1_LVT U4822 ( .A1(n4845), .A2(n4844), .Y(n2968) );
  AND2X1_LVT U4823 ( .A1(n5067), .A2(io_fpu_inst[4]), .Y(n5106) );
  AND3X2_LVT U4824 ( .A1(n6973), .A2(n6926), .A3(n2983), .Y(n9029) );
  NAND2X0_LVT U4825 ( .A1(n7910), .A2(n7911), .Y(n9047) );
  AND3X1_LVT U4826 ( .A1(n7389), .A2(n7388), .A3(n7387), .Y(n2970) );
  AND3X1_LVT U4827 ( .A1(n7383), .A2(n7384), .A3(n7385), .Y(n2971) );
  AND3X1_LVT U4828 ( .A1(n7381), .A2(n7380), .A3(n7379), .Y(n2972) );
  AND3X1_LVT U4829 ( .A1(n7222), .A2(n7221), .A3(n7220), .Y(n2973) );
  AND3X1_LVT U4830 ( .A1(n7214), .A2(n7213), .A3(n7212), .Y(n2974) );
  AND3X1_LVT U4831 ( .A1(n7167), .A2(n7166), .A3(n7165), .Y(n2975) );
  AND3X1_LVT U4832 ( .A1(n7161), .A2(n7162), .A3(n7163), .Y(n2976) );
  AND3X1_LVT U4833 ( .A1(n7159), .A2(n7158), .A3(n7157), .Y(n2977) );
  AND3X1_LVT U4834 ( .A1(n7050), .A2(n7049), .A3(n7048), .Y(n2978) );
  AND3X1_LVT U4835 ( .A1(n7043), .A2(n7042), .A3(n7041), .Y(n2979) );
  OR2X1_LVT U4836 ( .A1(n2069), .A2(n2980), .Y(n8246) );
  AND3X1_LVT U4837 ( .A1(n6964), .A2(n6963), .A3(n2627), .Y(n7910) );
  IBUFFX2_LVT U4838 ( .A(n3012), .Y(n2985) );
  IBUFFX2_LVT U4839 ( .A(n3012), .Y(n2986) );
  AND3X1_LVT U4840 ( .A1(n8954), .A2(n8953), .A3(n8952), .Y(n2988) );
  AND3X1_LVT U4841 ( .A1(n8950), .A2(n8949), .A3(n8948), .Y(n2989) );
  AND2X1_LVT U4842 ( .A1(n2990), .A2(n2991), .Y(n3738) );
  AND3X1_LVT U4843 ( .A1(n8509), .A2(n8508), .A3(n8507), .Y(n2990) );
  AND3X1_LVT U4844 ( .A1(n8505), .A2(n8504), .A3(n8503), .Y(n2991) );
  AND2X1_LVT U4845 ( .A1(n2992), .A2(n2993), .Y(n3034) );
  AND3X1_LVT U4846 ( .A1(n8303), .A2(n8304), .A3(n8305), .Y(n2992) );
  AND3X1_LVT U4847 ( .A1(n8301), .A2(n8300), .A3(n8299), .Y(n2993) );
  AND2X1_LVT U4848 ( .A1(n2994), .A2(n2995), .Y(n3731) );
  AND3X1_LVT U4849 ( .A1(n8827), .A2(n8826), .A3(n8825), .Y(n2994) );
  AND3X1_LVT U4850 ( .A1(n8823), .A2(n8822), .A3(n8821), .Y(n2995) );
  AND2X1_LVT U4851 ( .A1(n2996), .A2(n2997), .Y(n3735) );
  AND3X1_LVT U4852 ( .A1(n8612), .A2(n8611), .A3(n8610), .Y(n2996) );
  AND3X1_LVT U4853 ( .A1(n8608), .A2(n8607), .A3(n8606), .Y(n2997) );
  NBUFFX2_LVT U4854 ( .A(n9008), .Y(n2998) );
  NAND3X0_LVT U4855 ( .A1(n3001), .A2(n3000), .A3(n2999), .Y(N699) );
  AND3X1_LVT U4856 ( .A1(n3680), .A2(n3681), .A3(n3682), .Y(n2999) );
  AND3X1_LVT U4857 ( .A1(n7511), .A2(n7510), .A3(n7509), .Y(n3000) );
  AND3X1_LVT U4858 ( .A1(n7507), .A2(n7506), .A3(n7505), .Y(n3001) );
  NAND3X0_LVT U4859 ( .A1(n3002), .A2(n3003), .A3(n3004), .Y(N709) );
  AND3X1_LVT U4860 ( .A1(n3057), .A2(n3058), .A3(n3059), .Y(n3002) );
  AND3X1_LVT U4861 ( .A1(n7827), .A2(n7826), .A3(n7825), .Y(n3003) );
  AND3X1_LVT U4862 ( .A1(n7823), .A2(n7822), .A3(n7821), .Y(n3004) );
  AND3X1_LVT U4863 ( .A1(n7856), .A2(n7855), .A3(n7854), .Y(n3005) );
  AND3X1_LVT U4864 ( .A1(n7852), .A2(n7851), .A3(n7850), .Y(n3006) );
  AND3X1_LVT U4865 ( .A1(n7478), .A2(n7477), .A3(n7476), .Y(n3007) );
  AND3X1_LVT U4866 ( .A1(n7474), .A2(n7473), .A3(n7472), .Y(n3008) );
  NAND3X0_LVT U4867 ( .A1(n3011), .A2(n3010), .A3(n3009), .Y(N703) );
  AND3X1_LVT U4868 ( .A1(n3066), .A2(n3067), .A3(n3068), .Y(n3009) );
  AND3X1_LVT U4869 ( .A1(n7634), .A2(n7633), .A3(n7632), .Y(n3010) );
  AND3X1_LVT U4870 ( .A1(n7630), .A2(n7629), .A3(n7628), .Y(n3011) );
  OA22X1_LVT U4871 ( .A1(n3993), .A2(n3524), .A3(n3178), .A4(n3988), .Y(n3568)
         );
  AND3X1_LVT U4872 ( .A1(n7697), .A2(n7696), .A3(n7695), .Y(n3013) );
  AND3X1_LVT U4873 ( .A1(n7693), .A2(n7692), .A3(n7691), .Y(n3014) );
  AND3X1_LVT U4874 ( .A1(n7730), .A2(n7729), .A3(n7728), .Y(n3015) );
  AND3X1_LVT U4875 ( .A1(n7726), .A2(n7725), .A3(n7724), .Y(n3016) );
  NAND3X0_LVT U4876 ( .A1(n3017), .A2(n3018), .A3(n3019), .Y(N700) );
  AND3X1_LVT U4877 ( .A1(n7540), .A2(n7539), .A3(n7538), .Y(n3018) );
  AND3X1_LVT U4878 ( .A1(n7536), .A2(n7535), .A3(n7534), .Y(n3019) );
  AND3X1_LVT U4879 ( .A1(n7450), .A2(n7449), .A3(n7448), .Y(n3020) );
  AND3X1_LVT U4880 ( .A1(n7446), .A2(n7445), .A3(n7444), .Y(n3021) );
  AND3X1_LVT U4881 ( .A1(n7571), .A2(n7570), .A3(n7569), .Y(n3022) );
  AND3X1_LVT U4882 ( .A1(n7567), .A2(n7566), .A3(n7565), .Y(n3023) );
  AND2X1_LVT U4883 ( .A1(n3024), .A2(n3025), .Y(n3728) );
  AND3X1_LVT U4884 ( .A1(n8859), .A2(n8858), .A3(n8857), .Y(n3024) );
  AND3X1_LVT U4885 ( .A1(n8861), .A2(n8862), .A3(n8863), .Y(n3025) );
  AND2X1_LVT U4886 ( .A1(n3026), .A2(n3027), .Y(n3748) );
  AND3X1_LVT U4887 ( .A1(n9011), .A2(n9010), .A3(n9009), .Y(n3026) );
  AND3X1_LVT U4888 ( .A1(n9017), .A2(n9018), .A3(n9019), .Y(n3027) );
  NAND3X0_LVT U4889 ( .A1(n3028), .A2(n3029), .A3(n3030), .Y(N702) );
  AND3X1_LVT U4890 ( .A1(n7603), .A2(n7602), .A3(n7601), .Y(n3029) );
  AND3X1_LVT U4891 ( .A1(n7599), .A2(n7598), .A3(n7597), .Y(n3030) );
  NAND2X0_LVT U4892 ( .A1(n9231), .A2(n3031), .Y(n3574) );
  AND2X1_LVT U4893 ( .A1(n3575), .A2(csr_io_status_isa[12]), .Y(n3031) );
  NAND2X0_LVT U4894 ( .A1(n3032), .A2(n3033), .Y(n8774) );
  AND3X1_LVT U4895 ( .A1(n8768), .A2(n8769), .A3(n8767), .Y(n3032) );
  AND3X1_LVT U4896 ( .A1(n8773), .A2(n8772), .A3(n8771), .Y(n3033) );
  NAND3X0_LVT U4897 ( .A1(n3034), .A2(n3036), .A3(n3035), .Y(N723) );
  NOR3X0_LVT U4898 ( .A1(n8329), .A2(n8328), .A3(n8327), .Y(n3036) );
  NAND2X0_LVT U4899 ( .A1(n3037), .A2(n3038), .Y(n8923) );
  AND3X1_LVT U4900 ( .A1(n8918), .A2(n8917), .A3(n8916), .Y(n3037) );
  AND3X1_LVT U4901 ( .A1(n8922), .A2(n8921), .A3(n8920), .Y(n3038) );
  IBUFFX2_LVT U4902 ( .A(n6877), .Y(n3879) );
  IBUFFX2_LVT U4903 ( .A(n3082), .Y(n3826) );
  IBUFFX2_LVT U4904 ( .A(n3082), .Y(n3825) );
  MUX21X1_LVT U4905 ( .A1(n3041), .A2(n5306), .S0(n9381), .Y(n3040) );
  IBUFFX2_LVT U4906 ( .A(n9529), .Y(n3044) );
  AND2X1_LVT U4907 ( .A1(n3044), .A2(n5074), .Y(n9076) );
  NAND3X0_LVT U4908 ( .A1(n4843), .A2(n3044), .A3(n4842), .Y(n4845) );
  NAND3X0_LVT U4909 ( .A1(n9091), .A2(n1867), .A3(n9090), .Y(n9092) );
  IBUFFX2_LVT U4910 ( .A(n5075), .Y(n9075) );
  OR3X1_LVT U4911 ( .A1(reset), .A2(n3046), .A3(n9380), .Y(N746) );
  INVX1_LVT U4912 ( .A(n5905), .Y(n6838) );
  XOR2X1_LVT U4913 ( .A1(n2037), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5425) );
  NAND3X0_LVT U4914 ( .A1(n9439), .A2(n2553), .A3(n5097), .Y(n5098) );
  AND3X2_LVT U4915 ( .A1(n6973), .A2(n6931), .A3(n3709), .Y(n9004) );
  AND3X2_LVT U4916 ( .A1(n6973), .A2(n6931), .A3(n3709), .Y(n3613) );
  XOR2X1_LVT U4917 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n2574), .Y(
        n5431) );
  MUX21X1_LVT U4918 ( .A1(n3199), .A2(n5426), .S0(n9381), .Y(n9403) );
  MUX21X1_LVT U4919 ( .A1(n3198), .A2(n5428), .S0(n9381), .Y(n9398) );
  AND2X1_LVT U4920 ( .A1(n4971), .A2(n4752), .Y(n6972) );
  INVX1_LVT U4921 ( .A(ibuf_io_inst_0_bits_inst_rs1[2]), .Y(n4752) );
  IBUFFX2_LVT U4922 ( .A(n9522), .Y(n9440) );
  IBUFFX2_LVT U4923 ( .A(n5099), .Y(n5138) );
  AND3X1_LVT U4924 ( .A1(n8958), .A2(n8957), .A3(n8956), .Y(n3050) );
  NOR2X4_LVT U4925 ( .A1(n2552), .A2(n9528), .Y(n9107) );
  AOI22X1_LVT U4926 ( .A1(n2570), .A2(io_fpu_inst[13]), .A3(io_fpu_inst[5]), 
        .A4(n9107), .Y(n4844) );
  IBUFFX2_LVT U4927 ( .A(n9526), .Y(n9105) );
  IBUFFX2_LVT U4928 ( .A(n9107), .Y(n9096) );
  AO22X1_LVT U4929 ( .A1(n5173), .A2(n5174), .A3(n9107), .A4(n9097), .Y(
        id_ctrl_wfd) );
  AND3X1_LVT U4930 ( .A1(n7802), .A2(n7801), .A3(n7800), .Y(n3051) );
  AND3X1_LVT U4931 ( .A1(n7815), .A2(n7813), .A3(n7814), .Y(n3052) );
  AND3X1_LVT U4932 ( .A1(n7798), .A2(n7797), .A3(n7796), .Y(n3053) );
  AND3X1_LVT U4933 ( .A1(n7890), .A2(n7889), .A3(n7888), .Y(n3054) );
  AND3X1_LVT U4934 ( .A1(n7903), .A2(n7902), .A3(n7901), .Y(n3055) );
  AND3X1_LVT U4935 ( .A1(n7886), .A2(n7885), .A3(n7884), .Y(n3056) );
  AND3X1_LVT U4936 ( .A1(n7835), .A2(n7834), .A3(n7833), .Y(n3057) );
  AND3X1_LVT U4937 ( .A1(n7831), .A2(n7830), .A3(n7829), .Y(n3058) );
  AND3X1_LVT U4938 ( .A1(n7848), .A2(n7847), .A3(n7846), .Y(n3059) );
  XNOR2X1_LVT U4939 ( .A1(n4813), .A2(n9390), .Y(n5424) );
  AND3X1_LVT U4940 ( .A1(n7770), .A2(n7769), .A3(n7768), .Y(n3061) );
  AND3X1_LVT U4941 ( .A1(n7783), .A2(n7782), .A3(n7781), .Y(n3062) );
  AND3X1_LVT U4942 ( .A1(n7766), .A2(n7765), .A3(n7764), .Y(n3063) );
  AND3X1_LVT U4943 ( .A1(n7875), .A2(n7874), .A3(n7873), .Y(n3064) );
  AND3X1_LVT U4944 ( .A1(n7859), .A2(n7858), .A3(n7857), .Y(n3065) );
  AND3X1_LVT U4945 ( .A1(n7642), .A2(n7641), .A3(n7640), .Y(n3066) );
  AND3X1_LVT U4946 ( .A1(n7655), .A2(n7654), .A3(n7653), .Y(n3067) );
  AND3X1_LVT U4947 ( .A1(n7638), .A2(n7637), .A3(n7636), .Y(n3068) );
  AND3X1_LVT U4948 ( .A1(n7486), .A2(n7485), .A3(n7484), .Y(n3069) );
  AND3X1_LVT U4949 ( .A1(n7499), .A2(n7498), .A3(n7497), .Y(n3070) );
  AND3X1_LVT U4950 ( .A1(n7482), .A2(n7481), .A3(n7480), .Y(n3071) );
  NAND2X0_LVT U4951 ( .A1(n4844), .A2(n4845), .Y(n3073) );
  NBUFFX2_LVT U4952 ( .A(n9524), .Y(io_fpu_inst[13]) );
  NAND3X2_LVT U4953 ( .A1(n2068), .A2(n6931), .A3(n3709), .Y(n9006) );
  AND3X2_LVT U4954 ( .A1(n6975), .A2(n6931), .A3(n2068), .Y(n3692) );
  AND2X1_LVT U4955 ( .A1(n3044), .A2(n5106), .Y(n9231) );
  INVX1_LVT U4956 ( .A(n9521), .Y(n9438) );
  IBUFFX2_LVT U4957 ( .A(n2981), .Y(n3877) );
  IBUFFX2_LVT U4958 ( .A(n6877), .Y(n3878) );
  MUX21X1_LVT U4959 ( .A1(n5249), .A2(div_io_resp_bits_tag[3]), .S0(n5403), 
        .Y(n5426) );
  MUX21X1_LVT U4960 ( .A1(n5228), .A2(div_io_resp_bits_tag[4]), .S0(n5403), 
        .Y(n5428) );
  MUX21X1_LVT U4961 ( .A1(n5185), .A2(div_io_resp_bits_tag[1]), .S0(n5403), 
        .Y(n5423) );
  MUX21X1_LVT U4962 ( .A1(io_fpu_dmem_resp_tag[0]), .A2(
        div_io_resp_bits_tag[0]), .S0(n5403), .Y(n5306) );
  INVX1_LVT U4963 ( .A(n3883), .Y(n3880) );
  NAND4X1_LVT U4964 ( .A1(n9114), .A2(io_fpu_inst[5]), .A3(n9113), .A4(n9112), 
        .Y(n9115) );
  INVX1_LVT U4965 ( .A(n3803), .Y(n3801) );
  INVX1_LVT U4966 ( .A(n3803), .Y(n3802) );
  INVX1_LVT U4967 ( .A(n3803), .Y(n6764) );
  XOR2X1_LVT U4968 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n9398), .Y(
        n5429) );
  MUX21X1_LVT U4969 ( .A1(n3103), .A2(n5423), .S0(n9381), .Y(n9390) );
  IBUFFX2_LVT U4970 ( .A(n6878), .Y(n3883) );
  IBUFFX2_LVT U4971 ( .A(io_dmem_resp_bits_tag[0]), .Y(n4685) );
  IBUFFX2_LVT U4972 ( .A(n3799), .Y(n3798) );
  IBUFFX2_LVT U4973 ( .A(n9028), .Y(n3717) );
  IBUFFX2_LVT U4974 ( .A(n9028), .Y(n4014) );
  IBUFFX2_LVT U4975 ( .A(n9028), .Y(n3716) );
  NAND3X2_LVT U4976 ( .A1(n6974), .A2(n6973), .A3(n6941), .Y(n9028) );
  IBUFFX2_LVT U4977 ( .A(n2069), .Y(n3744) );
  NBUFFX2_LVT U4978 ( .A(n9518), .Y(n3078) );
  NBUFFX2_LVT U4979 ( .A(n9518), .Y(n3079) );
  INVX1_LVT U4980 ( .A(ibuf_io_inst_0_bits_inst_rs2[1]), .Y(n4813) );
  XOR2X1_LVT U4981 ( .A1(n3781), .A2(n9403), .Y(n5432) );
  IBUFFX2_LVT U4982 ( .A(n9036), .Y(n4017) );
  IBUFFX2_LVT U4983 ( .A(n3012), .Y(n3991) );
  IBUFFX2_LVT U4984 ( .A(n9036), .Y(n4016) );
  IBUFFX2_LVT U4985 ( .A(n2825), .Y(n6956) );
  IBUFFX2_LVT U4986 ( .A(n9523), .Y(n9445) );
  IBUFFX2_LVT U4987 ( .A(n9047), .Y(n3683) );
  IBUFFX2_LVT U4988 ( .A(n9047), .Y(n4053) );
  INVX1_LVT U4989 ( .A(n3658), .Y(n4007) );
  INVX1_LVT U4990 ( .A(n3658), .Y(n4006) );
  INVX1_LVT U4991 ( .A(n3715), .Y(n3747) );
  IBUFFX2_LVT U4992 ( .A(n3012), .Y(n3992) );
  IBUFFX2_LVT U4993 ( .A(n3683), .Y(n3632) );
  IBUFFX2_LVT U4994 ( .A(n3683), .Y(n3656) );
  IBUFFX2_LVT U4995 ( .A(n9529), .Y(n9104) );
  NAND3X2_LVT U4996 ( .A1(n2068), .A2(n6957), .A3(n3709), .Y(n3653) );
  AND3X2_LVT U4997 ( .A1(n3773), .A2(n6948), .A3(n6940), .Y(n9022) );
  IBUFFX2_LVT U4998 ( .A(n6763), .Y(n3799) );
  AND2X1_LVT U4999 ( .A1(n5450), .A2(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(
        n6794) );
  IBUFFX2_LVT U5000 ( .A(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(n3782) );
  IBUFFX2_LVT U5001 ( .A(n4040), .Y(n4036) );
  NBUFFX2_LVT U5002 ( .A(net34650), .Y(n4080) );
  NBUFFX2_LVT U5003 ( .A(net34650), .Y(n4082) );
  NBUFFX2_LVT U5004 ( .A(net34650), .Y(n4084) );
  NBUFFX2_LVT U5005 ( .A(net34650), .Y(n4081) );
  NBUFFX2_LVT U5006 ( .A(net34650), .Y(n4083) );
  NBUFFX2_LVT U5007 ( .A(net34535), .Y(n4223) );
  NBUFFX2_LVT U5008 ( .A(net34575), .Y(n4173) );
  NBUFFX2_LVT U5009 ( .A(net34535), .Y(n4222) );
  NBUFFX2_LVT U5010 ( .A(net34535), .Y(n4219) );
  NBUFFX2_LVT U5011 ( .A(net34535), .Y(n4221) );
  NBUFFX2_LVT U5012 ( .A(net34535), .Y(n4220) );
  NBUFFX2_LVT U5013 ( .A(net34565), .Y(n4183) );
  NBUFFX2_LVT U5014 ( .A(net34525), .Y(n4234) );
  NBUFFX2_LVT U5015 ( .A(net34525), .Y(n4235) );
  NBUFFX2_LVT U5016 ( .A(net34565), .Y(n4184) );
  NBUFFX2_LVT U5017 ( .A(net34565), .Y(n4185) );
  NBUFFX2_LVT U5018 ( .A(net34565), .Y(n4187) );
  NBUFFX2_LVT U5019 ( .A(net34565), .Y(n4186) );
  NBUFFX2_LVT U5020 ( .A(net34575), .Y(n4174) );
  NBUFFX2_LVT U5021 ( .A(net34575), .Y(n4175) );
  NBUFFX2_LVT U5022 ( .A(net34525), .Y(n4231) );
  NBUFFX2_LVT U5023 ( .A(net34570), .Y(n4177) );
  NBUFFX2_LVT U5024 ( .A(net34555), .Y(n4195) );
  NBUFFX2_LVT U5025 ( .A(net34525), .Y(n4232) );
  NBUFFX2_LVT U5026 ( .A(net34570), .Y(n4178) );
  NBUFFX2_LVT U5027 ( .A(net34570), .Y(n4179) );
  NBUFFX2_LVT U5028 ( .A(net34570), .Y(n4180) );
  NBUFFX2_LVT U5029 ( .A(net34525), .Y(n4233) );
  NBUFFX2_LVT U5030 ( .A(net34570), .Y(n4181) );
  NBUFFX2_LVT U5031 ( .A(net34545), .Y(n4210) );
  NBUFFX2_LVT U5032 ( .A(net34615), .Y(n4123) );
  NBUFFX2_LVT U5033 ( .A(net34615), .Y(n4124) );
  NBUFFX2_LVT U5034 ( .A(net34615), .Y(n4125) );
  NBUFFX2_LVT U5035 ( .A(net34555), .Y(n4198) );
  NBUFFX2_LVT U5036 ( .A(net34615), .Y(n4126) );
  NBUFFX2_LVT U5037 ( .A(net34615), .Y(n4127) );
  NBUFFX2_LVT U5038 ( .A(net34555), .Y(n4197) );
  NBUFFX2_LVT U5039 ( .A(net34545), .Y(n4209) );
  NBUFFX2_LVT U5040 ( .A(net34555), .Y(n4196) );
  NBUFFX2_LVT U5041 ( .A(net34605), .Y(n4135) );
  NBUFFX2_LVT U5042 ( .A(net34605), .Y(n4136) );
  NBUFFX2_LVT U5043 ( .A(net34605), .Y(n4137) );
  NBUFFX2_LVT U5044 ( .A(net34635), .Y(n4102) );
  NBUFFX2_LVT U5045 ( .A(net34635), .Y(n4099) );
  NBUFFX2_LVT U5046 ( .A(net34635), .Y(n4103) );
  NBUFFX2_LVT U5047 ( .A(net34545), .Y(n4208) );
  NBUFFX2_LVT U5048 ( .A(net34635), .Y(n4100) );
  NBUFFX2_LVT U5049 ( .A(net34545), .Y(n4207) );
  NBUFFX2_LVT U5050 ( .A(net34625), .Y(n4111) );
  NBUFFX2_LVT U5051 ( .A(net34625), .Y(n4112) );
  NBUFFX2_LVT U5052 ( .A(net34625), .Y(n4113) );
  NBUFFX2_LVT U5053 ( .A(net34625), .Y(n4114) );
  NBUFFX2_LVT U5054 ( .A(net34625), .Y(n4115) );
  NBUFFX2_LVT U5055 ( .A(net34555), .Y(n4199) );
  NBUFFX2_LVT U5056 ( .A(net34545), .Y(n4211) );
  NBUFFX2_LVT U5057 ( .A(net34635), .Y(n4101) );
  NBUFFX2_LVT U5058 ( .A(net34595), .Y(n4151) );
  NBUFFX2_LVT U5059 ( .A(net34645), .Y(n4089) );
  NBUFFX2_LVT U5060 ( .A(net34645), .Y(n4088) );
  NBUFFX2_LVT U5061 ( .A(net34645), .Y(n4087) );
  NBUFFX2_LVT U5062 ( .A(net34645), .Y(n4086) );
  NBUFFX2_LVT U5063 ( .A(net34585), .Y(n4159) );
  NBUFFX2_LVT U5064 ( .A(net34585), .Y(n4160) );
  NBUFFX2_LVT U5065 ( .A(net34585), .Y(n4161) );
  NBUFFX2_LVT U5066 ( .A(net34585), .Y(n4162) );
  NBUFFX2_LVT U5067 ( .A(net34585), .Y(n4163) );
  NBUFFX2_LVT U5068 ( .A(net34575), .Y(n4171) );
  NBUFFX2_LVT U5069 ( .A(net34575), .Y(n4172) );
  NBUFFX2_LVT U5070 ( .A(net34595), .Y(n4150) );
  NBUFFX2_LVT U5071 ( .A(net34595), .Y(n4149) );
  NBUFFX2_LVT U5072 ( .A(net34595), .Y(n4148) );
  NBUFFX2_LVT U5073 ( .A(net34645), .Y(n4090) );
  NBUFFX2_LVT U5074 ( .A(net34605), .Y(n4138) );
  NBUFFX2_LVT U5075 ( .A(net34605), .Y(n4139) );
  NBUFFX2_LVT U5076 ( .A(net34595), .Y(n4147) );
  NBUFFX2_LVT U5077 ( .A(net34640), .Y(n4098) );
  NAND3X0_LVT U5078 ( .A1(n9244), .A2(n9243), .A3(n9242), .Y(n9245) );
  NBUFFX2_LVT U5079 ( .A(net34540), .Y(n4217) );
  NBUFFX2_LVT U5080 ( .A(net34540), .Y(n4216) );
  NBUFFX2_LVT U5081 ( .A(net34655), .Y(n4078) );
  NBUFFX2_LVT U5082 ( .A(net34520), .Y(n4239) );
  NBUFFX2_LVT U5083 ( .A(net34540), .Y(n4215) );
  NBUFFX2_LVT U5084 ( .A(net34540), .Y(n4214) );
  NBUFFX2_LVT U5085 ( .A(net34530), .Y(n4228) );
  NBUFFX2_LVT U5086 ( .A(net34530), .Y(n4227) );
  NBUFFX2_LVT U5087 ( .A(net34530), .Y(n4226) );
  NBUFFX2_LVT U5088 ( .A(net34530), .Y(n4229) );
  NBUFFX2_LVT U5089 ( .A(net34530), .Y(n4225) );
  NBUFFX2_LVT U5090 ( .A(net34655), .Y(n4076) );
  NBUFFX2_LVT U5091 ( .A(net34655), .Y(n4074) );
  NBUFFX2_LVT U5092 ( .A(net34520), .Y(n4241) );
  NBUFFX2_LVT U5093 ( .A(net34655), .Y(n4077) );
  NBUFFX2_LVT U5094 ( .A(net34655), .Y(n4075) );
  NBUFFX2_LVT U5095 ( .A(net34560), .Y(n4190) );
  NBUFFX2_LVT U5096 ( .A(net34600), .Y(n4145) );
  NBUFFX2_LVT U5097 ( .A(net34560), .Y(n4191) );
  NBUFFX2_LVT U5098 ( .A(net34600), .Y(n4144) );
  NBUFFX2_LVT U5099 ( .A(net34600), .Y(n4143) );
  NBUFFX2_LVT U5100 ( .A(net34560), .Y(n4192) );
  NBUFFX2_LVT U5101 ( .A(net34600), .Y(n4142) );
  NBUFFX2_LVT U5102 ( .A(net34600), .Y(n4141) );
  NBUFFX2_LVT U5103 ( .A(net34560), .Y(n4193) );
  NBUFFX2_LVT U5104 ( .A(net34610), .Y(n4133) );
  NBUFFX2_LVT U5105 ( .A(net34610), .Y(n4132) );
  NBUFFX2_LVT U5106 ( .A(net34610), .Y(n4131) );
  NBUFFX2_LVT U5107 ( .A(net34580), .Y(n4167) );
  NBUFFX2_LVT U5108 ( .A(net34580), .Y(n4166) );
  NBUFFX2_LVT U5109 ( .A(net34580), .Y(n4165) );
  NBUFFX2_LVT U5110 ( .A(net34630), .Y(n4105) );
  NBUFFX2_LVT U5111 ( .A(net34630), .Y(n4106) );
  NBUFFX2_LVT U5112 ( .A(net34580), .Y(n4169) );
  NBUFFX2_LVT U5113 ( .A(net34580), .Y(n4168) );
  NBUFFX2_LVT U5114 ( .A(net34630), .Y(n4107) );
  NBUFFX2_LVT U5115 ( .A(net34520), .Y(n4240) );
  NBUFFX2_LVT U5116 ( .A(net34590), .Y(n4157) );
  NBUFFX2_LVT U5117 ( .A(net34590), .Y(n4156) );
  NBUFFX2_LVT U5118 ( .A(net34590), .Y(n4155) );
  NBUFFX2_LVT U5119 ( .A(net34630), .Y(n4108) );
  NBUFFX2_LVT U5120 ( .A(net34590), .Y(n4154) );
  NBUFFX2_LVT U5121 ( .A(net34520), .Y(n4238) );
  NBUFFX2_LVT U5122 ( .A(net34630), .Y(n4109) );
  NBUFFX2_LVT U5123 ( .A(net34560), .Y(n4189) );
  NBUFFX2_LVT U5124 ( .A(net34590), .Y(n4153) );
  NBUFFX2_LVT U5125 ( .A(net34520), .Y(n4237) );
  NBUFFX2_LVT U5126 ( .A(net34550), .Y(n4204) );
  NBUFFX2_LVT U5127 ( .A(net34620), .Y(n4119) );
  NBUFFX2_LVT U5128 ( .A(net34550), .Y(n4202) );
  NBUFFX2_LVT U5129 ( .A(net34550), .Y(n4203) );
  NBUFFX2_LVT U5130 ( .A(net34620), .Y(n4120) );
  NBUFFX2_LVT U5131 ( .A(net34620), .Y(n4121) );
  NBUFFX2_LVT U5132 ( .A(net34540), .Y(n4213) );
  NBUFFX2_LVT U5133 ( .A(net34610), .Y(n4130) );
  NBUFFX2_LVT U5134 ( .A(net34610), .Y(n4129) );
  NBUFFX2_LVT U5135 ( .A(net34620), .Y(n4117) );
  NBUFFX2_LVT U5136 ( .A(net34550), .Y(n4201) );
  NBUFFX2_LVT U5137 ( .A(net34550), .Y(n4205) );
  NBUFFX2_LVT U5138 ( .A(net34620), .Y(n4118) );
  NBUFFX2_LVT U5139 ( .A(net34640), .Y(n4093) );
  NBUFFX2_LVT U5140 ( .A(net34640), .Y(n4095) );
  NBUFFX2_LVT U5141 ( .A(net34640), .Y(n4094) );
  NBUFFX2_LVT U5142 ( .A(net34640), .Y(n4096) );
  NBUFFX2_LVT U5143 ( .A(net34640), .Y(n4097) );
  NBUFFX2_LVT U5144 ( .A(net34640), .Y(n4092) );
  MUX21X1_LVT U5145 ( .A1(n9252), .A2(wb_cause[3]), .S0(wb_cause[1]), .Y(n9255) );
  INVX1_LVT U5146 ( .A(n5260), .Y(n5287) );
  OR2X1_LVT U5147 ( .A1(n5259), .A2(n5270), .Y(n5276) );
  OR2X1_LVT U5148 ( .A1(n5259), .A2(n5280), .Y(n5266) );
  INVX1_LVT U5149 ( .A(n9164), .Y(n9144) );
  OR2X1_LVT U5150 ( .A1(io_fpu_dmem_resp_tag[2]), .A2(n5244), .Y(n5237) );
  NBUFFX2_LVT U5151 ( .A(n711), .Y(n4066) );
  NBUFFX2_LVT U5152 ( .A(n711), .Y(n4067) );
  NBUFFX2_LVT U5153 ( .A(n_T_427__T_1136_data[16]), .Y(n4362) );
  NBUFFX2_LVT U5154 ( .A(n_T_427__T_1136_data[16]), .Y(n4363) );
  NBUFFX2_LVT U5155 ( .A(n_T_427__T_1136_data[54]), .Y(n4468) );
  NBUFFX2_LVT U5156 ( .A(n_T_427__T_1136_data[54]), .Y(n4467) );
  NBUFFX2_LVT U5157 ( .A(n_T_427__T_1136_data[36]), .Y(n4415) );
  NBUFFX2_LVT U5158 ( .A(n_T_427__T_1136_data[36]), .Y(n4414) );
  NBUFFX2_LVT U5159 ( .A(n_T_427__T_1136_data[49]), .Y(n4453) );
  NBUFFX2_LVT U5160 ( .A(n_T_427__T_1136_data[52]), .Y(n4462) );
  NBUFFX2_LVT U5161 ( .A(n_T_427__T_1136_data[56]), .Y(n4474) );
  NBUFFX2_LVT U5162 ( .A(n_T_427__T_1136_data[29]), .Y(n4396) );
  NBUFFX2_LVT U5163 ( .A(n_T_427__T_1136_data[30]), .Y(n4399) );
  NBUFFX2_LVT U5164 ( .A(n_T_427__T_1136_data[49]), .Y(n4452) );
  NBUFFX2_LVT U5165 ( .A(n_T_427__T_1136_data[41]), .Y(n4429) );
  NBUFFX2_LVT U5166 ( .A(n_T_427__T_1136_data[29]), .Y(n4397) );
  NBUFFX2_LVT U5167 ( .A(n_T_427__T_1136_data[56]), .Y(n4473) );
  NBUFFX2_LVT U5168 ( .A(n_T_427__T_1136_data[30]), .Y(n4400) );
  NBUFFX2_LVT U5169 ( .A(n_T_427__T_1136_data[41]), .Y(n4428) );
  NBUFFX2_LVT U5170 ( .A(n_T_427__T_1136_data[52]), .Y(n4461) );
  NBUFFX2_LVT U5171 ( .A(n_T_427__T_1136_data[27]), .Y(n4391) );
  NBUFFX2_LVT U5172 ( .A(n_T_427__T_1136_data[27]), .Y(n4392) );
  NBUFFX2_LVT U5173 ( .A(n_T_427__T_1136_data[58]), .Y(n4480) );
  NBUFFX2_LVT U5174 ( .A(n_T_427__T_1136_data[58]), .Y(n4479) );
  NBUFFX2_LVT U5175 ( .A(n_T_427__T_1136_data[62]), .Y(n4491) );
  NBUFFX2_LVT U5176 ( .A(n_T_427__T_1136_data[60]), .Y(n4485) );
  NBUFFX2_LVT U5177 ( .A(n_T_427__T_1136_data[62]), .Y(n4492) );
  NBUFFX2_LVT U5178 ( .A(n_T_427__T_1136_data[60]), .Y(n4486) );
  NBUFFX2_LVT U5179 ( .A(n_T_427__T_1136_data[53]), .Y(n4465) );
  NBUFFX2_LVT U5180 ( .A(n_T_427__T_1136_data[53]), .Y(n4464) );
  NBUFFX2_LVT U5181 ( .A(n_T_427__T_1136_data[59]), .Y(n4483) );
  NBUFFX2_LVT U5182 ( .A(n_T_427__T_1136_data[59]), .Y(n4482) );
  NBUFFX2_LVT U5183 ( .A(n_T_427__T_1136_data[1]), .Y(n4320) );
  NBUFFX2_LVT U5184 ( .A(n_T_427__T_1136_data[1]), .Y(n4319) );
  NBUFFX2_LVT U5185 ( .A(n_T_427__T_1136_data[50]), .Y(n4456) );
  NBUFFX2_LVT U5186 ( .A(n_T_427__T_1136_data[50]), .Y(n4455) );
  NBUFFX2_LVT U5187 ( .A(n_T_427__T_1136_data[61]), .Y(n4489) );
  NBUFFX2_LVT U5188 ( .A(n_T_427__T_1136_data[61]), .Y(n4488) );
  NBUFFX2_LVT U5189 ( .A(n_T_427__T_1136_data[57]), .Y(n4477) );
  NBUFFX2_LVT U5190 ( .A(n_T_427__T_1136_data[55]), .Y(n4470) );
  NBUFFX2_LVT U5191 ( .A(n_T_427__T_1136_data[55]), .Y(n4471) );
  NBUFFX2_LVT U5192 ( .A(n_T_427__T_1136_data[57]), .Y(n4476) );
  NBUFFX2_LVT U5193 ( .A(n_T_427__T_1136_data[19]), .Y(n4372) );
  NBUFFX2_LVT U5194 ( .A(n_T_427__T_1136_data[20]), .Y(n4375) );
  NBUFFX2_LVT U5195 ( .A(n_T_427__T_1136_data[19]), .Y(n4371) );
  NBUFFX2_LVT U5196 ( .A(n_T_427__T_1136_data[24]), .Y(n4385) );
  NBUFFX2_LVT U5197 ( .A(n_T_427__T_1136_data[0]), .Y(n4317) );
  NBUFFX2_LVT U5198 ( .A(n_T_427__T_1136_data[24]), .Y(n4384) );
  NBUFFX2_LVT U5199 ( .A(n_T_427__T_1136_data[0]), .Y(n4316) );
  NBUFFX2_LVT U5200 ( .A(n_T_427__T_1136_data[18]), .Y(n4368) );
  NBUFFX2_LVT U5201 ( .A(n_T_427__T_1136_data[18]), .Y(n4369) );
  NBUFFX2_LVT U5202 ( .A(n_T_427__T_1136_data[20]), .Y(n4374) );
  NBUFFX2_LVT U5203 ( .A(n_T_427__T_1136_data[63]), .Y(n4495) );
  NBUFFX2_LVT U5204 ( .A(n_T_427__T_1136_data[63]), .Y(n4494) );
  NBUFFX2_LVT U5205 ( .A(n_T_427__T_1136_data[37]), .Y(n4417) );
  NBUFFX2_LVT U5206 ( .A(n_T_427__T_1136_data[37]), .Y(n4418) );
  NBUFFX2_LVT U5207 ( .A(n_T_427__T_1136_data[44]), .Y(n4437) );
  NBUFFX2_LVT U5208 ( .A(n_T_427__T_1136_data[32]), .Y(n4404) );
  NBUFFX2_LVT U5209 ( .A(n_T_427__T_1136_data[34]), .Y(n4410) );
  NBUFFX2_LVT U5210 ( .A(n_T_427__T_1136_data[46]), .Y(n4444) );
  NBUFFX2_LVT U5211 ( .A(n_T_427__T_1136_data[46]), .Y(n4443) );
  NBUFFX2_LVT U5212 ( .A(n_T_427__T_1136_data[39]), .Y(n4423) );
  NBUFFX2_LVT U5213 ( .A(n_T_427__T_1136_data[32]), .Y(n4405) );
  NBUFFX2_LVT U5214 ( .A(n_T_427__T_1136_data[44]), .Y(n4438) );
  NBUFFX2_LVT U5215 ( .A(n_T_427__T_1136_data[34]), .Y(n4409) );
  NBUFFX2_LVT U5216 ( .A(n_T_427__T_1136_data[39]), .Y(n4422) );
  NBUFFX2_LVT U5217 ( .A(n_T_427__T_1136_data[17]), .Y(n4365) );
  NBUFFX2_LVT U5218 ( .A(n_T_427__T_1136_data[23]), .Y(n4381) );
  NBUFFX2_LVT U5219 ( .A(n_T_427__T_1136_data[23]), .Y(n4382) );
  NBUFFX2_LVT U5220 ( .A(n_T_427__T_1136_data[17]), .Y(n4366) );
  NBUFFX2_LVT U5221 ( .A(n_T_427__T_1136_data[40]), .Y(n4425) );
  NBUFFX2_LVT U5222 ( .A(n_T_427__T_1136_data[47]), .Y(n4447) );
  NBUFFX2_LVT U5223 ( .A(n_T_427__T_1136_data[48]), .Y(n4450) );
  NBUFFX2_LVT U5224 ( .A(n_T_427__T_1136_data[48]), .Y(n4449) );
  NBUFFX2_LVT U5225 ( .A(n_T_427__T_1136_data[47]), .Y(n4446) );
  NBUFFX2_LVT U5226 ( .A(n_T_427__T_1136_data[40]), .Y(n4426) );
  NBUFFX2_LVT U5227 ( .A(n_T_427__T_1136_data[45]), .Y(n4441) );
  NBUFFX2_LVT U5228 ( .A(n_T_427__T_1136_data[45]), .Y(n4440) );
  NBUFFX2_LVT U5229 ( .A(n_T_427__T_1136_data[51]), .Y(n4458) );
  NBUFFX2_LVT U5230 ( .A(n_T_427__T_1136_data[43]), .Y(n4434) );
  NBUFFX2_LVT U5231 ( .A(n_T_427__T_1136_data[42]), .Y(n4431) );
  NBUFFX2_LVT U5232 ( .A(n_T_427__T_1136_data[51]), .Y(n4459) );
  NBUFFX2_LVT U5233 ( .A(n_T_427__T_1136_data[43]), .Y(n4435) );
  NBUFFX2_LVT U5234 ( .A(n_T_427__T_1136_data[42]), .Y(n4432) );
  AND3X1_LVT U5235 ( .A1(io_imem_bht_update_bits_mispredict), .A2(
        io_imem_bht_update_valid), .A3(n9329), .Y(io_imem_btb_update_valid) );
  NAND3X0_LVT U5236 ( .A1(n9231), .A2(n2618), .A3(n9079), .Y(n9080) );
  XOR2X1_LVT U5237 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n591), .Y(n5032)
         );
  XOR2X1_LVT U5238 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n589), .Y(n5030)
         );
  XOR2X1_LVT U5239 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n592), .Y(n5035)
         );
  XOR2X1_LVT U5240 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n3201), .Y(n5017) );
  XOR2X1_LVT U5241 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n3103), .Y(n5018) );
  XOR2X1_LVT U5242 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n3199), .Y(n5014) );
  XOR2X1_LVT U5243 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n3198), .Y(n5015) );
  XOR2X1_LVT U5244 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n3102), .Y(n5016) );
  NAND4X0_LVT U5245 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n5437), .Y(n4910) );
  NAND4X0_LVT U5246 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n5437), .Y(n4914) );
  OA21X1_LVT U5247 ( .A1(n3264), .A2(n6422), .A3(n5434), .Y(n4883) );
  MUX21X1_LVT U5248 ( .A1(n4812), .A2(n4811), .S0(
        ibuf_io_inst_0_bits_inst_rs3_4_), .Y(n4839) );
  NAND2X0_LVT U5249 ( .A1(n4782), .A2(ibuf_io_inst_0_bits_raw[27]), .Y(n4803)
         );
  NAND2X0_LVT U5250 ( .A1(n4781), .A2(ibuf_io_inst_0_bits_raw[28]), .Y(n4801)
         );
  XOR2X1_LVT U5251 ( .A1(ibuf_io_inst_0_bits_inst_rs3_2_), .A2(n3200), .Y(
        n4624) );
  XOR2X1_LVT U5252 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n596), .Y(n4619)
         );
  XOR2X1_LVT U5253 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n595), .Y(n4620)
         );
  XOR2X1_LVT U5254 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n3200), .Y(n4621) );
  INVX1_LVT U5255 ( .A(ibuf_io_pc[34]), .Y(n4557) );
  XOR2X1_LVT U5256 ( .A1(n9484), .A2(ibuf_io_pc[5]), .Y(n4541) );
  XOR2X1_LVT U5257 ( .A1(n9334), .A2(n4532), .Y(n4535) );
  XOR2X1_LVT U5258 ( .A1(n9503), .A2(ibuf_io_pc[3]), .Y(n4537) );
  XOR2X1_LVT U5259 ( .A1(n9499), .A2(ibuf_io_pc[7]), .Y(n4543) );
  INVX1_LVT U5260 ( .A(ibuf_io_pc[16]), .Y(n4518) );
  NBUFFX2_LVT U5261 ( .A(n711), .Y(n4065) );
  OR2X1_LVT U5262 ( .A1(csr_io_exception), .A2(csr_io_eret), .Y(n711) );
  NBUFFX2_LVT U5263 ( .A(n6898), .Y(n3957) );
  NBUFFX2_LVT U5264 ( .A(n6886), .Y(n3908) );
  NBUFFX2_LVT U5265 ( .A(n6838), .Y(n3840) );
  NBUFFX2_LVT U5266 ( .A(n6865), .Y(n3859) );
  NBUFFX2_LVT U5267 ( .A(n6868), .Y(n3867) );
  NBUFFX2_LVT U5268 ( .A(n6870), .Y(n3871) );
  NBUFFX2_LVT U5269 ( .A(n6898), .Y(n3958) );
  INVX1_LVT U5270 ( .A(n5546), .Y(n6870) );
  INVX1_LVT U5271 ( .A(n4814), .Y(n4901) );
  NAND2X0_LVT U5272 ( .A1(n5452), .A2(n2878), .Y(n3083) );
  NBUFFX2_LVT U5273 ( .A(n6715), .Y(n3796) );
  NBUFFX2_LVT U5274 ( .A(n6869), .Y(n3868) );
  NBUFFX2_LVT U5275 ( .A(n6837), .Y(n3836) );
  NAND2X0_LVT U5276 ( .A1(n5449), .A2(n5436), .Y(n6766) );
  NBUFFX2_LVT U5277 ( .A(n6795), .Y(n3812) );
  AND2X1_LVT U5278 ( .A1(n4027), .A2(n2135), .Y(n3661) );
  NBUFFX2_LVT U5279 ( .A(n9038), .Y(n4027) );
  NBUFFX2_LVT U5280 ( .A(n8900), .Y(n3960) );
  NBUFFX2_LVT U5281 ( .A(n8981), .Y(n3979) );
  NBUFFX2_LVT U5282 ( .A(n8932), .Y(n3972) );
  NBUFFX2_LVT U5283 ( .A(n8931), .Y(n3968) );
  NBUFFX2_LVT U5284 ( .A(n8982), .Y(n3983) );
  NBUFFX2_LVT U5285 ( .A(n8980), .Y(n3976) );
  NAND2X0_LVT U5286 ( .A1(n6939), .A2(n6936), .Y(n3625) );
  NBUFFX2_LVT U5287 ( .A(n9042), .Y(n4051) );
  INVX1_LVT U5288 ( .A(n3184), .Y(n4026) );
  INVX1_LVT U5289 ( .A(n6945), .Y(n9042) );
  INVX1_LVT U5290 ( .A(n4017), .Y(n4015) );
  XOR2X1_LVT U5291 ( .A1(ibuf_io_inst_0_bits_inst_rs1[3]), .A2(n9403), .Y(
        n6908) );
  XOR2X1_LVT U5292 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n9398), .Y(
        n6909) );
  XOR2X1_LVT U5293 ( .A1(n3040), .A2(n2098), .Y(n6910) );
  XOR2X1_LVT U5294 ( .A1(n3042), .A2(n2038), .Y(n6911) );
  XOR2X1_LVT U5295 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n588), .Y(n5010) );
  XOR2X1_LVT U5296 ( .A1(ibuf_io_inst_0_bits_inst_rs1[2]), .A2(n590), .Y(n5012) );
  XOR2X1_LVT U5297 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n595), .Y(n4617) );
  OAI21X1_LVT U5298 ( .A1(n2618), .A2(n3079), .A3(n9522), .Y(n3180) );
  XOR2X1_LVT U5299 ( .A1(n9495), .A2(ibuf_io_pc[4]), .Y(n4540) );
  INVX1_LVT U5300 ( .A(ibuf_io_pc[2]), .Y(n4532) );
  XOR2X1_LVT U5301 ( .A1(n9512), .A2(ibuf_io_pc[1]), .Y(n4534) );
  NBUFFX2_LVT U5302 ( .A(n8901), .Y(n3964) );
  OA22X1_LVT U5303 ( .A1(n3269), .A2(n5906), .A3(n3128), .A4(n5905), .Y(n4882)
         );
  AO22X1_LVT U5304 ( .A1(n_T_698[3]), .A2(n9101), .A3(io_fpu_fromint_data[3]), 
        .A4(n9103), .Y(alu_io_in1[3]) );
  AO22X1_LVT U5305 ( .A1(n_T_698[4]), .A2(n9101), .A3(io_fpu_fromint_data[4]), 
        .A4(n9103), .Y(alu_io_in1[4]) );
  AO22X1_LVT U5306 ( .A1(n_T_698[2]), .A2(n4054), .A3(io_fpu_fromint_data[2]), 
        .A4(n9103), .Y(alu_io_in1[2]) );
  AO22X1_LVT U5307 ( .A1(n_T_698[6]), .A2(n4054), .A3(io_fpu_fromint_data[6]), 
        .A4(n9103), .Y(alu_io_in1[6]) );
  AO22X1_LVT U5308 ( .A1(n_T_698[0]), .A2(n9101), .A3(io_fpu_fromint_data[0]), 
        .A4(n9103), .Y(alu_io_in1[0]) );
  AO22X1_LVT U5309 ( .A1(n_T_698[7]), .A2(n4054), .A3(io_fpu_fromint_data[7]), 
        .A4(n9103), .Y(alu_io_in1[7]) );
  AO22X1_LVT U5310 ( .A1(n_T_698[10]), .A2(n4054), .A3(io_fpu_fromint_data[10]), .A4(n9103), .Y(alu_io_in1[10]) );
  AO22X1_LVT U5311 ( .A1(n_T_698[12]), .A2(n4054), .A3(io_fpu_fromint_data[12]), .A4(n9103), .Y(alu_io_in1[12]) );
  AO22X1_LVT U5312 ( .A1(n_T_698[13]), .A2(n4054), .A3(io_fpu_fromint_data[13]), .A4(n9103), .Y(alu_io_in1[13]) );
  AO22X1_LVT U5313 ( .A1(n_T_698[14]), .A2(n4054), .A3(io_fpu_fromint_data[14]), .A4(n9103), .Y(alu_io_in1[14]) );
  AO22X1_LVT U5314 ( .A1(n_T_698[15]), .A2(n4054), .A3(io_fpu_fromint_data[15]), .A4(n9103), .Y(alu_io_in1[15]) );
  AO22X1_LVT U5315 ( .A1(n_T_698[16]), .A2(n4054), .A3(io_fpu_fromint_data[16]), .A4(n9103), .Y(alu_io_in1[16]) );
  AO22X1_LVT U5316 ( .A1(n4054), .A2(n_T_698[17]), .A3(io_fpu_fromint_data[17]), .A4(n9103), .Y(alu_io_in1[17]) );
  AO22X1_LVT U5317 ( .A1(n_T_698[18]), .A2(n4054), .A3(io_fpu_fromint_data[18]), .A4(n9103), .Y(alu_io_in1[18]) );
  AO22X1_LVT U5318 ( .A1(n_T_698[19]), .A2(n4054), .A3(io_fpu_fromint_data[19]), .A4(n9103), .Y(alu_io_in1[19]) );
  AO22X1_LVT U5319 ( .A1(n9101), .A2(n_T_698[20]), .A3(io_fpu_fromint_data[20]), .A4(n9103), .Y(alu_io_in1[20]) );
  AO22X1_LVT U5320 ( .A1(n_T_698[21]), .A2(n9101), .A3(io_fpu_fromint_data[21]), .A4(n9103), .Y(alu_io_in1[21]) );
  AO22X1_LVT U5321 ( .A1(n_T_698[22]), .A2(n9101), .A3(io_fpu_fromint_data[22]), .A4(n9103), .Y(alu_io_in1[22]) );
  AO22X1_LVT U5322 ( .A1(n_T_698[29]), .A2(n4054), .A3(io_fpu_fromint_data[29]), .A4(n9103), .Y(alu_io_in1[29]) );
  AO22X1_LVT U5323 ( .A1(n9101), .A2(n_T_698[30]), .A3(io_fpu_fromint_data[30]), .A4(n9103), .Y(alu_io_in1[30]) );
  AO22X1_LVT U5324 ( .A1(n_T_698[23]), .A2(n9101), .A3(io_fpu_fromint_data[23]), .A4(n9103), .Y(alu_io_in1[23]) );
  AO22X1_LVT U5325 ( .A1(n_T_698[24]), .A2(n9101), .A3(io_fpu_fromint_data[24]), .A4(n9103), .Y(alu_io_in1[24]) );
  AO22X1_LVT U5326 ( .A1(n4054), .A2(n_T_698[33]), .A3(io_fpu_fromint_data[33]), .A4(n9103), .Y(alu_io_in1[33]) );
  AO22X1_LVT U5327 ( .A1(n_T_698[35]), .A2(n9101), .A3(io_fpu_fromint_data[35]), .A4(n9103), .Y(alu_io_in1[35]) );
  AO22X1_LVT U5328 ( .A1(n_T_698[32]), .A2(n9101), .A3(io_fpu_fromint_data[32]), .A4(n9103), .Y(alu_io_in1[32]) );
  AO22X1_LVT U5329 ( .A1(n_T_698[34]), .A2(n4054), .A3(io_fpu_fromint_data[34]), .A4(n9103), .Y(alu_io_in1[34]) );
  AO22X1_LVT U5330 ( .A1(n4054), .A2(n_T_698[36]), .A3(io_fpu_fromint_data[36]), .A4(n9103), .Y(alu_io_in1[36]) );
  AO22X1_LVT U5331 ( .A1(n9101), .A2(n_T_698[37]), .A3(io_fpu_fromint_data[37]), .A4(n9103), .Y(alu_io_in1[37]) );
  AO22X1_LVT U5332 ( .A1(n4054), .A2(n_T_698[38]), .A3(io_fpu_fromint_data[38]), .A4(n9103), .Y(alu_io_in1[38]) );
  NAND2X0_LVT U5333 ( .A1(mem_br_target_39_), .A2(n6249), .Y(n6857) );
  AND2X1_LVT U5334 ( .A1(n5409), .A2(n5410), .Y(n6855) );
  INVX1_LVT U5335 ( .A(n5410), .Y(n6856) );
  AND2X1_LVT U5336 ( .A1(n5407), .A2(n5406), .Y(n6249) );
  INVX1_LVT U5337 ( .A(n9292), .Y(n9301) );
  INVX1_LVT U5338 ( .A(n3234), .Y(n4058) );
  NAND2X0_LVT U5339 ( .A1(io_dmem_req_bits_size[0]), .A2(
        io_dmem_req_bits_size[1]), .Y(n3234) );
  NOR2X0_LVT U5340 ( .A1(io_dmem_req_bits_size[1]), .A2(
        io_dmem_req_bits_size[0]), .Y(n9291) );
  OR2X1_LVT U5341 ( .A1(io_fpu_sboard_clra[4]), .A2(io_fpu_sboard_clra[3]), 
        .Y(n5193) );
  MUX21X1_LVT U5342 ( .A1(n7016), .A2(io_fpu_dmem_resp_data[0]), .S0(n9064), 
        .Y(io_fpu_fromint_data[0]) );
  OR2X1_LVT U5343 ( .A1(n9201), .A2(n9173), .Y(n9164) );
  OR2X1_LVT U5344 ( .A1(n9201), .A2(n9172), .Y(n9163) );
  OR2X1_LVT U5345 ( .A1(ex_ctrl_sel_imm[2]), .A2(n546), .Y(n9178) );
  AND3X1_LVT U5346 ( .A1(n9173), .A2(n9179), .A3(ex_reg_inst_31_), .Y(n9226)
         );
  AND2X1_LVT U5347 ( .A1(n9101), .A2(n_T_698[39]), .Y(n9102) );
  NOR2X0_LVT U5348 ( .A1(ex_ctrl_sel_alu1_0_), .A2(n561), .Y(n9101) );
  AND2X1_LVT U5349 ( .A1(n561), .A2(ex_ctrl_sel_alu1_0_), .Y(n9103) );
  MUX21X1_LVT U5350 ( .A1(io_fpu_inst[3]), .A2(io_fpu_inst[2]), .S0(n2553), 
        .Y(id_ctrl_sel_imm[1]) );
  INVX1_LVT U5351 ( .A(n5282), .Y(n5381) );
  INVX1_LVT U5352 ( .A(n5272), .Y(n5365) );
  AND2X1_LVT U5353 ( .A1(n5210), .A2(n3043), .Y(n5317) );
  AND2X1_LVT U5354 ( .A1(n5227), .A2(wb_waddr[3]), .Y(n5382) );
  INVX1_LVT U5355 ( .A(n5298), .Y(n5362) );
  INVX1_LVT U5356 ( .A(ex_reg_rs_bypass_1), .Y(n6901) );
  AND2X1_LVT U5357 ( .A1(n5484), .A2(ex_reg_rs_bypass_1), .Y(n6900) );
  AND2X1_LVT U5358 ( .A1(n7017), .A2(n569), .Y(n9065) );
  OR2X1_LVT U5359 ( .A1(mem_reg_xcpt), .A2(mem_reg_xcpt_interrupt), .Y(n1279)
         );
  MUX21X1_LVT U5360 ( .A1(io_fpu_inst[13]), .A2(n5421), .S0(n9287), .Y(N370)
         );
  MUX21X1_LVT U5361 ( .A1(n2618), .A2(n9288), .S0(n9287), .Y(N369) );
  MUX21X1_LVT U5362 ( .A1(n3226), .A2(n4592), .S0(n3792), .Y(n9505) );
  MUX21X1_LVT U5363 ( .A1(n3219), .A2(n4586), .S0(n3792), .Y(n9492) );
  MUX21X1_LVT U5364 ( .A1(n3110), .A2(n4581), .S0(n3792), .Y(n9497) );
  MUX21X1_LVT U5365 ( .A1(n3210), .A2(n4580), .S0(n4591), .Y(n9493) );
  MUX21X1_LVT U5366 ( .A1(n3216), .A2(n4579), .S0(n3792), .Y(n9501) );
  MUX21X1_LVT U5367 ( .A1(n3224), .A2(n4578), .S0(n3792), .Y(n9486) );
  MUX21X1_LVT U5368 ( .A1(n_T_918[28]), .A2(mem_br_target_28_), .S0(n3792), 
        .Y(n9368) );
  MUX21X1_LVT U5369 ( .A1(n_T_918[24]), .A2(mem_br_target_24_), .S0(n3792), 
        .Y(n9364) );
  MUX21X1_LVT U5370 ( .A1(n4573), .A2(mem_br_target_39_), .S0(n3792), .Y(n9377) );
  MUX21X1_LVT U5371 ( .A1(n3212), .A2(n4572), .S0(n3792), .Y(n9510) );
  MUX21X1_LVT U5372 ( .A1(n_T_918[21]), .A2(mem_br_target_21_), .S0(n3792), 
        .Y(n9361) );
  MUX21X1_LVT U5373 ( .A1(n3211), .A2(n4571), .S0(n3792), .Y(n9490) );
  MUX21X1_LVT U5374 ( .A1(n3106), .A2(n4570), .S0(n3792), .Y(n9500) );
  MUX21X1_LVT U5375 ( .A1(n3225), .A2(n4569), .S0(n3792), .Y(n9509) );
  MUX21X1_LVT U5376 ( .A1(n_T_918[15]), .A2(mem_br_target_15_), .S0(n3792), 
        .Y(n9355) );
  MUX21X1_LVT U5377 ( .A1(n3111), .A2(n4568), .S0(n3792), .Y(n9504) );
  MUX21X1_LVT U5378 ( .A1(n3528), .A2(n4567), .S0(n3792), .Y(n9494) );
  MUX21X1_LVT U5379 ( .A1(n3105), .A2(n4562), .S0(n4591), .Y(n9502) );
  MUX21X1_LVT U5380 ( .A1(n_T_918[34]), .A2(mem_br_target_34_), .S0(n3792), 
        .Y(n9373) );
  MUX21X1_LVT U5381 ( .A1(n3107), .A2(n4550), .S0(n4591), .Y(n9487) );
  MUX21X1_LVT U5382 ( .A1(n3207), .A2(n4533), .S0(n4591), .Y(n9512) );
  MUX21X1_LVT U5383 ( .A1(n3221), .A2(n4527), .S0(n4591), .Y(n9491) );
  MUX21X1_LVT U5384 ( .A1(n3223), .A2(n4526), .S0(n3792), .Y(n9506) );
  MUX21X1_LVT U5385 ( .A1(n3220), .A2(n4525), .S0(n4591), .Y(n9496) );
  MUX21X1_LVT U5386 ( .A1(n3213), .A2(n4524), .S0(n3792), .Y(n9488) );
  MUX21X1_LVT U5387 ( .A1(n3209), .A2(n4523), .S0(n4591), .Y(n9489) );
  MUX21X1_LVT U5388 ( .A1(n3227), .A2(n4522), .S0(n3792), .Y(n9508) );
  MUX21X1_LVT U5389 ( .A1(n3218), .A2(n4517), .S0(n3792), .Y(n9483) );
  NBUFFX2_LVT U5390 ( .A(n4591), .Y(n3792) );
  MUX21X1_LVT U5391 ( .A1(n3205), .A2(n4516), .S0(n4591), .Y(n9498) );
  AND2X1_LVT U5392 ( .A1(n3230), .A2(n5080), .Y(n5083) );
  AND2X1_LVT U5393 ( .A1(n_T_844_10_), .A2(n5082), .Y(n9427) );
  NAND3X2_LVT U5394 ( .A1(n2068), .A2(n6972), .A3(n3709), .Y(n3684) );
  NAND3X2_LVT U5395 ( .A1(n6975), .A2(n6957), .A3(n2068), .Y(n3658) );
  NAND3X2_LVT U5396 ( .A1(n3773), .A2(n6954), .A3(n2068), .Y(n3601) );
  OR2X2_LVT U5397 ( .A1(n9113), .A2(n9104), .Y(n1699) );
  OR2X2_LVT U5398 ( .A1(n4848), .A2(n4847), .Y(n6991) );
  NAND2X0_LVT U5399 ( .A1(n5408), .A2(n3251), .Y(n5410) );
  NBUFFX2_LVT U5400 ( .A(net34475), .Y(n4311) );
  NBUFFX2_LVT U5401 ( .A(n9276), .Y(n4056) );
  NBUFFX2_LVT U5402 ( .A(n9276), .Y(n4057) );
  NBUFFX2_LVT U5403 ( .A(n9276), .Y(n4055) );
  NBUFFX2_LVT U5404 ( .A(n5296), .Y(n3794) );
  NBUFFX2_LVT U5405 ( .A(n5296), .Y(n3793) );
  AND2X1_LVT U5406 ( .A1(n4498), .A2(n9379), .Y(n5296) );
  NBUFFX2_LVT U5407 ( .A(n9378), .Y(n4059) );
  NBUFFX2_LVT U5408 ( .A(n9414), .Y(n4062) );
  NBUFFX2_LVT U5409 ( .A(n9378), .Y(n4060) );
  NBUFFX2_LVT U5410 ( .A(n9414), .Y(n4063) );
  NBUFFX2_LVT U5411 ( .A(n9378), .Y(n4061) );
  NBUFFX2_LVT U5412 ( .A(n9414), .Y(n4064) );
  NAND2X0_LVT U5413 ( .A1(n5481), .A2(n_T_635[1]), .Y(n5483) );
  OR2X1_LVT U5414 ( .A1(n9330), .A2(n4065), .Y(n9332) );
  NBUFFX2_LVT U5415 ( .A(n6860), .Y(n3853) );
  AND3X2_LVT U5416 ( .A1(n3709), .A2(n6957), .A3(n6940), .Y(n3770) );
  NBUFFX2_LVT U5417 ( .A(n6861), .Y(n3857) );
  NBUFFX2_LVT U5418 ( .A(n6859), .Y(n3847) );
  NBUFFX2_LVT U5419 ( .A(n6861), .Y(n3854) );
  NBUFFX2_LVT U5420 ( .A(n6859), .Y(n3846) );
  NBUFFX2_LVT U5421 ( .A(n6861), .Y(n3856) );
  NBUFFX2_LVT U5422 ( .A(n6860), .Y(n3852) );
  NBUFFX2_LVT U5423 ( .A(n6861), .Y(n3855) );
  AND2X1_LVT U5424 ( .A1(n5411), .A2(n5415), .Y(n6858) );
  AND2X1_LVT U5425 ( .A1(n5412), .A2(n5413), .Y(n5411) );
  OR3X1_LVT U5426 ( .A1(wb_ctrl_csr[1]), .A2(wb_ctrl_csr[0]), .A3(
        wb_ctrl_csr[2]), .Y(n5412) );
  AO21X1_LVT U5427 ( .A1(n9249), .A2(n4515), .A3(n9240), .Y(csr_io_exception)
         );
  AO21X1_LVT U5428 ( .A1(n4514), .A2(n9249), .A3(n3262), .Y(n9240) );
  NBUFFX2_LVT U5429 ( .A(n9525), .Y(n3593) );
  NBUFFX2_LVT U5430 ( .A(clock), .Y(n4499) );
  AND2X1_LVT U5431 ( .A1(n5416), .A2(n5415), .Y(n6859) );
  NBUFFX2_LVT U5432 ( .A(n9526), .Y(n3590) );
  NBUFFX2_LVT U5433 ( .A(n9526), .Y(io_fpu_inst[5]) );
  NOR4X1_LVT U5434 ( .A1(n_T_904[6]), .A2(n_T_904[4]), .A3(n_T_904[7]), .A4(
        n3104), .Y(n9513) );
  NBUFFX2_LVT U5435 ( .A(net34660), .Y(n4073) );
  NBUFFX2_LVT U5436 ( .A(net34660), .Y(n4071) );
  NBUFFX2_LVT U5437 ( .A(net34660), .Y(n4072) );
  NBUFFX2_LVT U5438 ( .A(net34480), .Y(n4294) );
  NBUFFX2_LVT U5439 ( .A(net34480), .Y(n4296) );
  NBUFFX2_LVT U5440 ( .A(net34480), .Y(n4292) );
  NBUFFX2_LVT U5441 ( .A(net34480), .Y(n4293) );
  NBUFFX2_LVT U5442 ( .A(net34480), .Y(n4297) );
  NBUFFX2_LVT U5443 ( .A(net34480), .Y(n4295) );
  NBUFFX2_LVT U5444 ( .A(net34480), .Y(n4299) );
  NBUFFX2_LVT U5445 ( .A(net34469), .Y(n4315) );
  NBUFFX2_LVT U5446 ( .A(net34510), .Y(n4254) );
  NBUFFX2_LVT U5447 ( .A(net34500), .Y(n4266) );
  NBUFFX2_LVT U5448 ( .A(net34515), .Y(n4248) );
  NBUFFX2_LVT U5449 ( .A(net34495), .Y(n4272) );
  NBUFFX2_LVT U5450 ( .A(net34505), .Y(n4260) );
  NBUFFX2_LVT U5451 ( .A(net34490), .Y(n4278) );
  NBUFFX2_LVT U5452 ( .A(net34485), .Y(n4284) );
  NBUFFX2_LVT U5453 ( .A(net34665), .Y(n4070) );
  NBUFFX2_LVT U5454 ( .A(net34665), .Y(n4069) );
  NBUFFX2_LVT U5455 ( .A(net34665), .Y(n4068) );
  NBUFFX2_LVT U5456 ( .A(net34645), .Y(n4091) );
  NBUFFX2_LVT U5457 ( .A(net34570), .Y(n4182) );
  NBUFFX2_LVT U5458 ( .A(net34525), .Y(n4236) );
  NBUFFX2_LVT U5459 ( .A(net34535), .Y(n4224) );
  NBUFFX2_LVT U5460 ( .A(net34635), .Y(n4104) );
  NBUFFX2_LVT U5461 ( .A(net34555), .Y(n4200) );
  NBUFFX2_LVT U5462 ( .A(net34575), .Y(n4176) );
  NBUFFX2_LVT U5463 ( .A(net34565), .Y(n4188) );
  NBUFFX2_LVT U5464 ( .A(net34585), .Y(n4164) );
  NBUFFX2_LVT U5465 ( .A(net34605), .Y(n4140) );
  NBUFFX2_LVT U5466 ( .A(net34545), .Y(n4212) );
  NBUFFX2_LVT U5467 ( .A(net34625), .Y(n4116) );
  NBUFFX2_LVT U5468 ( .A(net34615), .Y(n4128) );
  NBUFFX2_LVT U5469 ( .A(net34595), .Y(n4152) );
  NBUFFX2_LVT U5470 ( .A(net34469), .Y(n4313) );
  NBUFFX2_LVT U5471 ( .A(net34469), .Y(n4314) );
  NBUFFX2_LVT U5472 ( .A(net34469), .Y(n4312) );
  NBUFFX2_LVT U5473 ( .A(net34490), .Y(n4273) );
  NBUFFX2_LVT U5474 ( .A(net34510), .Y(n4249) );
  NBUFFX2_LVT U5475 ( .A(net34495), .Y(n4267) );
  NBUFFX2_LVT U5476 ( .A(net34510), .Y(n4253) );
  NBUFFX2_LVT U5477 ( .A(net34510), .Y(n4252) );
  NBUFFX2_LVT U5478 ( .A(net34510), .Y(n4251) );
  NBUFFX2_LVT U5479 ( .A(net34510), .Y(n4250) );
  NBUFFX2_LVT U5480 ( .A(net34500), .Y(n4261) );
  NBUFFX2_LVT U5481 ( .A(net34490), .Y(n4277) );
  NBUFFX2_LVT U5482 ( .A(net34500), .Y(n4263) );
  NBUFFX2_LVT U5483 ( .A(net34485), .Y(n4281) );
  NBUFFX2_LVT U5484 ( .A(net34505), .Y(n4258) );
  NBUFFX2_LVT U5485 ( .A(net34505), .Y(n4257) );
  NBUFFX2_LVT U5486 ( .A(net34505), .Y(n4256) );
  NBUFFX2_LVT U5487 ( .A(net34515), .Y(n4243) );
  NBUFFX2_LVT U5488 ( .A(net34505), .Y(n4255) );
  NBUFFX2_LVT U5489 ( .A(net34515), .Y(n4244) );
  NBUFFX2_LVT U5490 ( .A(net34500), .Y(n4264) );
  NBUFFX2_LVT U5491 ( .A(net34515), .Y(n4245) );
  NBUFFX2_LVT U5492 ( .A(net34505), .Y(n4259) );
  NBUFFX2_LVT U5493 ( .A(net34515), .Y(n4247) );
  NBUFFX2_LVT U5494 ( .A(net34495), .Y(n4271) );
  NBUFFX2_LVT U5495 ( .A(net34485), .Y(n4279) );
  NBUFFX2_LVT U5496 ( .A(net34500), .Y(n4262) );
  NBUFFX2_LVT U5497 ( .A(net34485), .Y(n4282) );
  NBUFFX2_LVT U5498 ( .A(net34485), .Y(n4283) );
  NBUFFX2_LVT U5499 ( .A(net34500), .Y(n4265) );
  NBUFFX2_LVT U5500 ( .A(net34490), .Y(n4274) );
  NBUFFX2_LVT U5501 ( .A(net34490), .Y(n4276) );
  NBUFFX2_LVT U5502 ( .A(net34495), .Y(n4268) );
  NBUFFX2_LVT U5503 ( .A(net34490), .Y(n4275) );
  NBUFFX2_LVT U5504 ( .A(net34515), .Y(n4246) );
  NBUFFX2_LVT U5505 ( .A(net34495), .Y(n4270) );
  NBUFFX2_LVT U5506 ( .A(net34495), .Y(n4269) );
  NBUFFX2_LVT U5507 ( .A(net34485), .Y(n4280) );
  NBUFFX2_LVT U5508 ( .A(n4285), .Y(n4288) );
  NBUFFX2_LVT U5509 ( .A(n4285), .Y(n4289) );
  NBUFFX2_LVT U5510 ( .A(n4285), .Y(n4290) );
  NBUFFX2_LVT U5511 ( .A(n4285), .Y(n4287) );
  NBUFFX2_LVT U5512 ( .A(n4285), .Y(n4291) );
  NBUFFX2_LVT U5513 ( .A(n4285), .Y(n4298) );
  NBUFFX2_LVT U5514 ( .A(n4285), .Y(n4286) );
  NBUFFX2_LVT U5515 ( .A(net34655), .Y(n4079) );
  NBUFFX2_LVT U5516 ( .A(net34630), .Y(n4110) );
  NBUFFX2_LVT U5517 ( .A(net34590), .Y(n4158) );
  NBUFFX2_LVT U5518 ( .A(net34530), .Y(n4230) );
  NBUFFX2_LVT U5519 ( .A(net34560), .Y(n4194) );
  NBUFFX2_LVT U5520 ( .A(net34600), .Y(n4146) );
  NBUFFX2_LVT U5521 ( .A(net34610), .Y(n4134) );
  NBUFFX2_LVT U5522 ( .A(net34520), .Y(n4242) );
  NBUFFX2_LVT U5523 ( .A(net34540), .Y(n4218) );
  NBUFFX2_LVT U5524 ( .A(net34620), .Y(n4122) );
  NBUFFX2_LVT U5525 ( .A(net34550), .Y(n4206) );
  NBUFFX2_LVT U5526 ( .A(net34580), .Y(n4170) );
  XOR2X1_LVT U5527 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(n592), .Y(n5038) );
  XOR2X1_LVT U5528 ( .A1(ibuf_io_inst_0_bits_inst_rs3_4_), .A2(n588), .Y(n5039) );
  XOR2X1_LVT U5529 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(n591), .Y(n5040) );
  XOR2X1_LVT U5530 ( .A1(n1859), .A2(io_dmem_req_bits_tag[4]), .Y(n5042) );
  XOR2X1_LVT U5531 ( .A1(ibuf_io_inst_0_bits_inst_rs3_2_), .A2(
        io_dmem_req_bits_tag[3]), .Y(n5043) );
  XOR2X1_LVT U5532 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n3102), .Y(
        n5025) );
  XOR2X1_LVT U5533 ( .A1(n3781), .A2(n3199), .Y(n5026) );
  XOR2X1_LVT U5534 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n3198), .Y(
        n5022) );
  XOR2X1_LVT U5535 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n3103), .Y(
        n5023) );
  XOR2X1_LVT U5536 ( .A1(n2072), .A2(n3201), .Y(n5024) );
  XOR2X1_LVT U5537 ( .A1(n2876), .A2(n5423), .Y(n5000) );
  XOR2X1_LVT U5538 ( .A1(n2825), .A2(n5426), .Y(n5001) );
  XOR2X1_LVT U5539 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n5428), .Y(
        n5002) );
  XOR2X1_LVT U5540 ( .A1(n2098), .A2(n5306), .Y(n5004) );
  XOR2X1_LVT U5541 ( .A1(n2038), .A2(n5313), .Y(n5005) );
  XOR2X1_LVT U5542 ( .A1(n2876), .A2(n3103), .Y(n4937) );
  XOR2X1_LVT U5543 ( .A1(n2825), .A2(n3199), .Y(n4938) );
  XOR2X1_LVT U5544 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n3198), .Y(
        n4939) );
  XOR2X1_LVT U5545 ( .A1(n2038), .A2(n3043), .Y(n4941) );
  XOR2X1_LVT U5546 ( .A1(n2098), .A2(n3041), .Y(n4942) );
  XOR2X1_LVT U5547 ( .A1(ibuf_io_inst_0_bits_inst_rs3_2_), .A2(n3102), .Y(
        n4920) );
  XOR2X1_LVT U5548 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(n3201), .Y(n4921)
         );
  XOR2X1_LVT U5549 ( .A1(ibuf_io_inst_0_bits_inst_rs3_4_), .A2(n3198), .Y(
        n4922) );
  XOR2X1_LVT U5550 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(wb_waddr[1]), .Y(
        n4924) );
  XOR2X1_LVT U5551 ( .A1(n1859), .A2(wb_waddr[3]), .Y(n4925) );
  XOR2X1_LVT U5552 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n5423), .Y(
        n4871) );
  XOR2X1_LVT U5553 ( .A1(n3781), .A2(n5426), .Y(n4872) );
  XOR2X1_LVT U5554 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n5428), .Y(
        n4868) );
  XOR2X1_LVT U5555 ( .A1(n2072), .A2(n5427), .Y(n4869) );
  XOR2X1_LVT U5556 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n2575), .Y(
        n4870) );
  XOR2X1_LVT U5557 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n5426), .Y(n4688) );
  XOR2X1_LVT U5558 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n5428), .Y(n4689) );
  XOR2X1_LVT U5559 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n5427), .Y(n4690) );
  XOR2X1_LVT U5560 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n2575), .Y(n4686) );
  XOR2X1_LVT U5561 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n5423), .Y(n4687) );
  XOR2X1_LVT U5562 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(n3202), .Y(n4623)
         );
  XOR2X1_LVT U5563 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(n598), .Y(n4625) );
  XOR2X1_LVT U5564 ( .A1(n1859), .A2(n2566), .Y(n4627) );
  XOR2X1_LVT U5565 ( .A1(ibuf_io_inst_0_bits_inst_rs3_4_), .A2(n_T_849[4]), 
        .Y(n4628) );
  XOR2X1_LVT U5566 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n598), .Y(n4622)
         );
  XOR2X1_LVT U5567 ( .A1(n9377), .A2(n_T_698[39]), .Y(n4606) );
  XOR2X1_LVT U5568 ( .A1(n9355), .A2(n124), .Y(n4602) );
  XOR2X1_LVT U5569 ( .A1(n9374), .A2(n104), .Y(n4605) );
  XOR2X1_LVT U5570 ( .A1(n9373), .A2(n_T_698[34]), .Y(n4609) );
  XOR2X1_LVT U5571 ( .A1(n9368), .A2(n_T_698[28]), .Y(n4597) );
  XOR2X1_LVT U5572 ( .A1(n9364), .A2(n_T_698[24]), .Y(n4598) );
  NOR4X1_LVT U5573 ( .A1(n_T_918[39]), .A2(n_T_918[40]), .A3(n_T_918[47]), 
        .A4(n_T_918[60]), .Y(n9464) );
  NOR4X1_LVT U5574 ( .A1(n_T_918[59]), .A2(n_T_918[48]), .A3(n_T_918[62]), 
        .A4(n_T_918[56]), .Y(n9465) );
  NOR4X1_LVT U5575 ( .A1(n_T_918[63]), .A2(n_T_918[46]), .A3(n_T_918[42]), 
        .A4(n_T_918[52]), .Y(n9460) );
  NOR4X1_LVT U5576 ( .A1(n_T_918[41]), .A2(n_T_918[53]), .A3(n_T_918[54]), 
        .A4(n_T_918[50]), .Y(n9461) );
  NOR4X1_LVT U5577 ( .A1(n_T_918[49]), .A2(n_T_918[45]), .A3(n_T_918[61]), 
        .A4(n_T_918[57]), .Y(n9462) );
  NOR4X1_LVT U5578 ( .A1(n_T_918[55]), .A2(n_T_918[58]), .A3(n_T_918[44]), 
        .A4(n_T_918[43]), .Y(n9463) );
  NOR4X1_LVT U5579 ( .A1(n9457), .A2(n9456), .A3(n9455), .A4(n9454), .Y(n9458)
         );
  NBUFFX2_LVT U5580 ( .A(n6830), .Y(n3835) );
  NBUFFX2_LVT U5581 ( .A(n6884), .Y(n3903) );
  NBUFFX2_LVT U5582 ( .A(n6897), .Y(n3956) );
  NBUFFX2_LVT U5583 ( .A(n6895), .Y(n3946) );
  NBUFFX2_LVT U5584 ( .A(n6893), .Y(n3936) );
  NBUFFX2_LVT U5585 ( .A(n6891), .Y(n3926) );
  NBUFFX2_LVT U5586 ( .A(n6812), .Y(n3821) );
  NBUFFX2_LVT U5587 ( .A(n6883), .Y(n3902) );
  NBUFFX2_LVT U5588 ( .A(n6897), .Y(n3955) );
  NBUFFX2_LVT U5589 ( .A(n6895), .Y(n3945) );
  NBUFFX2_LVT U5590 ( .A(n6893), .Y(n3935) );
  NBUFFX2_LVT U5591 ( .A(n6891), .Y(n3925) );
  NBUFFX2_LVT U5592 ( .A(n6882), .Y(n3895) );
  NBUFFX2_LVT U5593 ( .A(n6773), .Y(n3806) );
  NBUFFX2_LVT U5594 ( .A(n6880), .Y(n3893) );
  NBUFFX2_LVT U5595 ( .A(n6795), .Y(n3814) );
  NBUFFX2_LVT U5596 ( .A(n6883), .Y(n3901) );
  NBUFFX2_LVT U5597 ( .A(n6870), .Y(n3873) );
  NBUFFX2_LVT U5598 ( .A(n6829), .Y(n3833) );
  NBUFFX2_LVT U5599 ( .A(n6884), .Y(n3904) );
  NBUFFX2_LVT U5600 ( .A(n6869), .Y(n3870) );
  NBUFFX2_LVT U5601 ( .A(n6812), .Y(n3820) );
  NBUFFX2_LVT U5602 ( .A(n6880), .Y(n3894) );
  NBUFFX2_LVT U5603 ( .A(n6837), .Y(n3838) );
  NBUFFX2_LVT U5604 ( .A(n6811), .Y(n3819) );
  NBUFFX2_LVT U5605 ( .A(n6896), .Y(n3951) );
  NBUFFX2_LVT U5606 ( .A(n6894), .Y(n3941) );
  NBUFFX2_LVT U5607 ( .A(n6892), .Y(n3931) );
  NBUFFX2_LVT U5608 ( .A(n6774), .Y(n3810) );
  NBUFFX2_LVT U5609 ( .A(n6813), .Y(n3823) );
  NBUFFX2_LVT U5610 ( .A(n6884), .Y(n3905) );
  NBUFFX2_LVT U5611 ( .A(n6882), .Y(n3896) );
  NBUFFX2_LVT U5612 ( .A(n6893), .Y(n3933) );
  NBUFFX2_LVT U5613 ( .A(n6774), .Y(n3809) );
  NBUFFX2_LVT U5614 ( .A(n6887), .Y(n3912) );
  NBUFFX2_LVT U5615 ( .A(n6795), .Y(n3813) );
  NBUFFX2_LVT U5616 ( .A(n6868), .Y(n3866) );
  NBUFFX2_LVT U5617 ( .A(n6715), .Y(n3795) );
  NBUFFX2_LVT U5618 ( .A(n6869), .Y(n3869) );
  NBUFFX2_LVT U5619 ( .A(n6882), .Y(n3897) );
  NBUFFX2_LVT U5620 ( .A(n6773), .Y(n3807) );
  NBUFFX2_LVT U5621 ( .A(n6883), .Y(n3899) );
  NBUFFX2_LVT U5622 ( .A(n6897), .Y(n3952) );
  NBUFFX2_LVT U5623 ( .A(n6895), .Y(n3942) );
  NBUFFX2_LVT U5624 ( .A(n6891), .Y(n3922) );
  NBUFFX2_LVT U5625 ( .A(n6880), .Y(n3890) );
  NBUFFX2_LVT U5626 ( .A(n6888), .Y(n3913) );
  NBUFFX2_LVT U5627 ( .A(n6887), .Y(n3911) );
  NBUFFX2_LVT U5628 ( .A(n6773), .Y(n3808) );
  OR2X1_LVT U5629 ( .A1(n8803), .A2(n2645), .Y(n8804) );
  NBUFFX2_LVT U5630 ( .A(n_T_427__T_1136_data[57]), .Y(n4478) );
  NBUFFX2_LVT U5631 ( .A(n6715), .Y(n3797) );
  NBUFFX2_LVT U5632 ( .A(n6837), .Y(n3837) );
  NBUFFX2_LVT U5633 ( .A(n6813), .Y(n3822) );
  NBUFFX2_LVT U5634 ( .A(n6890), .Y(n3917) );
  NBUFFX2_LVT U5635 ( .A(n6891), .Y(n3923) );
  NBUFFX2_LVT U5636 ( .A(n6893), .Y(n3932) );
  NBUFFX2_LVT U5637 ( .A(n6880), .Y(n3891) );
  NBUFFX2_LVT U5638 ( .A(n6879), .Y(n3885) );
  NBUFFX2_LVT U5639 ( .A(n6829), .Y(n3831) );
  NBUFFX2_LVT U5640 ( .A(n6896), .Y(n3947) );
  NBUFFX2_LVT U5641 ( .A(n6897), .Y(n3953) );
  NBUFFX2_LVT U5642 ( .A(n6883), .Y(n3898) );
  NBUFFX2_LVT U5643 ( .A(n6895), .Y(n3943) );
  NBUFFX2_LVT U5644 ( .A(n6894), .Y(n3937) );
  NBUFFX2_LVT U5645 ( .A(n_T_427__T_1136_data[51]), .Y(n4460) );
  NBUFFX2_LVT U5646 ( .A(n_T_427__T_1136_data[53]), .Y(n4466) );
  NBUFFX2_LVT U5647 ( .A(n_T_427__T_1136_data[54]), .Y(n4469) );
  NBUFFX2_LVT U5648 ( .A(n_T_427__T_1136_data[60]), .Y(n4487) );
  OR2X1_LVT U5649 ( .A1(n8878), .A2(n2155), .Y(n8879) );
  NBUFFX2_LVT U5650 ( .A(n_T_427__T_1136_data[59]), .Y(n4484) );
  NBUFFX2_LVT U5651 ( .A(n_T_427__T_1136_data[45]), .Y(n4442) );
  NBUFFX2_LVT U5652 ( .A(n_T_427__T_1136_data[16]), .Y(n4364) );
  NBUFFX2_LVT U5653 ( .A(n_T_427__T_1136_data[24]), .Y(n4386) );
  NAND3X0_LVT U5654 ( .A1(n3731), .A2(n3732), .A3(n3733), .Y(N738) );
  NBUFFX2_LVT U5655 ( .A(n_T_427__T_1136_data[58]), .Y(n4481) );
  NBUFFX2_LVT U5656 ( .A(n_T_427__T_1136_data[47]), .Y(n4448) );
  OA21X1_LVT U5657 ( .A1(n3477), .A2(n3753), .A3(n8442), .Y(n8445) );
  NBUFFX2_LVT U5658 ( .A(n_T_427__T_1136_data[49]), .Y(n4454) );
  NBUFFX2_LVT U5659 ( .A(n6829), .Y(n3832) );
  NBUFFX2_LVT U5660 ( .A(n6883), .Y(n3900) );
  NBUFFX2_LVT U5661 ( .A(n6896), .Y(n3949) );
  AND2X1_LVT U5662 ( .A1(n5457), .A2(n5455), .Y(n6896) );
  NBUFFX2_LVT U5663 ( .A(n6897), .Y(n3954) );
  NBUFFX2_LVT U5664 ( .A(n6894), .Y(n3939) );
  AND2X1_LVT U5665 ( .A1(n5457), .A2(n2034), .Y(n6894) );
  NBUFFX2_LVT U5666 ( .A(n6895), .Y(n3944) );
  NBUFFX2_LVT U5667 ( .A(n6892), .Y(n3929) );
  AND2X1_LVT U5668 ( .A1(n5457), .A2(n5451), .Y(n6892) );
  NBUFFX2_LVT U5669 ( .A(n6893), .Y(n3934) );
  NBUFFX2_LVT U5670 ( .A(n6890), .Y(n3919) );
  AND2X1_LVT U5671 ( .A1(n5457), .A2(n5449), .Y(n6890) );
  NBUFFX2_LVT U5672 ( .A(n6891), .Y(n3924) );
  NBUFFX2_LVT U5673 ( .A(n6879), .Y(n3886) );
  AND2X1_LVT U5674 ( .A1(n5446), .A2(n5454), .Y(n6879) );
  NBUFFX2_LVT U5675 ( .A(n6880), .Y(n3892) );
  AND2X1_LVT U5676 ( .A1(n5437), .A2(n5449), .Y(n3579) );
  NBUFFX2_LVT U5677 ( .A(n6870), .Y(n3872) );
  NBUFFX2_LVT U5678 ( .A(n6865), .Y(n3860) );
  NBUFFX2_LVT U5679 ( .A(n6889), .Y(n3915) );
  NBUFFX2_LVT U5680 ( .A(n6811), .Y(n3818) );
  NBUFFX2_LVT U5681 ( .A(n6887), .Y(n3910) );
  NBUFFX2_LVT U5682 ( .A(n6830), .Y(n3834) );
  XOR2X1_LVT U5683 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n592), .Y(n4861) );
  XOR2X1_LVT U5684 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n588), .Y(n4862) );
  XOR2X1_LVT U5685 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n590), .Y(n4863) );
  XOR2X1_LVT U5686 ( .A1(n3781), .A2(n589), .Y(n4864) );
  XOR2X1_LVT U5687 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n591), .Y(n5044) );
  XOR2X1_LVT U5688 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n3200), .Y(
        n4629) );
  XOR2X1_LVT U5689 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n598), .Y(n4630) );
  XOR2X1_LVT U5690 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n595), .Y(n4631) );
  XOR2X1_LVT U5691 ( .A1(n3781), .A2(n596), .Y(n4632) );
  XOR2X1_LVT U5692 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n_T_849[11]), 
        .Y(n4860) );
  NBUFFX2_LVT U5693 ( .A(n_T_427__T_1136_data[55]), .Y(n4472) );
  NBUFFX2_LVT U5694 ( .A(n_T_427__T_1136_data[32]), .Y(n4406) );
  NBUFFX2_LVT U5695 ( .A(n_T_427__T_1136_data[50]), .Y(n4457) );
  NBUFFX2_LVT U5696 ( .A(n_T_427__T_1136_data[40]), .Y(n4427) );
  NBUFFX2_LVT U5697 ( .A(n_T_427__T_1136_data[1]), .Y(n4321) );
  NBUFFX2_LVT U5698 ( .A(n_T_427__T_1136_data[43]), .Y(n4436) );
  NAND3X0_LVT U5699 ( .A1(n3735), .A2(n3736), .A3(n3737), .Y(N732) );
  OR2X1_LVT U5700 ( .A1(n8624), .A2(n3656), .Y(n8625) );
  NBUFFX2_LVT U5701 ( .A(n_T_427__T_1136_data[52]), .Y(n4463) );
  NAND3X0_LVT U5702 ( .A1(n3748), .A2(n3749), .A3(n3750), .Y(N743) );
  OR2X1_LVT U5703 ( .A1(n9048), .A2(n3632), .Y(n9049) );
  NBUFFX2_LVT U5704 ( .A(n_T_427__T_1136_data[63]), .Y(n4496) );
  NBUFFX2_LVT U5705 ( .A(n_T_427__T_1136_data[19]), .Y(n4373) );
  NBUFFX2_LVT U5706 ( .A(n_T_427__T_1136_data[56]), .Y(n4475) );
  NBUFFX2_LVT U5707 ( .A(n_T_427__T_1136_data[44]), .Y(n4439) );
  NBUFFX2_LVT U5708 ( .A(n_T_427__T_1136_data[37]), .Y(n4419) );
  NBUFFX2_LVT U5709 ( .A(n_T_427__T_1136_data[48]), .Y(n4451) );
  NBUFFX2_LVT U5710 ( .A(n8932), .Y(n3975) );
  OR2X1_LVT U5711 ( .A1(n8987), .A2(n2155), .Y(n8988) );
  NBUFFX2_LVT U5712 ( .A(n_T_427__T_1136_data[62]), .Y(n4493) );
  NBUFFX2_LVT U5713 ( .A(n_T_427__T_1136_data[41]), .Y(n4430) );
  OA21X1_LVT U5714 ( .A1(n3475), .A2(n3601), .A3(n8246), .Y(n8249) );
  NBUFFX2_LVT U5715 ( .A(n3182), .Y(n4048) );
  NBUFFX2_LVT U5716 ( .A(n_T_427__T_1136_data[39]), .Y(n4424) );
  NBUFFX2_LVT U5717 ( .A(n_T_427__T_1136_data[36]), .Y(n4416) );
  NBUFFX2_LVT U5718 ( .A(n8901), .Y(n3967) );
  NBUFFX2_LVT U5719 ( .A(n_T_427__T_1136_data[46]), .Y(n4445) );
  NBUFFX2_LVT U5720 ( .A(n6858), .Y(n3845) );
  NBUFFX2_LVT U5721 ( .A(n9037), .Y(n4021) );
  NBUFFX2_LVT U5722 ( .A(n9041), .Y(n4044) );
  NBUFFX2_LVT U5723 ( .A(n8982), .Y(n3986) );
  NBUFFX2_LVT U5724 ( .A(n_T_427__T_1136_data[34]), .Y(n4411) );
  AND2X1_LVT U5725 ( .A1(n3712), .A2(n_T_427[993]), .Y(n3763) );
  NBUFFX2_LVT U5726 ( .A(n9029), .Y(n3641) );
  NBUFFX2_LVT U5727 ( .A(n_T_427__T_1136_data[61]), .Y(n4490) );
  NBUFFX2_LVT U5728 ( .A(n9016), .Y(n4001) );
  NBUFFX2_LVT U5729 ( .A(n_T_427__T_1136_data[17]), .Y(n4367) );
  NBUFFX2_LVT U5730 ( .A(n_T_427__T_1136_data[20]), .Y(n4376) );
  NBUFFX2_LVT U5731 ( .A(n9042), .Y(n4052) );
  NBUFFX2_LVT U5732 ( .A(n8931), .Y(n3971) );
  NBUFFX2_LVT U5733 ( .A(n9037), .Y(n4022) );
  NBUFFX2_LVT U5734 ( .A(n9039), .Y(n4035) );
  NBUFFX2_LVT U5735 ( .A(n_T_427__T_1136_data[42]), .Y(n4433) );
  NBUFFX2_LVT U5736 ( .A(n9016), .Y(n4002) );
  INVX1_LVT U5737 ( .A(n9014), .Y(n3995) );
  NBUFFX2_LVT U5738 ( .A(n9039), .Y(n4031) );
  NBUFFX2_LVT U5739 ( .A(n8900), .Y(n3961) );
  NBUFFX2_LVT U5740 ( .A(n8981), .Y(n3980) );
  INVX1_LVT U5741 ( .A(n9006), .Y(n3990) );
  NBUFFX2_LVT U5742 ( .A(n9015), .Y(n4000) );
  NBUFFX2_LVT U5743 ( .A(n_T_427__T_1136_data[0]), .Y(n4318) );
  NBUFFX2_LVT U5744 ( .A(n6858), .Y(n3841) );
  NBUFFX2_LVT U5745 ( .A(n9041), .Y(n4041) );
  NBUFFX2_LVT U5746 ( .A(n3182), .Y(n4045) );
  NBUFFX2_LVT U5747 ( .A(n9039), .Y(n4032) );
  NBUFFX2_LVT U5748 ( .A(n9038), .Y(n4030) );
  NBUFFX2_LVT U5749 ( .A(n9037), .Y(n4018) );
  NBUFFX2_LVT U5750 ( .A(n9042), .Y(n4049) );
  NBUFFX2_LVT U5751 ( .A(n_T_427__T_1136_data[30]), .Y(n4401) );
  NBUFFX2_LVT U5752 ( .A(n8900), .Y(n3963) );
  NBUFFX2_LVT U5753 ( .A(n8981), .Y(n3982) );
  NBUFFX2_LVT U5754 ( .A(n6859), .Y(n3848) );
  NBUFFX2_LVT U5755 ( .A(n_T_427__T_1136_data[27]), .Y(n4393) );
  NBUFFX2_LVT U5756 ( .A(n_T_427__T_1136_data[23]), .Y(n4383) );
  NBUFFX2_LVT U5757 ( .A(n6861), .Y(n3858) );
  NBUFFX2_LVT U5758 ( .A(n6858), .Y(n3844) );
  NBUFFX2_LVT U5759 ( .A(n9041), .Y(n4043) );
  NBUFFX2_LVT U5760 ( .A(n3182), .Y(n4047) );
  NBUFFX2_LVT U5761 ( .A(n8932), .Y(n3974) );
  NBUFFX2_LVT U5762 ( .A(n8901), .Y(n3966) );
  NBUFFX2_LVT U5763 ( .A(n8931), .Y(n3970) );
  NBUFFX2_LVT U5764 ( .A(n8982), .Y(n3985) );
  NBUFFX2_LVT U5765 ( .A(n9039), .Y(n4034) );
  NBUFFX2_LVT U5766 ( .A(n9038), .Y(n4028) );
  NBUFFX2_LVT U5767 ( .A(n9037), .Y(n4020) );
  NBUFFX2_LVT U5768 ( .A(n_T_427__T_1136_data[29]), .Y(n4398) );
  NBUFFX2_LVT U5769 ( .A(n6860), .Y(n3851) );
  NBUFFX2_LVT U5770 ( .A(n9016), .Y(n4003) );
  NBUFFX2_LVT U5771 ( .A(n9015), .Y(n3998) );
  NBUFFX2_LVT U5772 ( .A(n9041), .Y(n4042) );
  NBUFFX2_LVT U5773 ( .A(n8900), .Y(n3962) );
  NBUFFX2_LVT U5774 ( .A(n3182), .Y(n4046) );
  NBUFFX2_LVT U5775 ( .A(n8981), .Y(n3981) );
  NBUFFX2_LVT U5776 ( .A(n8932), .Y(n3973) );
  NBUFFX2_LVT U5777 ( .A(n8901), .Y(n3965) );
  NBUFFX2_LVT U5778 ( .A(n8931), .Y(n3969) );
  NBUFFX2_LVT U5779 ( .A(n8982), .Y(n3984) );
  NBUFFX2_LVT U5780 ( .A(n9039), .Y(n4033) );
  NBUFFX2_LVT U5781 ( .A(n9038), .Y(n4029) );
  NBUFFX2_LVT U5782 ( .A(n8980), .Y(n3977) );
  NBUFFX2_LVT U5783 ( .A(n9037), .Y(n4019) );
  NBUFFX2_LVT U5784 ( .A(n9042), .Y(n4050) );
  NBUFFX2_LVT U5785 ( .A(n_T_427__T_1136_data[18]), .Y(n4370) );
  NBUFFX2_LVT U5786 ( .A(n6859), .Y(n3849) );
  NBUFFX2_LVT U5787 ( .A(n6858), .Y(n3843) );
  INVX1_LVT U5788 ( .A(n9008), .Y(n3993) );
  XOR2X1_LVT U5789 ( .A1(io_fpu_inst[20]), .A2(n9522), .Y(n5142) );
  INVX1_LVT U5790 ( .A(n5394), .Y(n3567) );
  OA21X1_LVT U5791 ( .A1(n5118), .A2(n3039), .A3(n5111), .Y(n5112) );
  XOR2X1_LVT U5792 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n592), .Y(n5011) );
  XOR2X1_LVT U5793 ( .A1(n2876), .A2(n598), .Y(n4615) );
  XOR2X1_LVT U5794 ( .A1(ibuf_io_inst_0_bits_inst_rs1[2]), .A2(n3200), .Y(
        n4616) );
  OA21X1_LVT U5795 ( .A1(io_fpu_inst[2]), .A2(n3076), .A3(n5165), .Y(n5109) );
  NBUFFX2_LVT U5796 ( .A(n6888), .Y(n3914) );
  NBUFFX2_LVT U5797 ( .A(n6885), .Y(n3907) );
  NBUFFX2_LVT U5798 ( .A(n6885), .Y(n3906) );
  NBUFFX2_LVT U5799 ( .A(n6838), .Y(n3839) );
  AND3X1_LVT U5800 ( .A1(n6118), .A2(n6117), .A3(n6116), .Y(n3091) );
  NAND2X0_LVT U5801 ( .A1(wb_cause[3]), .A2(n9252), .Y(n3100) );
  NBUFFX2_LVT U5802 ( .A(n9015), .Y(n3997) );
  NBUFFX2_LVT U5803 ( .A(n9015), .Y(n3996) );
  NBUFFX2_LVT U5804 ( .A(n9015), .Y(n3999) );
  NBUFFX2_LVT U5805 ( .A(n9016), .Y(n4004) );
  NBUFFX2_LVT U5806 ( .A(n9016), .Y(n4005) );
  NBUFFX2_LVT U5807 ( .A(n6886), .Y(n3909) );
  NBUFFX2_LVT U5808 ( .A(n6889), .Y(n3916) );
  AND4X1_LVT U5809 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .Y(n3181)
         );
  NBUFFX2_LVT U5810 ( .A(n6796), .Y(n3816) );
  NBUFFX2_LVT U5811 ( .A(n6796), .Y(n3815) );
  NBUFFX2_LVT U5812 ( .A(n6898), .Y(n3959) );
  NBUFFX2_LVT U5813 ( .A(n6892), .Y(n3927) );
  NBUFFX2_LVT U5814 ( .A(n6892), .Y(n3930) );
  NBUFFX2_LVT U5815 ( .A(n6892), .Y(n3928) );
  NBUFFX2_LVT U5816 ( .A(n6890), .Y(n3920) );
  NBUFFX2_LVT U5817 ( .A(n6890), .Y(n3918) );
  NBUFFX2_LVT U5818 ( .A(n6890), .Y(n3921) );
  NBUFFX2_LVT U5819 ( .A(n6894), .Y(n3938) );
  NBUFFX2_LVT U5820 ( .A(n6894), .Y(n3940) );
  NBUFFX2_LVT U5821 ( .A(n6896), .Y(n3948) );
  NBUFFX2_LVT U5822 ( .A(n6896), .Y(n3950) );
  NBUFFX2_LVT U5823 ( .A(n6879), .Y(n3889) );
  NBUFFX2_LVT U5824 ( .A(n6879), .Y(n3888) );
  NBUFFX2_LVT U5825 ( .A(n6879), .Y(n3887) );
  NBUFFX2_LVT U5826 ( .A(n8980), .Y(n3978) );
  AND3X1_LVT U5827 ( .A1(n6166), .A2(n6165), .A3(n6164), .Y(n3183) );
  NAND2X0_LVT U5828 ( .A1(n6946), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n3184) );
  NBUFFX2_LVT U5829 ( .A(n6810), .Y(n3817) );
  NBUFFX2_LVT U5830 ( .A(n6859), .Y(n3850) );
  NBUFFX2_LVT U5831 ( .A(n6858), .Y(n3842) );
  NBUFFX2_LVT U5832 ( .A(n9101), .Y(n4054) );
  AND4X1_LVT U5833 ( .A1(n9481), .A2(n9480), .A3(n9479), .A4(n9478), .Y(n3204)
         );
  AND2X1_LVT U5834 ( .A1(n3078), .A2(n9105), .Y(n3566) );
  OA22X1_LVT U5835 ( .A1(n5115), .A2(n3571), .A3(n3570), .A4(n1699), .Y(n3576)
         );
  OR2X1_LVT U5836 ( .A1(csr_io_status_isa[3]), .A2(n3039), .Y(n3571) );
  AND4X1_LVT U5837 ( .A1(n3576), .A2(n5112), .A3(n5121), .A4(n5120), .Y(n3572)
         );
  AND2X1_LVT U5838 ( .A1(n3574), .A2(n5113), .Y(n3573) );
  NAND2X0_LVT U5839 ( .A1(n9231), .A2(n3575), .Y(n9413) );
  AO22X1_LVT U5840 ( .A1(n1853), .A2(n3577), .A3(n1867), .A4(n1891), .Y(
        id_ctrl_sel_imm[0]) );
  NAND4X0_LVT U5841 ( .A1(n4616), .A2(n4615), .A3(n4617), .A4(n3581), .Y(n4847) );
  NAND2X0_LVT U5842 ( .A1(n5446), .A2(n5450), .Y(n6878) );
  AND2X1_LVT U5843 ( .A1(n9446), .A2(io_fpu_inst[12]), .Y(n9230) );
  AND2X1_LVT U5844 ( .A1(n9446), .A2(n3077), .Y(n5101) );
  NAND2X0_LVT U5845 ( .A1(n3583), .A2(io_fpu_inst[14]), .Y(n5105) );
  NAND2X0_LVT U5846 ( .A1(n2547), .A2(n2131), .Y(n5122) );
  NAND2X0_LVT U5847 ( .A1(n5077), .A2(n5076), .Y(n3584) );
  AND2X1_LVT U5848 ( .A1(n9440), .A2(io_fpu_inst[28]), .Y(n3585) );
  OA22X1_LVT U5849 ( .A1(n5443), .A2(n3586), .A3(n3490), .A4(n3880), .Y(n5445)
         );
  OA22X1_LVT U5850 ( .A1(n6695), .A2(n3586), .A3(n3491), .A4(n3882), .Y(n6698)
         );
  OA22X1_LVT U5851 ( .A1(n6720), .A2(n3586), .A3(n3492), .A4(n3882), .Y(n6723)
         );
  OA22X1_LVT U5852 ( .A1(n6739), .A2(n3586), .A3(n3493), .A4(n3882), .Y(n6743)
         );
  OA22X1_LVT U5853 ( .A1(n6801), .A2(n3586), .A3(n3483), .A4(n3882), .Y(n6805)
         );
  OA22X1_LVT U5854 ( .A1(n6843), .A2(n3586), .A3(n3484), .A4(n3882), .Y(n6846)
         );
  NBUFFX2_LVT U5855 ( .A(net34650), .Y(n4085) );
  NAND2X0_LVT U5856 ( .A1(n9253), .A2(csr_io_exception), .Y(n9254) );
  AND2X1_LVT U5857 ( .A1(n3100), .A2(n3589), .Y(n9253) );
  INVX1_LVT U5858 ( .A(wb_cause[63]), .Y(n3589) );
  AND3X1_LVT U5918 ( .A1(n7138), .A2(n7137), .A3(n7136), .Y(n3598) );
  AND3X1_LVT U5919 ( .A1(n7131), .A2(n7130), .A3(n7129), .Y(n3599) );
  NBUFFX2_LVT U5920 ( .A(n9053), .Y(n3789) );
  NBUFFX2_LVT U5921 ( .A(n3613), .Y(n3602) );
  NBUFFX2_LVT U5922 ( .A(n9004), .Y(n3603) );
  NBUFFX2_LVT U5923 ( .A(n9004), .Y(n3604) );
  NBUFFX2_LVT U5924 ( .A(n9004), .Y(n3605) );
  NBUFFX2_LVT U5925 ( .A(n3613), .Y(n3606) );
  NBUFFX2_LVT U5926 ( .A(n9004), .Y(n3607) );
  NBUFFX2_LVT U5927 ( .A(n3613), .Y(n3608) );
  NBUFFX2_LVT U5928 ( .A(n3613), .Y(n3609) );
  NBUFFX2_LVT U5929 ( .A(n9004), .Y(n3611) );
  NBUFFX2_LVT U5930 ( .A(n9047), .Y(n3612) );
  NBUFFX2_LVT U5931 ( .A(n9021), .Y(n3615) );
  NBUFFX2_LVT U5932 ( .A(n9021), .Y(n3616) );
  NBUFFX2_LVT U5933 ( .A(n9021), .Y(n3617) );
  NBUFFX2_LVT U5934 ( .A(n9021), .Y(n3618) );
  NBUFFX2_LVT U5935 ( .A(n9021), .Y(n3619) );
  NBUFFX2_LVT U5936 ( .A(n9021), .Y(n3620) );
  NBUFFX2_LVT U5937 ( .A(n9021), .Y(n3621) );
  AND3X1_LVT U5938 ( .A1(n8006), .A2(n8007), .A3(n8008), .Y(n3622) );
  AND3X1_LVT U5939 ( .A1(n8005), .A2(n8004), .A3(n8003), .Y(n3623) );
  NBUFFX2_LVT U5940 ( .A(n9058), .Y(n3624) );
  NBUFFX2_LVT U5941 ( .A(n9007), .Y(n3626) );
  NBUFFX2_LVT U5942 ( .A(n9007), .Y(n3627) );
  NBUFFX2_LVT U5943 ( .A(n9007), .Y(n3628) );
  NBUFFX2_LVT U5944 ( .A(n9007), .Y(n3629) );
  NBUFFX2_LVT U5945 ( .A(n9007), .Y(n3630) );
  AND3X1_LVT U5946 ( .A1(n8942), .A2(n8941), .A3(n8940), .Y(n3634) );
  NBUFFX2_LVT U5947 ( .A(n9029), .Y(n3635) );
  NBUFFX2_LVT U5948 ( .A(n9029), .Y(n3636) );
  NBUFFX2_LVT U5949 ( .A(n9029), .Y(n3638) );
  NBUFFX2_LVT U5950 ( .A(n9029), .Y(n3639) );
  NBUFFX2_LVT U5951 ( .A(n9029), .Y(n3640) );
  OR2X1_LVT U5952 ( .A1(n4016), .A2(n3644), .Y(n8753) );
  OR2X1_LVT U5953 ( .A1(n2090), .A2(n3645), .Y(n7874) );
  OR2X1_LVT U5954 ( .A1(n9412), .A2(n3646), .Y(n6971) );
  NBUFFX2_LVT U5955 ( .A(n8944), .Y(n3647) );
  NBUFFX2_LVT U5956 ( .A(n9022), .Y(n3648) );
  NBUFFX2_LVT U5957 ( .A(n9022), .Y(n3650) );
  NBUFFX2_LVT U5958 ( .A(n9022), .Y(n3651) );
  NBUFFX2_LVT U5959 ( .A(n9022), .Y(n3652) );
  OR2X1_LVT U5960 ( .A1(n2069), .A2(n3655), .Y(n7966) );
  NBUFFX2_LVT U5961 ( .A(n9012), .Y(n3657) );
  OR2X1_LVT U5962 ( .A1(n2089), .A2(n3659), .Y(n8389) );
  OR2X1_LVT U5963 ( .A1(n2090), .A2(n3660), .Y(n8426) );
  OR2X1_LVT U5964 ( .A1(n4016), .A2(n3090), .Y(n7814) );
  AND3X1_LVT U5965 ( .A1(n8725), .A2(n8724), .A3(n8723), .Y(n3662) );
  NBUFFX2_LVT U5966 ( .A(n9030), .Y(n3668) );
  NBUFFX2_LVT U5967 ( .A(n9030), .Y(n3669) );
  NBUFFX2_LVT U5968 ( .A(n3666), .Y(n3670) );
  NBUFFX2_LVT U5969 ( .A(n3666), .Y(n3671) );
  NBUFFX2_LVT U5970 ( .A(n3666), .Y(n3672) );
  NBUFFX2_LVT U5971 ( .A(n9030), .Y(n3673) );
  NBUFFX2_LVT U5972 ( .A(n9030), .Y(n3674) );
  NBUFFX2_LVT U5973 ( .A(n9030), .Y(n3675) );
  AND3X1_LVT U5974 ( .A1(n8037), .A2(n8036), .A3(n8038), .Y(n3676) );
  AND3X1_LVT U5975 ( .A1(n8041), .A2(n8040), .A3(n8039), .Y(n3677) );
  AND3X1_LVT U5976 ( .A1(n8736), .A2(n8735), .A3(n8737), .Y(n3678) );
  OR2X1_LVT U5977 ( .A1(n4016), .A2(n3679), .Y(n6943) );
  AND3X1_LVT U5978 ( .A1(n7532), .A2(n7531), .A3(n7530), .Y(n3680) );
  AND3X1_LVT U5979 ( .A1(n7515), .A2(n7514), .A3(n7513), .Y(n3681) );
  AND3X1_LVT U5980 ( .A1(n7517), .A2(n7518), .A3(n7519), .Y(n3682) );
  OR2X1_LVT U5981 ( .A1(n2069), .A2(n3685), .Y(n8131) );
  OA21X1_LVT U5982 ( .A1(n3412), .A2(n3753), .A3(n8591), .Y(n8594) );
  OA21X1_LVT U5983 ( .A1(n3413), .A2(n3751), .A3(n8374), .Y(n8377) );
  OR2X1_LVT U5984 ( .A1(n2090), .A2(n3686), .Y(n6997) );
  OR2X1_LVT U5985 ( .A1(n2089), .A2(n3687), .Y(n8072) );
  OR2X1_LVT U5986 ( .A1(n2090), .A2(n3688), .Y(n8321) );
  OA21X1_LVT U5987 ( .A1(n3414), .A2(n3753), .A3(n8488), .Y(n8491) );
  OA21X1_LVT U5988 ( .A1(n3415), .A2(n3753), .A3(n8358), .Y(n8361) );
  AND3X1_LVT U5989 ( .A1(n8024), .A2(n8025), .A3(n8026), .Y(n3690) );
  NBUFFX2_LVT U5990 ( .A(n3708), .Y(n3691) );
  AND3X1_LVT U5991 ( .A1(n7705), .A2(n7704), .A3(n7703), .Y(n3693) );
  AND3X1_LVT U5992 ( .A1(n7701), .A2(n7700), .A3(n7699), .Y(n3694) );
  AND3X1_LVT U5993 ( .A1(n7718), .A2(n7717), .A3(n7716), .Y(n3695) );
  AND3X1_LVT U5994 ( .A1(n7454), .A2(n7453), .A3(n7452), .Y(n3696) );
  AND3X1_LVT U5995 ( .A1(n7470), .A2(n7469), .A3(n7468), .Y(n3697) );
  AND3X1_LVT U5996 ( .A1(n7738), .A2(n7737), .A3(n7736), .Y(n3698) );
  AND3X1_LVT U5997 ( .A1(n7734), .A2(n7733), .A3(n7732), .Y(n3699) );
  AND3X1_LVT U5998 ( .A1(n7751), .A2(n7750), .A3(n7749), .Y(n3700) );
  AND3X1_LVT U5999 ( .A1(n7607), .A2(n7606), .A3(n7605), .Y(n3701) );
  AND3X1_LVT U6000 ( .A1(n7622), .A2(n7621), .A3(n7620), .Y(n3702) );
  AND3X1_LVT U6001 ( .A1(n7544), .A2(n7543), .A3(n7542), .Y(n3703) );
  AND3X1_LVT U6002 ( .A1(n7559), .A2(n7558), .A3(n7557), .Y(n3704) );
  AND3X1_LVT U6003 ( .A1(n7575), .A2(n7574), .A3(n7573), .Y(n3705) );
  AND3X1_LVT U6004 ( .A1(n7591), .A2(n7590), .A3(n7589), .Y(n3706) );
  NBUFFX2_LVT U6005 ( .A(n8994), .Y(n3707) );
  NAND2X0_LVT U6006 ( .A1(n3182), .A2(n8105), .Y(n3708) );
  OR2X1_LVT U6007 ( .A1(n4016), .A2(n3710), .Y(n7441) );
  OR2X1_LVT U6008 ( .A1(n4016), .A2(n3711), .Y(n7847) );
  NBUFFX2_LVT U6009 ( .A(n9059), .Y(n3713) );
  NBUFFX2_LVT U6010 ( .A(n9059), .Y(n3714) );
  NBUFFX2_LVT U6011 ( .A(n9059), .Y(n3791) );
  AND3X1_LVT U6012 ( .A1(n8696), .A2(n8695), .A3(n8694), .Y(n3718) );
  AND3X1_LVT U6013 ( .A1(n8692), .A2(n8691), .A3(n8690), .Y(n3720) );
  AND3X1_LVT U6014 ( .A1(n8660), .A2(n8659), .A3(n8658), .Y(n3721) );
  AND3X1_LVT U6015 ( .A1(n8654), .A2(n8653), .A3(n8652), .Y(n3722) );
  AND2X1_LVT U6016 ( .A1(n8910), .A2(n8909), .Y(n3723) );
  AND3X1_LVT U6017 ( .A1(n8908), .A2(n8907), .A3(n8906), .Y(n3724) );
  AND2X1_LVT U6018 ( .A1(n8588), .A2(n8587), .Y(n3726) );
  AND3X1_LVT U6019 ( .A1(n8586), .A2(n8585), .A3(n8584), .Y(n3727) );
  NAND3X0_LVT U6020 ( .A1(n3728), .A2(n3729), .A3(n3730), .Y(N739) );
  NOR3X0_LVT U6021 ( .A1(n8849), .A2(n8850), .A3(n8851), .Y(n3733) );
  NOR3X0_LVT U6022 ( .A1(n8813), .A2(n8814), .A3(n8815), .Y(n3734) );
  NAND3X0_LVT U6023 ( .A1(n3738), .A2(n3739), .A3(n3740), .Y(N729) );
  NAND3X0_LVT U6024 ( .A1(n3741), .A2(n3742), .A3(n3743), .Y(N727) );
  NBUFFX2_LVT U6025 ( .A(n9058), .Y(n3745) );
  XOR2X1_LVT U6026 ( .A1(n2876), .A2(n9390), .Y(n6907) );
  NBUFFX2_LVT U6027 ( .A(n9014), .Y(n3751) );
  NBUFFX2_LVT U6028 ( .A(n9028), .Y(n3752) );
  NBUFFX2_LVT U6029 ( .A(n9014), .Y(n3753) );
  AND3X1_LVT U6030 ( .A1(n8241), .A2(n8240), .A3(n8239), .Y(n3754) );
  NBUFFX2_LVT U6031 ( .A(n9026), .Y(n3755) );
  AND3X1_LVT U6032 ( .A1(n7993), .A2(n7992), .A3(n7991), .Y(n3762) );
  AOI21X1_LVT U6033 ( .A1(n3716), .A2(n_T_427[1057]), .A3(n3763), .Y(n8008) );
  INVX1_LVT U6034 ( .A(n9006), .Y(n3764) );
  AND2X1_LVT U6035 ( .A1(n6962), .A2(n6965), .Y(n3765) );
  AND3X1_LVT U6036 ( .A1(n7989), .A2(n7988), .A3(n7987), .Y(n3766) );
  NBUFFX2_LVT U6037 ( .A(n9006), .Y(n3767) );
  OR2X1_LVT U6038 ( .A1(n3653), .A2(n3774), .Y(n8492) );
  AOI21X1_LVT U6039 ( .A1(n4014), .A2(n_T_427[1058]), .A3(n3775), .Y(n8041) );
  AND2X1_LVT U6040 ( .A1(n3712), .A2(n_T_427[994]), .Y(n3775) );
  AND2X1_LVT U6041 ( .A1(n3712), .A2(n_T_427[1014]), .Y(n3776) );
  AND2X1_LVT U6042 ( .A1(n3712), .A2(n_T_427[1000]), .Y(n3777) );
  AND3X1_LVT U6043 ( .A1(n8237), .A2(n8236), .A3(n8235), .Y(n3778) );
  AND3X1_LVT U6044 ( .A1(n8022), .A2(n8021), .A3(n8020), .Y(n3779) );
  AND3X1_LVT U6045 ( .A1(n8720), .A2(n8719), .A3(n8718), .Y(n3780) );
  NBUFFX2_LVT U6046 ( .A(n9035), .Y(n3786) );
  NBUFFX2_LVT U6047 ( .A(n9035), .Y(n3787) );
  NBUFFX2_LVT U6048 ( .A(n9035), .Y(n3788) );
  NBUFFX2_LVT U6049 ( .A(n9053), .Y(n3790) );
  NBUFFX2_LVT U6050 ( .A(net34475), .Y(n4300) );
  NBUFFX2_LVT U6051 ( .A(net34475), .Y(n4301) );
  NBUFFX2_LVT U6052 ( .A(net34475), .Y(n4302) );
  NBUFFX2_LVT U6053 ( .A(net34475), .Y(n4303) );
  NBUFFX2_LVT U6054 ( .A(net34475), .Y(n4304) );
  NBUFFX2_LVT U6055 ( .A(net34475), .Y(n4305) );
  NBUFFX2_LVT U6056 ( .A(net34475), .Y(n4306) );
  NBUFFX2_LVT U6057 ( .A(net34475), .Y(n4307) );
  NBUFFX2_LVT U6058 ( .A(net34475), .Y(n4308) );
  NBUFFX2_LVT U6059 ( .A(net34475), .Y(n4309) );
  NBUFFX2_LVT U6060 ( .A(net34475), .Y(n4310) );
  AND2X1_LVT U6061 ( .A1(n9529), .A2(n3590), .Y(n4507) );
  INVX1_LVT U6062 ( .A(n9520), .Y(n9437) );
  NAND2X0_LVT U6063 ( .A1(n3593), .A2(io_fpu_inst[4]), .Y(n9111) );
  INVX1_LVT U6064 ( .A(io_fpu_inst[10]), .Y(n9447) );
  AO21X1_LVT U6065 ( .A1(n9446), .A2(n9105), .A3(n9445), .Y(n4505) );
  NAND2X0_LVT U6066 ( .A1(n9529), .A2(n9446), .Y(n5086) );
  AND2X1_LVT U6067 ( .A1(n2137), .A2(n4507), .Y(n4510) );
  NAND2X0_LVT U6068 ( .A1(n9435), .A2(n9524), .Y(n4508) );
  NAND2X0_LVT U6069 ( .A1(n9438), .A2(n5394), .Y(n5149) );
  AND2X1_LVT U6070 ( .A1(wb_ctrl_mem), .A2(wb_reg_valid), .Y(n9249) );
  OR2X1_LVT U6071 ( .A1(io_dmem_s2_xcpt_pf_st), .A2(io_dmem_s2_xcpt_pf_ld), 
        .Y(n9239) );
  OR3X1_LVT U6072 ( .A1(io_dmem_s2_xcpt_ae_ld), .A2(io_dmem_s2_xcpt_ae_st), 
        .A3(n9239), .Y(n4515) );
  OR2X1_LVT U6073 ( .A1(io_dmem_s2_xcpt_ma_st), .A2(io_dmem_s2_xcpt_ma_ld), 
        .Y(n4514) );
  INVX1_LVT U6074 ( .A(mem_br_target_38_), .Y(n4516) );
  INVX1_LVT U6075 ( .A(mem_br_target_26_), .Y(n4517) );
  MUX21X1_LVT U6076 ( .A1(n_T_918[16]), .A2(mem_br_target_16_), .S0(n4591), 
        .Y(n9356) );
  AND3X1_LVT U6077 ( .A1(n4521), .A2(n4520), .A3(n4519), .Y(n4566) );
  INVX1_LVT U6078 ( .A(mem_br_target_36_), .Y(n4522) );
  INVX1_LVT U6079 ( .A(mem_br_target_27_), .Y(n4523) );
  INVX1_LVT U6080 ( .A(mem_br_target_23_), .Y(n4524) );
  INVX1_LVT U6081 ( .A(mem_br_target_18_), .Y(n4525) );
  INVX1_LVT U6082 ( .A(mem_br_target_14_), .Y(n4526) );
  INVX1_LVT U6083 ( .A(mem_br_target_12_), .Y(n4527) );
  INVX1_LVT U6084 ( .A(mem_br_target_8_), .Y(n4528) );
  MUX21X1_LVT U6085 ( .A1(n3222), .A2(n4528), .S0(n3792), .Y(n9511) );
  INVX1_LVT U6086 ( .A(mem_br_target_7_), .Y(n4529) );
  MUX21X1_LVT U6087 ( .A1(n3214), .A2(n4529), .S0(n4591), .Y(n9499) );
  INVX1_LVT U6088 ( .A(mem_br_target_3_), .Y(n4530) );
  MUX21X1_LVT U6089 ( .A1(n3208), .A2(n4530), .S0(n4591), .Y(n9503) );
  INVX1_LVT U6090 ( .A(ibuf_io_pc[0]), .Y(n4531) );
  OA21X1_LVT U6091 ( .A1(io_imem_resp_valid), .A2(ibuf_io_inst_0_valid), .A3(
        n4531), .Y(n4536) );
  MUX21X1_LVT U6092 ( .A1(n_T_918[2]), .A2(mem_br_target_2_), .S0(n3792), .Y(
        n9334) );
  INVX1_LVT U6093 ( .A(mem_br_target_1_), .Y(n4533) );
  AND4X1_LVT U6094 ( .A1(n4537), .A2(n4536), .A3(n4535), .A4(n4534), .Y(n4542)
         );
  INVX1_LVT U6095 ( .A(mem_br_target_5_), .Y(n4538) );
  MUX21X1_LVT U6096 ( .A1(n3109), .A2(n4538), .S0(n4591), .Y(n9484) );
  INVX1_LVT U6097 ( .A(mem_br_target_4_), .Y(n4539) );
  MUX21X1_LVT U6098 ( .A1(n3112), .A2(n4539), .S0(n3792), .Y(n9495) );
  AND4X1_LVT U6099 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .Y(n4548)
         );
  INVX1_LVT U6100 ( .A(mem_br_target_9_), .Y(n4544) );
  MUX21X1_LVT U6101 ( .A1(n3108), .A2(n4544), .S0(n4591), .Y(n9507) );
  INVX1_LVT U6102 ( .A(mem_br_target_6_), .Y(n4545) );
  MUX21X1_LVT U6103 ( .A1(n3217), .A2(n4545), .S0(n3792), .Y(n9485) );
  AND4X1_LVT U6104 ( .A1(n4549), .A2(n4548), .A3(n4547), .A4(n4546), .Y(n4552)
         );
  INVX1_LVT U6105 ( .A(mem_br_target_17_), .Y(n4550) );
  AND2X1_LVT U6106 ( .A1(n4552), .A2(n4551), .Y(n4553) );
  AND4X1_LVT U6107 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .Y(n4559)
         );
  AND4X1_LVT U6108 ( .A1(n4561), .A2(n4560), .A3(n4559), .A4(n4558), .Y(n4564)
         );
  INVX1_LVT U6109 ( .A(mem_br_target_31_), .Y(n4562) );
  AND4X1_LVT U6110 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .Y(n4596)
         );
  INVX1_LVT U6111 ( .A(mem_br_target_37_), .Y(n4567) );
  MUX21X1_LVT U6112 ( .A1(n_T_918[35]), .A2(mem_br_target_35_), .S0(n4591), 
        .Y(n9374) );
  INVX1_LVT U6113 ( .A(mem_br_target_29_), .Y(n4568) );
  INVX1_LVT U6114 ( .A(mem_br_target_10_), .Y(n4569) );
  INVX1_LVT U6115 ( .A(mem_br_target_13_), .Y(n4570) );
  INVX1_LVT U6116 ( .A(mem_br_target_11_), .Y(n4571) );
  INVX1_LVT U6117 ( .A(mem_br_target_19_), .Y(n4572) );
  MUX21X1_LVT U6118 ( .A1(n_T_918[39]), .A2(n3205), .S0(n9470), .Y(n4573) );
  NOR4X1_LVT U6119 ( .A1(n4577), .A2(n4576), .A3(n4575), .A4(n4574), .Y(n4595)
         );
  INVX1_LVT U6120 ( .A(mem_br_target_20_), .Y(n4578) );
  INVX1_LVT U6121 ( .A(mem_br_target_22_), .Y(n4579) );
  INVX1_LVT U6122 ( .A(mem_br_target_33_), .Y(n4580) );
  INVX1_LVT U6123 ( .A(mem_br_target_25_), .Y(n4581) );
  NAND4X0_LVT U6124 ( .A1(n4585), .A2(n4584), .A3(n4583), .A4(n4582), .Y(n4588) );
  INVX1_LVT U6125 ( .A(mem_br_target_30_), .Y(n4586) );
  NOR4X1_LVT U6126 ( .A1(n4590), .A2(n4589), .A3(n4588), .A4(n4587), .Y(n4594)
         );
  INVX1_LVT U6127 ( .A(mem_br_target_32_), .Y(n4592) );
  NAND4X0_LVT U6128 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .Y(n4614) );
  NOR3X0_LVT U6129 ( .A1(n4598), .A2(n4597), .A3(n9482), .Y(n4612) );
  OA21X1_LVT U6130 ( .A1(n_T_698[31]), .A2(n9502), .A3(n4600), .Y(n4601) );
  OA21X1_LVT U6131 ( .A1(n_T_698[32]), .A2(n9505), .A3(n4601), .Y(n4611) );
  OAI22X1_LVT U6132 ( .A1(n_T_698[27]), .A2(n9489), .A3(n_T_698[29]), .A4(
        n9504), .Y(n4608) );
  OA22X1_LVT U6133 ( .A1(n_T_698[19]), .A2(n9510), .A3(n_T_698[25]), .A4(n9497), .Y(n4604) );
  NAND4X0_LVT U6134 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .Y(n4607) );
  NOR4X1_LVT U6135 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .Y(n4610)
         );
  NAND4X0_LVT U6136 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n3204), .Y(n4613) );
  NOR3X0_LVT U6137 ( .A1(ex_reg_valid), .A2(ex_reg_replay), .A3(
        ex_reg_xcpt_interrupt), .Y(n9426) );
  INVX1_LVT U6138 ( .A(n9426), .Y(n5089) );
  MUX21X1_LVT U6139 ( .A1(n4614), .A2(n4613), .S0(n5089), .Y(
        io_imem_bht_update_bits_mispredict) );
  AND2X1_LVT U6140 ( .A1(ibuf_io_inst_0_valid), .A2(n9418), .Y(n9417) );
  NAND3X0_LVT U6141 ( .A1(n4618), .A2(io_fpu_dec_ren1), .A3(n4846), .Y(n4638)
         );
  AND4X1_LVT U6142 ( .A1(n4622), .A2(n4621), .A3(n4620), .A4(n4619), .Y(n4947)
         );
  NAND3X0_LVT U6143 ( .A1(n4947), .A2(io_fpu_dec_wen), .A3(n4946), .Y(n4637)
         );
  NAND4X0_LVT U6144 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(io_fpu_dec_ren3), 
        .Y(n4626) );
  OR3X1_LVT U6145 ( .A1(n4628), .A2(n4627), .A3(n4626), .Y(n4636) );
  NAND4X0_LVT U6146 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .Y(n4858) );
  NAND3X0_LVT U6147 ( .A1(n4634), .A2(io_fpu_dec_ren2), .A3(n4633), .Y(n4635)
         );
  NAND4X0_LVT U6148 ( .A1(n4638), .A2(n4637), .A3(n4636), .A4(n4635), .Y(n4639) );
  AO21X1_LVT U6149 ( .A1(mem_ctrl_wfd), .A2(n4639), .A3(csr_io_singleStep), 
        .Y(n4640) );
  NAND2X0_LVT U6150 ( .A1(n4640), .A2(mem_reg_valid), .Y(n4746) );
  OA22X1_LVT U6151 ( .A1(n3124), .A2(n4708), .A3(n3086), .A4(n4675), .Y(n4645)
         );
  NAND2X0_LVT U6152 ( .A1(n4729), .A2(n_T_1298[2]), .Y(n4644) );
  NAND2X0_LVT U6153 ( .A1(n4731), .A2(n_T_1298[0]), .Y(n4643) );
  NAND3X0_LVT U6154 ( .A1(n4645), .A2(n4644), .A3(n4643), .Y(n4650) );
  OA22X1_LVT U6155 ( .A1(n3125), .A2(n4708), .A3(n3088), .A4(n4675), .Y(n4648)
         );
  NAND2X0_LVT U6156 ( .A1(n4729), .A2(n_T_1298[6]), .Y(n4647) );
  NAND2X0_LVT U6157 ( .A1(n4731), .A2(n_T_1298[4]), .Y(n4646) );
  NAND3X0_LVT U6158 ( .A1(n4648), .A2(n4647), .A3(n4646), .Y(n4649) );
  MUX21X1_LVT U6159 ( .A1(n4650), .A2(n4649), .S0(
        ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4661) );
  NAND2X0_LVT U6160 ( .A1(n4731), .A2(n_T_1298[8]), .Y(n4652) );
  NAND2X0_LVT U6161 ( .A1(n4732), .A2(n_T_1298[9]), .Y(n4651) );
  NAND4X0_LVT U6162 ( .A1(n4652), .A2(n4651), .A3(n4733), .A4(n4719), .Y(n4659) );
  AO22X1_LVT U6163 ( .A1(n_T_1298[11]), .A2(n4730), .A3(n4729), .A4(
        n_T_1298[10]), .Y(n4658) );
  AO22X1_LVT U6164 ( .A1(n_T_1298[15]), .A2(n4730), .A3(n4731), .A4(
        n_T_1298[12]), .Y(n4656) );
  NAND2X0_LVT U6165 ( .A1(n4732), .A2(n_T_1298[13]), .Y(n4654) );
  NAND2X0_LVT U6166 ( .A1(n4729), .A2(n_T_1298[14]), .Y(n4653) );
  NAND3X0_LVT U6167 ( .A1(n4654), .A2(ibuf_io_inst_0_bits_inst_rd[2]), .A3(
        n4653), .Y(n4655) );
  OA21X1_LVT U6168 ( .A1(n4656), .A2(n4655), .A3(
        ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4657) );
  OA22X1_LVT U6169 ( .A1(n4659), .A2(n4658), .A3(
        ibuf_io_inst_0_bits_inst_rd[4]), .A4(n4657), .Y(n4660) );
  AO21X1_LVT U6170 ( .A1(n4662), .A2(n4661), .A3(n4660), .Y(n4683) );
  OA22X1_LVT U6171 ( .A1(n3126), .A2(n4708), .A3(n3087), .A4(n4675), .Y(n4665)
         );
  AND2X1_LVT U6172 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n4662), .Y(n4666) );
  AND2X1_LVT U6173 ( .A1(n4666), .A2(n4733), .Y(n4717) );
  NAND2X0_LVT U6174 ( .A1(n4731), .A2(n_T_1298[16]), .Y(n4664) );
  NAND2X0_LVT U6175 ( .A1(n4729), .A2(n_T_1298[18]), .Y(n4663) );
  NAND4X0_LVT U6176 ( .A1(n4665), .A2(n4717), .A3(n4664), .A4(n4663), .Y(n4671) );
  OA22X1_LVT U6177 ( .A1(n3239), .A2(n4708), .A3(n3114), .A4(n4675), .Y(n4669)
         );
  AND2X1_LVT U6178 ( .A1(n4666), .A2(ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4698) );
  NAND2X0_LVT U6179 ( .A1(n4731), .A2(n_T_1298[20]), .Y(n4668) );
  NAND2X0_LVT U6180 ( .A1(n4729), .A2(n_T_1298[22]), .Y(n4667) );
  NAND4X0_LVT U6181 ( .A1(n4669), .A2(n4698), .A3(n4668), .A4(n4667), .Y(n4670) );
  NAND2X0_LVT U6182 ( .A1(n1699), .A2(n3039), .Y(n9286) );
  AND4X1_LVT U6183 ( .A1(n4671), .A2(n4670), .A3(io_fpu_dec_wen), .A4(n9286), 
        .Y(n4682) );
  OA22X1_LVT U6184 ( .A1(n3085), .A2(n4708), .A3(n3116), .A4(n4675), .Y(n4674)
         );
  AND2X1_LVT U6185 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(
        ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4676) );
  AND2X1_LVT U6186 ( .A1(n4733), .A2(n4676), .Y(n4711) );
  NAND2X0_LVT U6187 ( .A1(n4731), .A2(n_T_1298[24]), .Y(n4673) );
  NAND2X0_LVT U6188 ( .A1(n4729), .A2(n_T_1298[26]), .Y(n4672) );
  NAND4X0_LVT U6189 ( .A1(n4674), .A2(n4711), .A3(n4673), .A4(n4672), .Y(n4681) );
  OA22X1_LVT U6190 ( .A1(n3241), .A2(n4708), .A3(n3084), .A4(n4675), .Y(n4679)
         );
  AND2X1_LVT U6191 ( .A1(n4676), .A2(ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4727) );
  NAND2X0_LVT U6192 ( .A1(n4731), .A2(n_T_1298[28]), .Y(n4678) );
  NAND2X0_LVT U6193 ( .A1(n4729), .A2(n_T_1298[30]), .Y(n4677) );
  NAND4X0_LVT U6194 ( .A1(n4679), .A2(n4727), .A3(n4678), .A4(n4677), .Y(n4680) );
  NAND4X0_LVT U6195 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .Y(n4745) );
  AND2X1_LVT U6196 ( .A1(n4700), .A2(n4733), .Y(n4691) );
  NAND2X0_LVT U6197 ( .A1(n4691), .A2(n4731), .Y(n4684) );
  AND2X1_LVT U6198 ( .A1(id_ctrl_wxd), .A2(n4684), .Y(n5054) );
  NAND2X0_LVT U6199 ( .A1(n4687), .A2(n4686), .Y(n4696) );
  NAND2X0_LVT U6200 ( .A1(wb_ctrl_wxd), .A2(wb_reg_valid), .Y(n5402) );
  NAND2X0_LVT U6201 ( .A1(div_io_resp_valid), .A2(n5402), .Y(n5415) );
  AO21X1_LVT U6202 ( .A1(n_T_1187[3]), .A2(n4730), .A3(n4692), .Y(n4694) );
  AO22X1_LVT U6203 ( .A1(n4729), .A2(n_T_1187[2]), .A3(n_T_1187[1]), .A4(n4732), .Y(n4693) );
  OA22X1_LVT U6204 ( .A1(n4696), .A2(n4695), .A3(n4694), .A4(n4693), .Y(n4715)
         );
  AO22X1_LVT U6205 ( .A1(n_T_1187[23]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[22]), .Y(n4706) );
  NAND2X0_LVT U6206 ( .A1(n4731), .A2(n_T_1187[20]), .Y(n4699) );
  NAND2X0_LVT U6207 ( .A1(n4732), .A2(n_T_1187[21]), .Y(n4697) );
  NAND3X0_LVT U6208 ( .A1(n4699), .A2(n4698), .A3(n4697), .Y(n4705) );
  AO22X1_LVT U6209 ( .A1(n_T_1187[7]), .A2(n4730), .A3(n4729), .A4(n_T_1187[6]), .Y(n4704) );
  NAND2X0_LVT U6210 ( .A1(n4731), .A2(n_T_1187[4]), .Y(n4702) );
  NAND2X0_LVT U6211 ( .A1(n4732), .A2(n_T_1187[5]), .Y(n4701) );
  NAND4X0_LVT U6212 ( .A1(n4702), .A2(n4701), .A3(
        ibuf_io_inst_0_bits_inst_rd[2]), .A4(n4700), .Y(n4703) );
  OA22X1_LVT U6213 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .Y(n4714)
         );
  OA22X1_LVT U6214 ( .A1(n3135), .A2(n4708), .A3(n3265), .A4(n4707), .Y(n4712)
         );
  NAND2X0_LVT U6215 ( .A1(n4732), .A2(n_T_1187[25]), .Y(n4710) );
  NAND2X0_LVT U6216 ( .A1(n4731), .A2(n_T_1187[24]), .Y(n4709) );
  NAND4X0_LVT U6217 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .Y(n4713) );
  AND4X1_LVT U6218 ( .A1(n5054), .A2(n4715), .A3(n4714), .A4(n4713), .Y(n4743)
         );
  AO22X1_LVT U6219 ( .A1(n_T_1187[19]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[18]), .Y(n4725) );
  NAND2X0_LVT U6220 ( .A1(n4731), .A2(n_T_1187[16]), .Y(n4718) );
  NAND2X0_LVT U6221 ( .A1(n4732), .A2(n_T_1187[17]), .Y(n4716) );
  NAND3X0_LVT U6222 ( .A1(n4718), .A2(n4717), .A3(n4716), .Y(n4724) );
  AO22X1_LVT U6223 ( .A1(n_T_1187[15]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[14]), .Y(n4723) );
  NAND2X0_LVT U6224 ( .A1(n4731), .A2(n_T_1187[12]), .Y(n4721) );
  NAND2X0_LVT U6225 ( .A1(n4732), .A2(n_T_1187[13]), .Y(n4720) );
  AND2X1_LVT U6226 ( .A1(n4719), .A2(ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4734) );
  NAND4X0_LVT U6227 ( .A1(n4721), .A2(n4720), .A3(
        ibuf_io_inst_0_bits_inst_rd[2]), .A4(n4734), .Y(n4722) );
  OA22X1_LVT U6228 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .Y(n4742)
         );
  AO22X1_LVT U6229 ( .A1(n_T_1187[31]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[30]), .Y(n4740) );
  NAND2X0_LVT U6230 ( .A1(n4731), .A2(n_T_1187[28]), .Y(n4728) );
  NAND2X0_LVT U6231 ( .A1(n4732), .A2(n_T_1187[29]), .Y(n4726) );
  NAND3X0_LVT U6232 ( .A1(n4728), .A2(n4727), .A3(n4726), .Y(n4739) );
  AO22X1_LVT U6233 ( .A1(n_T_1187[11]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[10]), .Y(n4738) );
  NAND2X0_LVT U6234 ( .A1(n4731), .A2(n_T_1187[8]), .Y(n4736) );
  NAND2X0_LVT U6235 ( .A1(n4732), .A2(n_T_1187[9]), .Y(n4735) );
  NAND4X0_LVT U6236 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .Y(n4737) );
  OA22X1_LVT U6237 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .Y(n4741)
         );
  NAND3X0_LVT U6238 ( .A1(n4743), .A2(n4742), .A3(n4741), .Y(n4744) );
  NAND3X0_LVT U6239 ( .A1(n4746), .A2(n4745), .A3(n4744), .Y(n9285) );
  AND2X1_LVT U6240 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n2877), .Y(
        n4971) );
  NAND2X0_LVT U6241 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n2790), .Y(
        n4968) );
  INVX1_LVT U6242 ( .A(n4968), .Y(n4749) );
  AO22X1_LVT U6243 ( .A1(n6972), .A2(n_T_1298[3]), .A3(n6974), .A4(n_T_1298[1]), .Y(n4756) );
  AND2X1_LVT U6244 ( .A1(n4747), .A2(n2876), .Y(n4970) );
  AO22X1_LVT U6245 ( .A1(n6946), .A2(n_T_1298[7]), .A3(n6931), .A4(n_T_1298[6]), .Y(n4755) );
  NAND2X0_LVT U6246 ( .A1(n6957), .A2(n_T_1298[0]), .Y(n4751) );
  NAND2X0_LVT U6247 ( .A1(n6954), .A2(n_T_1298[5]), .Y(n4750) );
  NAND4X0_LVT U6248 ( .A1(n4751), .A2(n6963), .A3(n4750), .A4(n6956), .Y(n4754) );
  AO22X1_LVT U6249 ( .A1(n6926), .A2(n_T_1298[4]), .A3(n6948), .A4(n_T_1298[2]), .Y(n4753) );
  AO22X1_LVT U6250 ( .A1(n6972), .A2(n_T_1298[11]), .A3(n6946), .A4(
        n_T_1298[15]), .Y(n4762) );
  AO22X1_LVT U6251 ( .A1(n6974), .A2(n_T_1298[9]), .A3(n6926), .A4(
        n_T_1298[12]), .Y(n4761) );
  AO22X1_LVT U6252 ( .A1(n6957), .A2(n_T_1298[8]), .A3(n6948), .A4(
        n_T_1298[10]), .Y(n4760) );
  NAND2X0_LVT U6253 ( .A1(n6931), .A2(n_T_1298[14]), .Y(n4758) );
  NAND2X0_LVT U6254 ( .A1(n6954), .A2(n_T_1298[13]), .Y(n4757) );
  AO22X1_LVT U6255 ( .A1(n6946), .A2(n_T_1298[23]), .A3(n6957), .A4(
        n_T_1298[16]), .Y(n4768) );
  AO22X1_LVT U6256 ( .A1(n6974), .A2(n_T_1298[17]), .A3(n6954), .A4(
        n_T_1298[21]), .Y(n4767) );
  OA22X1_LVT U6257 ( .A1(n3238), .A2(n6955), .A3(n3117), .A4(n6947), .Y(n4765)
         );
  AND2X1_LVT U6258 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n6956), .Y(
        n6924) );
  NAND2X0_LVT U6259 ( .A1(n6948), .A2(n_T_1298[18]), .Y(n4764) );
  NAND2X0_LVT U6260 ( .A1(n6972), .A2(n_T_1298[19]), .Y(n4763) );
  OR3X1_LVT U6261 ( .A1(n4766), .A2(n4767), .A3(n4768), .Y(n4780) );
  NAND2X0_LVT U6262 ( .A1(n6974), .A2(n_T_1298[25]), .Y(n4770) );
  AND2X1_LVT U6263 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n2825), .Y(
        n6917) );
  NAND2X0_LVT U6264 ( .A1(n6946), .A2(n_T_1298[31]), .Y(n4769) );
  AND3X1_LVT U6265 ( .A1(n4770), .A2(n6917), .A3(n4769), .Y(n4778) );
  OA22X1_LVT U6266 ( .A1(n3237), .A2(n4771), .A3(n3123), .A4(n6955), .Y(n4777)
         );
  OA22X1_LVT U6267 ( .A1(n3084), .A2(n4772), .A3(n3118), .A4(n6947), .Y(n4776)
         );
  OA22X1_LVT U6268 ( .A1(n4774), .A2(n3085), .A3(n3232), .A4(n4773), .Y(n4775)
         );
  NAND4X0_LVT U6269 ( .A1(n4778), .A2(n4777), .A3(n4776), .A4(n4775), .Y(n4779) );
  NAND2X0_LVT U6270 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(
        ibuf_io_inst_0_bits_raw[27]), .Y(n4802) );
  OA22X1_LVT U6271 ( .A1(n3124), .A2(n4802), .A3(n3247), .A4(n4801), .Y(n4784)
         );
  OA22X1_LVT U6272 ( .A1(n3254), .A2(n4804), .A3(n3086), .A4(n4803), .Y(n4783)
         );
  AND2X1_LVT U6273 ( .A1(n4784), .A2(n4783), .Y(n4794) );
  OA22X1_LVT U6274 ( .A1(n3240), .A2(n4802), .A3(n3115), .A4(n4801), .Y(n4786)
         );
  OA22X1_LVT U6275 ( .A1(n3242), .A2(n4804), .A3(n3119), .A4(n4803), .Y(n4785)
         );
  AND2X1_LVT U6276 ( .A1(n4786), .A2(n4785), .Y(n4793) );
  OA22X1_LVT U6277 ( .A1(n3125), .A2(n4802), .A3(n3248), .A4(n4801), .Y(n4788)
         );
  OA22X1_LVT U6278 ( .A1(n3253), .A2(n4804), .A3(n3088), .A4(n4803), .Y(n4787)
         );
  AND2X1_LVT U6279 ( .A1(n4788), .A2(n4787), .Y(n4792) );
  OA22X1_LVT U6280 ( .A1(n3236), .A2(n4802), .A3(n3121), .A4(n4801), .Y(n4790)
         );
  OA22X1_LVT U6281 ( .A1(n3235), .A2(n4804), .A3(n3120), .A4(n4803), .Y(n4789)
         );
  AND2X1_LVT U6282 ( .A1(n4790), .A2(n4789), .Y(n4791) );
  MUX41X1_LVT U6283 ( .A1(n4794), .A3(n4793), .A2(n4792), .A4(n4791), .S0(
        n1859), .S1(ibuf_io_inst_0_bits_inst_rs3_2_), .Y(n4812) );
  OA22X1_LVT U6284 ( .A1(n3126), .A2(n4802), .A3(n3250), .A4(n4801), .Y(n4796)
         );
  OA22X1_LVT U6285 ( .A1(n3252), .A2(n4804), .A3(n3087), .A4(n4803), .Y(n4795)
         );
  AND2X1_LVT U6286 ( .A1(n4796), .A2(n4795), .Y(n4810) );
  OA22X1_LVT U6287 ( .A1(n3085), .A2(n4802), .A3(n3232), .A4(n4801), .Y(n4798)
         );
  OA22X1_LVT U6288 ( .A1(n3237), .A2(n4804), .A3(n3116), .A4(n4803), .Y(n4797)
         );
  AND2X1_LVT U6289 ( .A1(n4798), .A2(n4797), .Y(n4809) );
  OA22X1_LVT U6290 ( .A1(n3239), .A2(n4802), .A3(n3117), .A4(n4801), .Y(n4800)
         );
  OA22X1_LVT U6291 ( .A1(n3238), .A2(n4804), .A3(n3114), .A4(n4803), .Y(n4799)
         );
  AND2X1_LVT U6292 ( .A1(n4800), .A2(n4799), .Y(n4808) );
  OA22X1_LVT U6293 ( .A1(n3241), .A2(n4802), .A3(n3118), .A4(n4801), .Y(n4806)
         );
  OA22X1_LVT U6294 ( .A1(n3123), .A2(n4804), .A3(n3084), .A4(n4803), .Y(n4805)
         );
  AND2X1_LVT U6295 ( .A1(n4806), .A2(n4805), .Y(n4807) );
  MUX41X1_LVT U6296 ( .A1(n4810), .A3(n4809), .A2(n4808), .A4(n4807), .S0(
        n1859), .S1(ibuf_io_inst_0_bits_raw[29]), .Y(n4811) );
  AND2X1_LVT U6297 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(
        ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n4889) );
  AO22X1_LVT U6298 ( .A1(n_T_1298[3]), .A2(n5452), .A3(n5455), .A4(n_T_1298[0]), .Y(n4820) );
  AND2X1_LVT U6299 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n4813), .Y(
        n4890) );
  AO22X1_LVT U6300 ( .A1(n_T_1298[7]), .A2(n5450), .A3(n5456), .A4(n_T_1298[1]), .Y(n4819) );
  AND2X1_LVT U6301 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n4815), .Y(
        n4900) );
  AO22X1_LVT U6302 ( .A1(n2034), .A2(n_T_1298[4]), .A3(n_T_1298[6]), .A4(n5449), .Y(n4818) );
  AO22X1_LVT U6303 ( .A1(n5451), .A2(n_T_1298[5]), .A3(n_T_1298[2]), .A4(n5454), .Y(n4817) );
  NOR4X1_LVT U6304 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .Y(n4835)
         );
  OA22X1_LVT U6305 ( .A1(n3236), .A2(n5438), .A3(n3119), .A4(n4905), .Y(n4824)
         );
  INVX1_LVT U6306 ( .A(n5453), .Y(n4880) );
  OA22X1_LVT U6307 ( .A1(n3235), .A2(n4880), .A3(n3115), .A4(n4873), .Y(n4823)
         );
  OA22X1_LVT U6308 ( .A1(n3240), .A2(n4906), .A3(n3120), .A4(n4894), .Y(n4822)
         );
  OA22X1_LVT U6309 ( .A1(n3242), .A2(n5435), .A3(n3121), .A4(n4874), .Y(n4821)
         );
  AO22X1_LVT U6310 ( .A1(n_T_1298[19]), .A2(n5452), .A3(n5454), .A4(
        n_T_1298[18]), .Y(n4828) );
  AO22X1_LVT U6311 ( .A1(n_T_1298[23]), .A2(n5450), .A3(n2034), .A4(
        n_T_1298[20]), .Y(n4827) );
  AO22X1_LVT U6312 ( .A1(n5455), .A2(n_T_1298[16]), .A3(n_T_1298[22]), .A4(
        n5449), .Y(n4826) );
  AO22X1_LVT U6313 ( .A1(n5451), .A2(n_T_1298[21]), .A3(n_T_1298[17]), .A4(
        n5456), .Y(n4825) );
  NOR4X1_LVT U6314 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), .Y(n4834)
         );
  AO22X1_LVT U6315 ( .A1(n_T_1298[27]), .A2(n5452), .A3(n5456), .A4(
        n_T_1298[25]), .Y(n4832) );
  AO22X1_LVT U6316 ( .A1(n_T_1298[31]), .A2(n5450), .A3(n5455), .A4(
        n_T_1298[24]), .Y(n4831) );
  AO22X1_LVT U6317 ( .A1(n2034), .A2(n_T_1298[28]), .A3(n_T_1298[30]), .A4(
        n5449), .Y(n4830) );
  AO22X1_LVT U6318 ( .A1(n5451), .A2(n_T_1298[29]), .A3(n_T_1298[26]), .A4(
        n5454), .Y(n4829) );
  NOR4X1_LVT U6319 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), .Y(n4833)
         );
  MUX41X1_LVT U6320 ( .A1(n4835), .A3(n3181), .A2(n4834), .A4(n4833), .S0(
        n3781), .S1(ibuf_io_inst_0_bits_inst_rs2[4]), .Y(n4836) );
  OA22X1_LVT U6321 ( .A1(n4839), .A2(n4838), .A3(n4837), .A4(n4836), .Y(n4849)
         );
  NAND2X0_LVT U6322 ( .A1(mem_ctrl_mem), .A2(mem_reg_slow_bypass), .Y(n4840)
         );
  NAND3X0_LVT U6323 ( .A1(n4840), .A2(n370), .A3(n3246), .Y(n4841) );
  NOR4X1_LVT U6324 ( .A1(mem_ctrl_csr[0]), .A2(mem_ctrl_csr[2]), .A3(n3279), 
        .A4(n4841), .Y(n4949) );
  NAND2X0_LVT U6325 ( .A1(n5163), .A2(io_fpu_inst[14]), .Y(n4842) );
  NAND2X0_LVT U6326 ( .A1(n2538), .A2(n9288), .Y(n9280) );
  AND2X1_LVT U6327 ( .A1(mem_ctrl_wxd), .A2(mem_reg_valid), .Y(n4948) );
  NAND2X0_LVT U6328 ( .A1(n4846), .A2(n4948), .Y(n4848) );
  OA22X1_LVT U6329 ( .A1(n2512), .A2(n4849), .A3(n4949), .A4(n5094), .Y(n4851)
         );
  NAND2X0_LVT U6330 ( .A1(n1612), .A2(n9432), .Y(n5087) );
  NAND3X0_LVT U6331 ( .A1(n5087), .A2(blocked), .A3(n5065), .Y(n4850) );
  AND3X1_LVT U6332 ( .A1(n4850), .A2(n4851), .A3(n4852), .Y(n4955) );
  AND2X1_LVT U6333 ( .A1(n5396), .A2(n2618), .Y(n1828) );
  NAND2X0_LVT U6334 ( .A1(n5087), .A2(id_reg_fence), .Y(n4854) );
  AND2X1_LVT U6335 ( .A1(ex_ctrl_mem), .A2(ex_reg_valid), .Y(io_dmem_req_valid) );
  INVX1_LVT U6336 ( .A(io_dmem_req_valid), .Y(n4853) );
  AND2X1_LVT U6337 ( .A1(n4853), .A2(io_dmem_ordered), .Y(n5063) );
  AO21X1_LVT U6338 ( .A1(n4855), .A2(n4854), .A3(n5063), .Y(n4954) );
  NAND2X0_LVT U6339 ( .A1(n4856), .A2(n3597), .Y(n4857) );
  NAND2X0_LVT U6340 ( .A1(n1531), .A2(n1532), .Y(n5466) );
  AND2X1_LVT U6341 ( .A1(n5466), .A2(n5421), .Y(n5021) );
  NOR3X0_LVT U6342 ( .A1(n4860), .A2(n4859), .A3(n4858), .Y(n5420) );
  NAND2X0_LVT U6343 ( .A1(n5021), .A2(n5420), .Y(n5093) );
  INVX1_LVT U6344 ( .A(n5044), .Y(n4867) );
  AND2X1_LVT U6345 ( .A1(ex_reg_valid), .A2(ex_ctrl_wxd), .Y(n5009) );
  AND4X1_LVT U6346 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .Y(n5045)
         );
  INVX1_LVT U6347 ( .A(n5045), .Y(n4865) );
  OR3X1_LVT U6348 ( .A1(n4867), .A2(n4866), .A3(n4865), .Y(n5419) );
  NAND2X0_LVT U6349 ( .A1(n4872), .A2(n4871), .Y(n4887) );
  OA22X1_LVT U6350 ( .A1(n3272), .A2(n4894), .A3(n3129), .A4(n4873), .Y(n4878)
         );
  OA22X1_LVT U6351 ( .A1(n3260), .A2(n4880), .A3(n3127), .A4(n4874), .Y(n4877)
         );
  OA22X1_LVT U6352 ( .A1(n4906), .A2(n3259), .A3(n3133), .A4(n4905), .Y(n4876)
         );
  OA22X1_LVT U6353 ( .A1(n5438), .A2(n3266), .A3(n3134), .A4(n5435), .Y(n4875)
         );
  NAND4X0_LVT U6354 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .Y(n4879) );
  AND2X1_LVT U6355 ( .A1(n4879), .A2(n2878), .Y(n4886) );
  NAND2X0_LVT U6356 ( .A1(n5451), .A2(n5436), .Y(n5546) );
  OA22X1_LVT U6357 ( .A1(n3271), .A2(n5546), .A3(n3136), .A4(n6766), .Y(n4884)
         );
  NAND2X0_LVT U6358 ( .A1(n5454), .A2(n5436), .Y(n6422) );
  NAND2X0_LVT U6359 ( .A1(n5452), .A2(n5436), .Y(n5906) );
  NAND2X0_LVT U6360 ( .A1(n5456), .A2(n5436), .Y(n5905) );
  NAND2X0_LVT U6361 ( .A1(n5450), .A2(n5436), .Y(n6767) );
  OA22X1_LVT U6362 ( .A1(n3270), .A2(n6767), .A3(n3132), .A4(n6423), .Y(n4881)
         );
  NAND4X0_LVT U6363 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n4881), .Y(n4885) );
  OAI22X1_LVT U6364 ( .A1(n4888), .A2(n4887), .A3(n4886), .A4(n4885), .Y(n4916) );
  OA22X1_LVT U6365 ( .A1(n4899), .A2(n3267), .A3(n3131), .A4(n4898), .Y(n4893)
         );
  NAND2X0_LVT U6366 ( .A1(n4901), .A2(n_T_1187[28]), .Y(n4892) );
  NAND2X0_LVT U6367 ( .A1(n4900), .A2(n_T_1187[30]), .Y(n4891) );
  OA22X1_LVT U6368 ( .A1(n5438), .A2(n3268), .A3(n3130), .A4(n4894), .Y(n4897)
         );
  NAND2X0_LVT U6369 ( .A1(n2034), .A2(n_T_1187[20]), .Y(n4896) );
  NAND2X0_LVT U6370 ( .A1(n5449), .A2(n_T_1187[22]), .Y(n4895) );
  NAND3X0_LVT U6371 ( .A1(n4897), .A2(n4896), .A3(n4895), .Y(n4913) );
  OA22X1_LVT U6372 ( .A1(n4899), .A2(n3135), .A3(n3089), .A4(n4898), .Y(n4904)
         );
  NAND2X0_LVT U6373 ( .A1(n4900), .A2(n_T_1187[26]), .Y(n4903) );
  NAND2X0_LVT U6374 ( .A1(n4901), .A2(n_T_1187[24]), .Y(n4902) );
  MUX21X1_LVT U6375 ( .A1(n4910), .A2(n4914), .S0(
        ibuf_io_inst_0_bits_inst_rs2[2]), .Y(n4912) );
  OA22X1_LVT U6376 ( .A1(n4906), .A2(n3258), .A3(n3113), .A4(n4905), .Y(n4909)
         );
  NAND2X0_LVT U6377 ( .A1(n5455), .A2(n_T_1187[16]), .Y(n4908) );
  NAND2X0_LVT U6378 ( .A1(n5454), .A2(n_T_1187[18]), .Y(n4907) );
  NAND3X0_LVT U6379 ( .A1(n4909), .A2(n4908), .A3(n4907), .Y(n4911) );
  AOI222X1_LVT U6380 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n5447), .A5(
        n4911), .A6(n4910), .Y(n4915) );
  OA22X1_LVT U6381 ( .A1(n5051), .A2(n5419), .A3(n4916), .A4(n4915), .Y(n4935)
         );
  AND2X1_LVT U6382 ( .A1(ex_reg_valid), .A2(ex_ctrl_div), .Y(n9422) );
  AO21X1_LVT U6383 ( .A1(n5415), .A2(n4917), .A3(n9422), .Y(n4932) );
  NOR2X0_LVT U6384 ( .A1(id_reg_pause), .A2(csr_io_csr_stall), .Y(n4928) );
  AND3X1_LVT U6385 ( .A1(wb_ctrl_wfd), .A2(wb_reg_valid), .A3(io_fpu_dec_ren3), 
        .Y(n4919) );
  NAND4X0_LVT U6386 ( .A1(n4922), .A2(n4921), .A3(n4920), .A4(n4919), .Y(n4923) );
  OR3X1_LVT U6387 ( .A1(n4925), .A2(n4924), .A3(n4923), .Y(n4927) );
  NAND2X0_LVT U6388 ( .A1(csr_io_singleStep), .A2(wb_reg_valid), .Y(n4926) );
  NAND4X0_LVT U6389 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .Y(n4930) );
  AOI21X1_LVT U6390 ( .A1(n4932), .A2(n4931), .A3(n4930), .Y(n4933) );
  OA21X1_LVT U6391 ( .A1(n4935), .A2(n4934), .A3(n4933), .Y(n4936) );
  OA21X1_LVT U6392 ( .A1(n4949), .A2(n5093), .A3(n4936), .Y(n4953) );
  NAND4X0_LVT U6393 ( .A1(n4939), .A2(n4938), .A3(n4937), .A4(wb_reg_valid), 
        .Y(n4940) );
  OR3X1_LVT U6394 ( .A1(n4942), .A2(n4941), .A3(n4940), .Y(n4951) );
  AND2X1_LVT U6395 ( .A1(n4943), .A2(wb_ctrl_mem), .Y(n5175) );
  OA21X1_LVT U6396 ( .A1(wb_ctrl_div), .A2(n5175), .A3(wb_ctrl_wxd), .Y(n5301)
         );
  OA22X1_LVT U6397 ( .A1(n4945), .A2(n3229), .A3(n4944), .A4(n9280), .Y(n4950)
         );
  NAND4X0_LVT U6398 ( .A1(n5054), .A2(n4948), .A3(n4947), .A4(n4946), .Y(n5092) );
  OA22X1_LVT U6399 ( .A1(n4951), .A2(n4950), .A3(n4949), .A4(n5092), .Y(n4952)
         );
  OA22X1_LVT U6400 ( .A1(n3261), .A2(n4969), .A3(n3113), .A4(n4968), .Y(n4958)
         );
  NAND2X0_LVT U6401 ( .A1(n4970), .A2(n_T_1187[18]), .Y(n4957) );
  NAND2X0_LVT U6402 ( .A1(n4971), .A2(n_T_1187[19]), .Y(n4956) );
  NAND3X0_LVT U6403 ( .A1(n4958), .A2(n4957), .A3(n4956), .Y(n4963) );
  OA22X1_LVT U6404 ( .A1(n3275), .A2(n4969), .A3(n3089), .A4(n4968), .Y(n4961)
         );
  NAND2X0_LVT U6405 ( .A1(n4970), .A2(n_T_1187[26]), .Y(n4960) );
  NAND2X0_LVT U6406 ( .A1(n4971), .A2(n_T_1187[27]), .Y(n4959) );
  NAND3X0_LVT U6407 ( .A1(n4961), .A2(n4960), .A3(n4959), .Y(n4962) );
  MUX21X1_LVT U6408 ( .A1(n4963), .A2(n4962), .S0(n2825), .Y(n4964) );
  OR2X1_LVT U6409 ( .A1(n6963), .A2(n4964), .Y(n4979) );
  OA22X1_LVT U6410 ( .A1(n3273), .A2(n4969), .A3(n3130), .A4(n4968), .Y(n4967)
         );
  NAND2X0_LVT U6411 ( .A1(n4970), .A2(n_T_1187[22]), .Y(n4966) );
  NAND2X0_LVT U6412 ( .A1(n4971), .A2(n_T_1187[23]), .Y(n4965) );
  NAND3X0_LVT U6413 ( .A1(n4967), .A2(n4966), .A3(n4965), .Y(n4976) );
  OA22X1_LVT U6414 ( .A1(n3274), .A2(n4969), .A3(n3131), .A4(n4968), .Y(n4974)
         );
  NAND2X0_LVT U6415 ( .A1(n4970), .A2(n_T_1187[30]), .Y(n4973) );
  NAND2X0_LVT U6416 ( .A1(n4971), .A2(n_T_1187[31]), .Y(n4972) );
  NAND3X0_LVT U6417 ( .A1(n4974), .A2(n4973), .A3(n4972), .Y(n4975) );
  MUX21X1_LVT U6418 ( .A1(n4976), .A2(n4975), .S0(n2825), .Y(n4977) );
  OR2X1_LVT U6419 ( .A1(n6963), .A2(n4977), .Y(n4978) );
  MUX21X1_LVT U6420 ( .A1(n4979), .A2(n4978), .S0(n2038), .Y(n5008) );
  OA21X1_LVT U6421 ( .A1(n3132), .A2(n6949), .A3(n6963), .Y(n4982) );
  NAND2X0_LVT U6422 ( .A1(n4044), .A2(n_T_1187[2]), .Y(n4981) );
  AND2X1_LVT U6423 ( .A1(n6946), .A2(n6956), .Y(n8931) );
  NAND2X0_LVT U6424 ( .A1(n3968), .A2(n_T_1187[7]), .Y(n4980) );
  NAND3X0_LVT U6425 ( .A1(n4982), .A2(n4980), .A3(n4981), .Y(n4999) );
  NAND2X0_LVT U6426 ( .A1(n6974), .A2(n6956), .Y(n6945) );
  NAND2X0_LVT U6427 ( .A1(n3972), .A2(n_T_1187[3]), .Y(n4983) );
  OA21X1_LVT U6428 ( .A1(n3128), .A2(n6945), .A3(n4983), .Y(n4986) );
  AND2X1_LVT U6429 ( .A1(n6954), .A2(n6956), .Y(n8901) );
  NAND2X0_LVT U6430 ( .A1(n3967), .A2(n_T_1187[5]), .Y(n4985) );
  NAND2X0_LVT U6431 ( .A1(n9040), .A2(n_T_1187[6]), .Y(n4984) );
  NAND3X0_LVT U6432 ( .A1(n4986), .A2(n4984), .A3(n4985), .Y(n4998) );
  NAND2X0_LVT U6433 ( .A1(n6972), .A2(n_T_1187[11]), .Y(n4987) );
  OA21X1_LVT U6434 ( .A1(n3127), .A2(n6947), .A3(n4987), .Y(n4990) );
  NAND2X0_LVT U6435 ( .A1(n6948), .A2(n_T_1187[10]), .Y(n4989) );
  NAND2X0_LVT U6436 ( .A1(n6974), .A2(n_T_1187[9]), .Y(n4988) );
  NAND3X0_LVT U6437 ( .A1(n4990), .A2(n4989), .A3(n4988), .Y(n4996) );
  NAND2X0_LVT U6438 ( .A1(n6946), .A2(n_T_1187[15]), .Y(n4991) );
  OA21X1_LVT U6439 ( .A1(n3260), .A2(n6955), .A3(n4991), .Y(n4994) );
  NAND2X0_LVT U6440 ( .A1(n6954), .A2(n_T_1187[13]), .Y(n4993) );
  NAND2X0_LVT U6441 ( .A1(n6957), .A2(n_T_1187[8]), .Y(n4992) );
  NAND3X0_LVT U6442 ( .A1(n4994), .A2(n4993), .A3(n4992), .Y(n4995) );
  OR3X1_LVT U6443 ( .A1(n4999), .A2(n4998), .A3(n4997), .Y(n5007) );
  OR3X1_LVT U6444 ( .A1(n5005), .A2(n5004), .A3(n5003), .Y(n5006) );
  NAND2X0_LVT U6445 ( .A1(n5037), .A2(n5009), .Y(n5013) );
  OA21X1_LVT U6446 ( .A1(n9280), .A2(n9281), .A3(n9385), .Y(n5029) );
  AO22X1_LVT U6447 ( .A1(wb_ctrl_wfd), .A2(io_fpu_dec_wen), .A3(n5054), .A4(
        n5301), .Y(n5020) );
  AND4X1_LVT U6448 ( .A1(n5016), .A2(wb_reg_valid), .A3(n5015), .A4(n5014), 
        .Y(n5019) );
  NAND4X0_LVT U6449 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .Y(n9278) );
  AO22X1_LVT U6450 ( .A1(io_fpu_dec_ren2), .A2(wb_ctrl_wfd), .A3(n5021), .A4(
        n5301), .Y(n5028) );
  AND4X1_LVT U6451 ( .A1(n5024), .A2(n5023), .A3(wb_reg_valid), .A4(n5022), 
        .Y(n5027) );
  NAND4X0_LVT U6452 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .Y(n9277) );
  AND3X1_LVT U6453 ( .A1(n5029), .A2(n9278), .A3(n9277), .Y(n5059) );
  AND2X1_LVT U6454 ( .A1(n5031), .A2(n5030), .Y(n5034) );
  AND4X1_LVT U6455 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5032), .Y(n5053)
         );
  NAND2X0_LVT U6456 ( .A1(n5053), .A2(io_fpu_dec_wen), .Y(n5049) );
  NAND3X0_LVT U6457 ( .A1(n2567), .A2(io_fpu_dec_ren1), .A3(n5037), .Y(n5048)
         );
  NAND4X0_LVT U6458 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(io_fpu_dec_ren3), 
        .Y(n5041) );
  OR3X1_LVT U6459 ( .A1(n5043), .A2(n5042), .A3(n5041), .Y(n5047) );
  NAND3X0_LVT U6460 ( .A1(n5045), .A2(io_fpu_dec_ren2), .A3(n5044), .Y(n5046)
         );
  NAND4X0_LVT U6461 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .Y(n5050) );
  NAND2X0_LVT U6462 ( .A1(n5050), .A2(ex_ctrl_wfd), .Y(n5057) );
  INVX1_LVT U6463 ( .A(csr_io_singleStep), .Y(n5056) );
  NAND4X0_LVT U6464 ( .A1(n5054), .A2(ex_ctrl_wxd), .A3(n5053), .A4(n5052), 
        .Y(n5055) );
  NAND3X0_LVT U6465 ( .A1(n5057), .A2(n5056), .A3(n5055), .Y(n5058) );
  NAND2X0_LVT U6466 ( .A1(n5058), .A2(ex_reg_valid), .Y(n9279) );
  NAND3X0_LVT U6467 ( .A1(n9279), .A2(n5059), .A3(n5060), .Y(n5061) );
  NOR3X0_LVT U6468 ( .A1(n5061), .A2(n9282), .A3(n9285), .Y(n5062) );
  NAND2X0_LVT U6469 ( .A1(io_dmem_req_valid), .A2(n5064), .Y(n5095) );
  NAND2X0_LVT U6470 ( .A1(n9521), .A2(io_fpu_inst[28]), .Y(n5154) );
  AND2X1_LVT U6471 ( .A1(n5066), .A2(io_fpu_inst[5]), .Y(n9431) );
  NAND2X0_LVT U6472 ( .A1(io_fpu_inst[3]), .A2(n5067), .Y(n9110) );
  AO21X1_LVT U6473 ( .A1(n9431), .A2(n5070), .A3(n5123), .Y(n9287) );
  NAND2X0_LVT U6474 ( .A1(n5071), .A2(n3597), .Y(n1628) );
  NAND2X0_LVT U6475 ( .A1(io_fpu_inst[13]), .A2(io_fpu_inst[4]), .Y(n9089) );
  AND2X1_LVT U6476 ( .A1(n2618), .A2(n5088), .Y(N286) );
  OA21X1_LVT U6477 ( .A1(n9105), .A2(n9520), .A3(n5072), .Y(n5073) );
  AND2X1_LVT U6478 ( .A1(n559), .A2(io_dmem_req_bits_cmd[0]), .Y(n5078) );
  NAND4X0_LVT U6479 ( .A1(ex_ctrl_mem), .A2(n5078), .A3(n3122), .A4(n3244), 
        .Y(n996) );
  AND3X1_LVT U6480 ( .A1(ex_ctrl_mem), .A2(n560), .A3(n3122), .Y(n5090) );
  OR2X1_LVT U6481 ( .A1(n559), .A2(io_dmem_req_bits_cmd[2]), .Y(n5079) );
  NAND3X0_LVT U6482 ( .A1(n5090), .A2(n3245), .A3(n5079), .Y(n882) );
  NAND2X0_LVT U6483 ( .A1(io_imem_bht_update_bits_branch), .A2(
        io_imem_bht_update_bits_taken), .Y(n5080) );
  AND2X1_LVT U6484 ( .A1(n555), .A2(n5080), .Y(n5084) );
  INVX1_LVT U6485 ( .A(n5080), .Y(n5085) );
  AND2X1_LVT U6486 ( .A1(n5085), .A2(n_T_844_10_), .Y(n5081) );
  AO21X1_LVT U6487 ( .A1(n5083), .A2(n_T_904[7]), .A3(n5081), .Y(n_T_914[19])
         );
  AO21X1_LVT U6488 ( .A1(n5083), .A2(n_T_904[6]), .A3(n5081), .Y(n_T_914[18])
         );
  AO21X1_LVT U6489 ( .A1(n5083), .A2(n_T_904[5]), .A3(n5081), .Y(n_T_914[17])
         );
  AO21X1_LVT U6490 ( .A1(n5083), .A2(n_T_904[4]), .A3(n5081), .Y(n_T_914[16])
         );
  AO21X1_LVT U6491 ( .A1(n5083), .A2(n_T_904[3]), .A3(n5081), .Y(n_T_914[15])
         );
  AO21X1_LVT U6492 ( .A1(n5083), .A2(n_T_904[2]), .A3(n5081), .Y(n_T_914[14])
         );
  AO21X1_LVT U6493 ( .A1(n5083), .A2(n_T_904[1]), .A3(n5081), .Y(n_T_914[13])
         );
  AO21X1_LVT U6494 ( .A1(n5083), .A2(n_T_904[0]), .A3(n5081), .Y(n_T_914[12])
         );
  AO22X1_LVT U6495 ( .A1(n5085), .A2(n_T_849[11]), .A3(n5083), .A4(n_T_911_11), 
        .Y(n_T_914[11]) );
  AND2X1_LVT U6496 ( .A1(n_T_849[10]), .A2(n5082), .Y(n_T_914[10]) );
  AND2X1_LVT U6497 ( .A1(n_T_849[9]), .A2(n5082), .Y(n_T_914[9]) );
  AND2X1_LVT U6498 ( .A1(n_T_849[8]), .A2(n5082), .Y(n_T_914[8]) );
  AND2X1_LVT U6499 ( .A1(n_T_849[7]), .A2(n5082), .Y(n_T_914[7]) );
  AND2X1_LVT U6500 ( .A1(n_T_849[6]), .A2(n5082), .Y(n_T_914[6]) );
  AND2X1_LVT U6501 ( .A1(n_T_849[5]), .A2(n5082), .Y(n_T_914[5]) );
  AO22X1_LVT U6502 ( .A1(n_T_911[4]), .A2(n5083), .A3(n5085), .A4(n_T_849[4]), 
        .Y(n_T_914[4]) );
  INVX1_LVT U6503 ( .A(io_fpu_inst[23]), .Y(n9441) );
  AO22X1_LVT U6504 ( .A1(n_T_911[3]), .A2(n5083), .A3(n5085), .A4(n2566), .Y(
        n_T_914[3]) );
  INVX1_LVT U6505 ( .A(io_fpu_inst[22]), .Y(n9442) );
  AO222X1_LVT U6506 ( .A1(n570), .A2(n5084), .A3(n_T_911[2]), .A4(n5083), .A5(
        n_T_849[2]), .A6(n5085), .Y(n_T_914[2]) );
  INVX1_LVT U6507 ( .A(io_fpu_inst[21]), .Y(n9443) );
  AO222X1_LVT U6508 ( .A1(n_T_849[1]), .A2(n5085), .A3(n5084), .A4(mem_reg_rvc), .A5(n5083), .A6(n_T_911[1]), .Y(n_T_914[1]) );
  NAND2X0_LVT U6509 ( .A1(mem_reg_valid), .A2(mem_reg_flush_pipe), .Y(n5091)
         );
  AND2X1_LVT U6510 ( .A1(n5089), .A2(n5091), .Y(N290) );
  AND2X1_LVT U6511 ( .A1(io_imem_req_bits_speculative), .A2(mem_reg_valid), 
        .Y(io_imem_bht_update_valid) );
  NAND2X0_LVT U6512 ( .A1(mem_ctrl_wxd), .A2(io_dmem_replay_next), .Y(n5404)
         );
  NAND2X0_LVT U6513 ( .A1(n2498), .A2(io_fpu_nack_mem), .Y(n5096) );
  AND2X1_LVT U6514 ( .A1(n5404), .A2(n5096), .Y(n5169) );
  NAND3X0_LVT U6515 ( .A1(n5102), .A2(n9075), .A3(n3578), .Y(n5103) );
  NAND2X0_LVT U6516 ( .A1(csr_io_decode_0_read_illegal), .A2(n5119), .Y(n5113)
         );
  NOR2X0_LVT U6517 ( .A1(io_fpu_illegal_rm), .A2(csr_io_decode_0_fp_illegal), 
        .Y(n5118) );
  OA21X1_LVT U6518 ( .A1(io_fpu_inst[28]), .A2(n5114), .A3(n9440), .Y(n5115)
         );
  NAND2X0_LVT U6519 ( .A1(csr_io_status_isa[0]), .A2(n5116), .Y(n5117) );
  OA21X1_LVT U6520 ( .A1(n5118), .A2(n1699), .A3(n5117), .Y(n5121) );
  OR2X1_LVT U6521 ( .A1(io_fpu_inst[18]), .A2(io_fpu_inst[17]), .Y(n5128) );
  OR2X1_LVT U6522 ( .A1(io_fpu_inst[15]), .A2(io_fpu_inst[16]), .Y(n5127) );
  OR3X1_LVT U6523 ( .A1(io_fpu_inst[10]), .A2(io_fpu_inst[19]), .A3(
        io_fpu_inst[11]), .Y(n5125) );
  OR3X1_LVT U6524 ( .A1(io_fpu_inst[8]), .A2(io_fpu_inst[9]), .A3(n5125), .Y(
        n5126) );
  OR3X1_LVT U6525 ( .A1(n5128), .A2(n5127), .A3(n5126), .Y(n5158) );
  INVX1_LVT U6526 ( .A(io_fpu_inst[24]), .Y(n5148) );
  NAND3X0_LVT U6527 ( .A1(n5132), .A2(n2565), .A3(n5131), .Y(n5141) );
  AND2X1_LVT U6528 ( .A1(io_fpu_inst[31]), .A2(n9445), .Y(n5136) );
  NAND4X0_LVT U6529 ( .A1(n5139), .A2(n3567), .A3(n5138), .A4(n5137), .Y(n5140) );
  OR3X1_LVT U6530 ( .A1(n5394), .A2(n5154), .A3(n5144), .Y(n5145) );
  NAND2X0_LVT U6531 ( .A1(n2537), .A2(n5146), .Y(n5147) );
  NAND2X0_LVT U6532 ( .A1(io_fpu_inst[22]), .A2(io_fpu_inst[21]), .Y(n5153) );
  OA21X1_LVT U6533 ( .A1(io_fpu_inst[22]), .A2(n9444), .A3(n5153), .Y(n5157)
         );
  NAND2X0_LVT U6534 ( .A1(n5154), .A2(n3079), .Y(n5155) );
  NAND3X0_LVT U6535 ( .A1(n5157), .A2(n5156), .A3(n5155), .Y(n5159) );
  OR3X1_LVT U6536 ( .A1(n5160), .A2(n5159), .A3(n5158), .Y(n5161) );
  NAND2X0_LVT U6537 ( .A1(n9430), .A2(n9118), .Y(n9243) );
  AND3X1_LVT U6538 ( .A1(n9418), .A2(ex_reg_valid), .A3(n9421), .Y(n407) );
  INVX1_LVT U6539 ( .A(n407), .Y(io_fpu_killx) );
  OR3X1_LVT U6540 ( .A1(mem_reg_sfence), .A2(csr_io_status_isa[2]), .A3(n9512), 
        .Y(n5405) );
  INVX1_LVT U6541 ( .A(n1279), .Y(n5168) );
  OA21X1_LVT U6542 ( .A1(n3206), .A2(n5405), .A3(n5168), .Y(n9425) );
  NAND3X0_LVT U6543 ( .A1(io_imem_bht_update_valid), .A2(n5169), .A3(n3251), 
        .Y(n5171) );
  AO22X1_LVT U6544 ( .A1(mem_reg_store), .A2(bpu_io_xcpt_st), .A3(
        bpu_io_xcpt_ld), .A4(mem_reg_load), .Y(n5170) );
  AO22X1_LVT U6545 ( .A1(mem_reg_store), .A2(bpu_io_debug_st), .A3(
        bpu_io_debug_ld), .A4(mem_reg_load), .Y(n9237) );
  OR2X1_LVT U6546 ( .A1(n5170), .A2(n9237), .Y(n5172) );
  OR2X1_LVT U6547 ( .A1(n5171), .A2(n5172), .Y(io_dmem_s1_kill) );
  NOR2X0_LVT U6548 ( .A1(n1281), .A2(io_dmem_s1_kill), .Y(n1829) );
  AO22X1_LVT U6549 ( .A1(io_imem_req_bits_speculative), .A2(n1281), .A3(n5172), 
        .A4(io_imem_bht_update_valid), .Y(N529) );
  AND2X1_LVT U6550 ( .A1(n3198), .A2(n3043), .Y(n5227) );
  AND2X1_LVT U6551 ( .A1(n5227), .A2(n3199), .Y(n5354) );
  AND2X1_LVT U6552 ( .A1(n3103), .A2(n3041), .Y(n5272) );
  AO21X1_LVT U6553 ( .A1(n5175), .A2(wb_ctrl_wfd), .A3(io_fpu_sboard_set), .Y(
        n5176) );
  AO21X1_LVT U6554 ( .A1(n5354), .A2(n5275), .A3(n_T_1298[5]), .Y(n5179) );
  AND3X1_LVT U6555 ( .A1(io_dmem_resp_bits_has_data), .A2(
        io_dmem_resp_bits_tag[0]), .A3(n2030), .Y(io_fpu_dmem_resp_val) );
  NAND2X0_LVT U6556 ( .A1(io_fpu_dmem_resp_val), .A2(io_dmem_resp_bits_replay), 
        .Y(n5191) );
  NAND3X0_LVT U6557 ( .A1(n5254), .A2(n5191), .A3(n5177), .Y(n9379) );
  NAND2X0_LVT U6558 ( .A1(n5183), .A2(io_fpu_sboard_clra[0]), .Y(n5271) );
  OR2X1_LVT U6559 ( .A1(n5257), .A2(n5271), .Y(n5277) );
  OA22X1_LVT U6560 ( .A1(n5277), .A2(n5193), .A3(n5192), .A4(n5276), .Y(n5178)
         );
  AND3X1_LVT U6561 ( .A1(n5179), .A2(n3794), .A3(n5178), .Y(N784) );
  AND2X1_LVT U6562 ( .A1(n3199), .A2(n3102), .Y(n5255) );
  AND2X1_LVT U6563 ( .A1(n5255), .A2(n3198), .Y(n5355) );
  AND2X1_LVT U6564 ( .A1(n3201), .A2(wb_waddr[1]), .Y(n5303) );
  AO21X1_LVT U6565 ( .A1(n5355), .A2(n5248), .A3(n_T_1298[2]), .Y(n5181) );
  AND2X1_LVT U6566 ( .A1(io_fpu_sboard_clr), .A2(io_fpu_sboard_clra[1]), .Y(
        n5190) );
  NAND2X0_LVT U6567 ( .A1(n5190), .A2(n5182), .Y(n5262) );
  OR2X1_LVT U6568 ( .A1(io_fpu_sboard_clra[2]), .A2(n5193), .Y(n5201) );
  OR2X1_LVT U6569 ( .A1(io_fpu_dmem_resp_tag[2]), .A2(n5192), .Y(n5200) );
  OA22X1_LVT U6570 ( .A1(n5262), .A2(n5201), .A3(n5200), .A4(n5261), .Y(n5180)
         );
  AND3X1_LVT U6571 ( .A1(n5181), .A2(n3793), .A3(n5180), .Y(N781) );
  AND2X1_LVT U6572 ( .A1(n3103), .A2(n3201), .Y(n5282) );
  AO21X1_LVT U6573 ( .A1(n5354), .A2(n5265), .A3(n_T_1298[4]), .Y(n5187) );
  NAND2X0_LVT U6574 ( .A1(n5183), .A2(n5182), .Y(n5281) );
  OR2X1_LVT U6575 ( .A1(n5257), .A2(n5281), .Y(n5267) );
  OA22X1_LVT U6576 ( .A1(n5193), .A2(n5267), .A3(n5192), .A4(n5266), .Y(n5186)
         );
  AND3X1_LVT U6577 ( .A1(n5187), .A2(n3793), .A3(n5186), .Y(N783) );
  AO21X1_LVT U6578 ( .A1(n5354), .A2(n5248), .A3(n_T_1298[6]), .Y(n5189) );
  OR2X1_LVT U6579 ( .A1(n5257), .A2(n5262), .Y(n5251) );
  OR2X1_LVT U6580 ( .A1(n5259), .A2(n5261), .Y(n5250) );
  OA22X1_LVT U6581 ( .A1(n5193), .A2(n5251), .A3(n5192), .A4(n5250), .Y(n5188)
         );
  AND3X1_LVT U6582 ( .A1(n5189), .A2(n3794), .A3(n5188), .Y(N785) );
  AND2X1_LVT U6583 ( .A1(n3041), .A2(wb_waddr[1]), .Y(n5298) );
  AO21X1_LVT U6584 ( .A1(n5354), .A2(n5285), .A3(n_T_1298[7]), .Y(n5195) );
  NAND2X0_LVT U6585 ( .A1(n5190), .A2(io_fpu_sboard_clra[0]), .Y(n5295) );
  OR2X1_LVT U6586 ( .A1(n5257), .A2(n5295), .Y(n5288) );
  OR2X1_LVT U6587 ( .A1(n5259), .A2(n5292), .Y(n5286) );
  OA22X1_LVT U6588 ( .A1(n5193), .A2(n5288), .A3(n5192), .A4(n5286), .Y(n5194)
         );
  AND3X1_LVT U6589 ( .A1(n5195), .A2(n3793), .A3(n5194), .Y(N786) );
  AO21X1_LVT U6590 ( .A1(n5355), .A2(n5275), .A3(n_T_1298[1]), .Y(n5197) );
  OA22X1_LVT U6591 ( .A1(n5271), .A2(n5201), .A3(n5200), .A4(n5270), .Y(n5196)
         );
  AND3X1_LVT U6592 ( .A1(n5197), .A2(n3793), .A3(n5196), .Y(N780) );
  AO21X1_LVT U6593 ( .A1(n5355), .A2(n5265), .A3(n_T_1298[0]), .Y(n5199) );
  OA22X1_LVT U6594 ( .A1(n5281), .A2(n5201), .A3(n5200), .A4(n5280), .Y(n5198)
         );
  AND3X1_LVT U6595 ( .A1(n5199), .A2(n3794), .A3(n5198), .Y(N779) );
  AO21X1_LVT U6596 ( .A1(n5355), .A2(n5285), .A3(n_T_1298[3]), .Y(n5203) );
  OA22X1_LVT U6597 ( .A1(n5295), .A2(n5201), .A3(n5200), .A4(n5292), .Y(n5202)
         );
  AND3X1_LVT U6598 ( .A1(n5203), .A2(n3794), .A3(n5202), .Y(N782) );
  AND2X1_LVT U6599 ( .A1(wb_waddr[4]), .A2(wb_waddr[3]), .Y(n5210) );
  AND2X1_LVT U6600 ( .A1(n5210), .A2(n3102), .Y(n5305) );
  AO21X1_LVT U6601 ( .A1(n5305), .A2(n5248), .A3(n_T_1298[26]), .Y(n5205) );
  AND2X1_LVT U6602 ( .A1(io_fpu_sboard_clra[3]), .A2(io_fpu_sboard_clra[4]), 
        .Y(n5211) );
  NAND2X0_LVT U6603 ( .A1(n5211), .A2(n5257), .Y(n5218) );
  AND2X1_LVT U6604 ( .A1(io_fpu_dmem_resp_tag[3]), .A2(io_fpu_dmem_resp_tag[4]), .Y(n5212) );
  NAND2X0_LVT U6605 ( .A1(n5212), .A2(n5259), .Y(n5217) );
  OA22X1_LVT U6606 ( .A1(n5262), .A2(n5218), .A3(n5217), .A4(n5261), .Y(n5204)
         );
  AND3X1_LVT U6607 ( .A1(n5205), .A2(n3794), .A3(n5204), .Y(N805) );
  AO21X1_LVT U6608 ( .A1(n5305), .A2(n5275), .A3(n_T_1298[25]), .Y(n5207) );
  OA22X1_LVT U6609 ( .A1(n5271), .A2(n5218), .A3(n5217), .A4(n5270), .Y(n5206)
         );
  AND3X1_LVT U6610 ( .A1(n5207), .A2(n3794), .A3(n5206), .Y(N804) );
  AO21X1_LVT U6611 ( .A1(n5305), .A2(n5285), .A3(n_T_1298[27]), .Y(n5209) );
  OA22X1_LVT U6612 ( .A1(n5295), .A2(n5218), .A3(n5217), .A4(n5292), .Y(n5208)
         );
  AND3X1_LVT U6613 ( .A1(n5209), .A2(n3794), .A3(n5208), .Y(N806) );
  AO21X1_LVT U6614 ( .A1(n5317), .A2(n5248), .A3(n_T_1298[30]), .Y(n5214) );
  INVX1_LVT U6615 ( .A(n5211), .Y(n5224) );
  INVX1_LVT U6616 ( .A(n5212), .Y(n5223) );
  OA22X1_LVT U6617 ( .A1(n5251), .A2(n5224), .A3(n5223), .A4(n5250), .Y(n5213)
         );
  AND3X1_LVT U6618 ( .A1(n5214), .A2(n3794), .A3(n5213), .Y(N809) );
  AO21X1_LVT U6619 ( .A1(n5317), .A2(n5275), .A3(n_T_1298[29]), .Y(n5216) );
  OA22X1_LVT U6620 ( .A1(n5277), .A2(n5224), .A3(n5223), .A4(n5276), .Y(n5215)
         );
  AND3X1_LVT U6621 ( .A1(n5216), .A2(n3794), .A3(n5215), .Y(N808) );
  AO21X1_LVT U6622 ( .A1(n5305), .A2(n5265), .A3(n_T_1298[24]), .Y(n5220) );
  OA22X1_LVT U6623 ( .A1(n5281), .A2(n5218), .A3(n5217), .A4(n5280), .Y(n5219)
         );
  AND3X1_LVT U6624 ( .A1(n5220), .A2(n3794), .A3(n5219), .Y(N803) );
  AO21X1_LVT U6625 ( .A1(n5317), .A2(n5265), .A3(n_T_1298[28]), .Y(n5222) );
  OA22X1_LVT U6626 ( .A1(n5267), .A2(n5224), .A3(n5223), .A4(n5266), .Y(n5221)
         );
  AND3X1_LVT U6627 ( .A1(n5222), .A2(n3794), .A3(n5221), .Y(N807) );
  AO21X1_LVT U6628 ( .A1(n5317), .A2(n5285), .A3(n_T_1298[31]), .Y(n5226) );
  OA22X1_LVT U6629 ( .A1(n5288), .A2(n5224), .A3(n5223), .A4(n5286), .Y(n5225)
         );
  AND3X1_LVT U6630 ( .A1(n5226), .A2(n3794), .A3(n5225), .Y(N810) );
  AO21X1_LVT U6631 ( .A1(n5382), .A2(n5285), .A3(n_T_1298[15]), .Y(n5230) );
  NAND2X0_LVT U6632 ( .A1(n5228), .A2(io_fpu_dmem_resp_tag[3]), .Y(n5244) );
  OA22X1_LVT U6633 ( .A1(n5245), .A2(n5288), .A3(n5244), .A4(n5286), .Y(n5229)
         );
  AND3X1_LVT U6634 ( .A1(n5230), .A2(n3794), .A3(n5229), .Y(N794) );
  AO21X1_LVT U6635 ( .A1(n5382), .A2(n5248), .A3(n_T_1298[14]), .Y(n5232) );
  OA22X1_LVT U6636 ( .A1(n5245), .A2(n5251), .A3(n5244), .A4(n5250), .Y(n5231)
         );
  AND3X1_LVT U6637 ( .A1(n5232), .A2(n3794), .A3(n5231), .Y(N793) );
  OR2X1_LVT U6638 ( .A1(io_fpu_sboard_clra[2]), .A2(n5245), .Y(n5238) );
  NAND3X0_LVT U6639 ( .A1(n3198), .A2(n3102), .A3(wb_waddr[3]), .Y(n5359) );
  NOR3X0_LVT U6640 ( .A1(reset), .A2(n5359), .A3(n5254), .Y(n5239) );
  OA22X1_LVT U6641 ( .A1(n5238), .A2(n5262), .A3(n5237), .A4(n5261), .Y(n5234)
         );
  AO22X1_LVT U6642 ( .A1(n5239), .A2(n5303), .A3(n_T_1298[10]), .A4(n3793), 
        .Y(n5233) );
  AND2X1_LVT U6643 ( .A1(n5234), .A2(n5233), .Y(N789) );
  OA22X1_LVT U6644 ( .A1(n5238), .A2(n5281), .A3(n5237), .A4(n5280), .Y(n5236)
         );
  AO22X1_LVT U6645 ( .A1(n5239), .A2(n5282), .A3(n_T_1298[8]), .A4(n3793), .Y(
        n5235) );
  AND2X1_LVT U6646 ( .A1(n5236), .A2(n5235), .Y(N787) );
  OA22X1_LVT U6647 ( .A1(n5238), .A2(n5271), .A3(n5237), .A4(n5270), .Y(n5241)
         );
  AO22X1_LVT U6648 ( .A1(n5239), .A2(n5272), .A3(n_T_1298[9]), .A4(n3793), .Y(
        n5240) );
  AND2X1_LVT U6649 ( .A1(n5241), .A2(n5240), .Y(N788) );
  AO21X1_LVT U6650 ( .A1(n5382), .A2(n5265), .A3(n_T_1298[12]), .Y(n5243) );
  OA22X1_LVT U6651 ( .A1(n5245), .A2(n5267), .A3(n5244), .A4(n5266), .Y(n5242)
         );
  AND3X1_LVT U6652 ( .A1(n5243), .A2(n5296), .A3(n5242), .Y(N791) );
  AO21X1_LVT U6653 ( .A1(n5382), .A2(n5275), .A3(n_T_1298[13]), .Y(n5247) );
  OA22X1_LVT U6654 ( .A1(n5245), .A2(n5277), .A3(n5244), .A4(n5276), .Y(n5246)
         );
  AND3X1_LVT U6655 ( .A1(n5247), .A2(n5296), .A3(n5246), .Y(N792) );
  AND3X1_LVT U6656 ( .A1(n3199), .A2(n3043), .A3(wb_waddr[4]), .Y(n5325) );
  AO21X1_LVT U6657 ( .A1(n5325), .A2(n5248), .A3(n_T_1298[22]), .Y(n5253) );
  INVX1_LVT U6658 ( .A(n5258), .Y(n5289) );
  AND2X1_LVT U6659 ( .A1(n5249), .A2(io_fpu_dmem_resp_tag[4]), .Y(n5260) );
  OA22X1_LVT U6660 ( .A1(n5289), .A2(n5251), .A3(n5287), .A4(n5250), .Y(n5252)
         );
  AND3X1_LVT U6661 ( .A1(n5253), .A2(n5296), .A3(n5252), .Y(N801) );
  AND2X1_LVT U6662 ( .A1(n5255), .A2(wb_waddr[4]), .Y(n5326) );
  AND3X1_LVT U6663 ( .A1(n5256), .A2(n5326), .A3(n4498), .Y(n5297) );
  AO22X1_LVT U6664 ( .A1(n5303), .A2(n5297), .A3(n3793), .A4(n_T_1298[18]), 
        .Y(n5264) );
  NAND2X0_LVT U6665 ( .A1(n5258), .A2(n5257), .Y(n5294) );
  NAND2X0_LVT U6666 ( .A1(n5260), .A2(n5259), .Y(n5293) );
  OA22X1_LVT U6667 ( .A1(n5262), .A2(n5294), .A3(n5293), .A4(n5261), .Y(n5263)
         );
  AND2X1_LVT U6668 ( .A1(n5264), .A2(n5263), .Y(N797) );
  AO21X1_LVT U6669 ( .A1(n5325), .A2(n5265), .A3(n_T_1298[20]), .Y(n5269) );
  OA22X1_LVT U6670 ( .A1(n5289), .A2(n5267), .A3(n5287), .A4(n5266), .Y(n5268)
         );
  AND3X1_LVT U6671 ( .A1(n5269), .A2(n5296), .A3(n5268), .Y(N799) );
  OA22X1_LVT U6672 ( .A1(n5271), .A2(n5294), .A3(n5293), .A4(n5270), .Y(n5274)
         );
  AO22X1_LVT U6673 ( .A1(n5272), .A2(n5297), .A3(n3793), .A4(n_T_1298[17]), 
        .Y(n5273) );
  AND2X1_LVT U6674 ( .A1(n5274), .A2(n5273), .Y(N796) );
  AO21X1_LVT U6675 ( .A1(n5325), .A2(n5275), .A3(n_T_1298[21]), .Y(n5279) );
  OA22X1_LVT U6676 ( .A1(n5289), .A2(n5277), .A3(n5287), .A4(n5276), .Y(n5278)
         );
  AND3X1_LVT U6677 ( .A1(n5279), .A2(n5296), .A3(n5278), .Y(N800) );
  OA22X1_LVT U6678 ( .A1(n5281), .A2(n5294), .A3(n5293), .A4(n5280), .Y(n5284)
         );
  AO22X1_LVT U6679 ( .A1(n5282), .A2(n5297), .A3(n3793), .A4(n_T_1298[16]), 
        .Y(n5283) );
  AND2X1_LVT U6680 ( .A1(n5284), .A2(n5283), .Y(N795) );
  AO21X1_LVT U6681 ( .A1(n5325), .A2(n5285), .A3(n_T_1298[23]), .Y(n5291) );
  OA22X1_LVT U6682 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .Y(n5290)
         );
  AND3X1_LVT U6683 ( .A1(n5291), .A2(n3793), .A3(n5290), .Y(N802) );
  OA22X1_LVT U6684 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .Y(n5300)
         );
  AO22X1_LVT U6685 ( .A1(n5298), .A2(n5297), .A3(n3793), .A4(n_T_1298[19]), 
        .Y(n5299) );
  AND2X1_LVT U6686 ( .A1(n5300), .A2(n5299), .Y(N798) );
  AND2X1_LVT U6687 ( .A1(n5301), .A2(csr_io_retire), .Y(n9380) );
  NAND2X0_LVT U6688 ( .A1(n3046), .A2(n4498), .Y(n5302) );
  AND2X1_LVT U6689 ( .A1(n5304), .A2(n5303), .Y(n5374) );
  NAND2X0_LVT U6690 ( .A1(n5378), .A2(n5305), .Y(n5310) );
  NAND2X0_LVT U6691 ( .A1(n5307), .A2(n5335), .Y(n5308) );
  NAND3X0_LVT U6692 ( .A1(n5308), .A2(n2572), .A3(n_T_1187[27]), .Y(n5309) );
  AND2X1_LVT U6693 ( .A1(n5379), .A2(n5313), .Y(n5367) );
  AND2X1_LVT U6694 ( .A1(n5339), .A2(n3046), .Y(n5363) );
  AND2X1_LVT U6695 ( .A1(n5313), .A2(n5363), .Y(n5385) );
  AND2X1_LVT U6696 ( .A1(n_T_1187[30]), .A2(n2572), .Y(n5312) );
  AND2X1_LVT U6697 ( .A1(n5356), .A2(n3046), .Y(n5390) );
  AND2X1_LVT U6698 ( .A1(n5313), .A2(n5390), .Y(n5371) );
  NAND2X0_LVT U6699 ( .A1(n5371), .A2(n5314), .Y(n5311) );
  AO22X1_LVT U6700 ( .A1(n5317), .A2(n5374), .A3(n5312), .A4(n5311), .Y(N776)
         );
  AND2X1_LVT U6701 ( .A1(n_T_1187[31]), .A2(n2572), .Y(n5316) );
  AND2X1_LVT U6702 ( .A1(n5335), .A2(n3046), .Y(n5360) );
  AND2X1_LVT U6703 ( .A1(n5360), .A2(n5313), .Y(n5375) );
  NAND2X0_LVT U6704 ( .A1(n5375), .A2(n5314), .Y(n5315) );
  AO22X1_LVT U6705 ( .A1(n5378), .A2(n5317), .A3(n5316), .A4(n5315), .Y(N777)
         );
  NAND2X0_LVT U6706 ( .A1(n5366), .A2(n5325), .Y(n5320) );
  NAND2X0_LVT U6707 ( .A1(n5367), .A2(n5328), .Y(n5318) );
  NAND3X0_LVT U6708 ( .A1(n5318), .A2(n_T_1187[20]), .A3(n2572), .Y(n5319) );
  NAND2X0_LVT U6709 ( .A1(n5320), .A2(n5319), .Y(N766) );
  AND2X1_LVT U6710 ( .A1(n_T_1187[22]), .A2(n2572), .Y(n5322) );
  NAND2X0_LVT U6711 ( .A1(n5371), .A2(n5328), .Y(n5321) );
  AO22X1_LVT U6712 ( .A1(n5325), .A2(n5374), .A3(n5322), .A4(n5321), .Y(N768)
         );
  AND2X1_LVT U6713 ( .A1(n_T_1187[23]), .A2(n2572), .Y(n5324) );
  NAND2X0_LVT U6714 ( .A1(n5375), .A2(n5328), .Y(n5323) );
  AO22X1_LVT U6715 ( .A1(n5378), .A2(n5325), .A3(n5324), .A4(n5323), .Y(N769)
         );
  AND2X1_LVT U6716 ( .A1(n5328), .A2(n2575), .Y(n5332) );
  AO21X1_LVT U6717 ( .A1(n5360), .A2(n5332), .A3(n3258), .Y(n5329) );
  OAI22X1_LVT U6718 ( .A1(n5334), .A2(n5362), .A3(n5329), .A4(n3185), .Y(N765)
         );
  AO21X1_LVT U6719 ( .A1(n5363), .A2(n5332), .A3(n3113), .Y(n5330) );
  OAI22X1_LVT U6720 ( .A1(n5334), .A2(n5365), .A3(n5330), .A4(n3185), .Y(N763)
         );
  AO21X1_LVT U6721 ( .A1(n5379), .A2(n5332), .A3(n3261), .Y(n5331) );
  OAI22X1_LVT U6722 ( .A1(n5381), .A2(n5334), .A3(n5331), .A4(n3185), .Y(N762)
         );
  AO21X1_LVT U6723 ( .A1(n5390), .A2(n5332), .A3(n3263), .Y(n5333) );
  OAI22X1_LVT U6724 ( .A1(n5334), .A2(n5392), .A3(n5333), .A4(n3185), .Y(N764)
         );
  NAND2X0_LVT U6725 ( .A1(n5378), .A2(n5355), .Y(n5338) );
  AND2X1_LVT U6726 ( .A1(n5426), .A2(n5428), .Y(n5351) );
  NAND2X0_LVT U6727 ( .A1(n5357), .A2(n5335), .Y(n5336) );
  NAND3X0_LVT U6728 ( .A1(n2572), .A2(n_T_1187[3]), .A3(n5336), .Y(n5337) );
  NAND2X0_LVT U6729 ( .A1(n5338), .A2(n5337), .Y(N749) );
  NAND2X0_LVT U6730 ( .A1(n5383), .A2(n5355), .Y(n5342) );
  NAND2X0_LVT U6731 ( .A1(n5357), .A2(n5339), .Y(n5340) );
  NAND3X0_LVT U6732 ( .A1(n2572), .A2(n_T_1187[1]), .A3(n5340), .Y(n5341) );
  NAND2X0_LVT U6733 ( .A1(n5342), .A2(n5341), .Y(N747) );
  NAND2X0_LVT U6734 ( .A1(n5383), .A2(n5354), .Y(n5345) );
  NAND2X0_LVT U6735 ( .A1(n5385), .A2(n5351), .Y(n5343) );
  NAND3X0_LVT U6736 ( .A1(n5343), .A2(n_T_1187[5]), .A3(n2572), .Y(n5344) );
  NAND2X0_LVT U6737 ( .A1(n5345), .A2(n5344), .Y(N751) );
  AND2X1_LVT U6738 ( .A1(n_T_1187[6]), .A2(n2572), .Y(n5347) );
  NAND2X0_LVT U6739 ( .A1(n5371), .A2(n5351), .Y(n5346) );
  AO22X1_LVT U6740 ( .A1(n5354), .A2(n5374), .A3(n5347), .A4(n5346), .Y(N752)
         );
  NAND2X0_LVT U6741 ( .A1(n5366), .A2(n5354), .Y(n5350) );
  NAND2X0_LVT U6742 ( .A1(n5367), .A2(n5351), .Y(n5348) );
  NAND3X0_LVT U6743 ( .A1(n5348), .A2(n_T_1187[4]), .A3(n2572), .Y(n5349) );
  NAND2X0_LVT U6744 ( .A1(n5350), .A2(n5349), .Y(N750) );
  AND2X1_LVT U6745 ( .A1(n_T_1187[7]), .A2(n2572), .Y(n5353) );
  NAND2X0_LVT U6746 ( .A1(n5375), .A2(n5351), .Y(n5352) );
  AO22X1_LVT U6747 ( .A1(n5378), .A2(n5354), .A3(n5353), .A4(n5352), .Y(N753)
         );
  AND2X1_LVT U6748 ( .A1(n5384), .A2(n2575), .Y(n5389) );
  AO21X1_LVT U6749 ( .A1(n5360), .A2(n5389), .A3(n3259), .Y(n5361) );
  OAI22X1_LVT U6750 ( .A1(n5393), .A2(n5362), .A3(n5361), .A4(n3185), .Y(N757)
         );
  AO21X1_LVT U6751 ( .A1(n5363), .A2(n5389), .A3(n3133), .Y(n5364) );
  OAI22X1_LVT U6752 ( .A1(n5393), .A2(n5365), .A3(n5364), .A4(n3185), .Y(N755)
         );
  NAND2X0_LVT U6753 ( .A1(n5366), .A2(n5382), .Y(n5370) );
  NAND2X0_LVT U6754 ( .A1(n5367), .A2(n5384), .Y(n5368) );
  NAND3X0_LVT U6755 ( .A1(n5368), .A2(n_T_1187[12]), .A3(n2572), .Y(n5369) );
  NAND2X0_LVT U6756 ( .A1(n5370), .A2(n5369), .Y(N758) );
  AND2X1_LVT U6757 ( .A1(n_T_1187[14]), .A2(n2572), .Y(n5373) );
  NAND2X0_LVT U6758 ( .A1(n5371), .A2(n5384), .Y(n5372) );
  AO22X1_LVT U6759 ( .A1(n5382), .A2(n5374), .A3(n5373), .A4(n5372), .Y(N760)
         );
  AND2X1_LVT U6760 ( .A1(n_T_1187[15]), .A2(n2572), .Y(n5377) );
  NAND2X0_LVT U6761 ( .A1(n5375), .A2(n5384), .Y(n5376) );
  AO22X1_LVT U6762 ( .A1(n5378), .A2(n5382), .A3(n5377), .A4(n5376), .Y(N761)
         );
  AO21X1_LVT U6763 ( .A1(n5379), .A2(n5389), .A3(n3134), .Y(n5380) );
  OAI22X1_LVT U6764 ( .A1(n5381), .A2(n5393), .A3(n5380), .A4(n3185), .Y(N754)
         );
  NAND2X0_LVT U6765 ( .A1(n5383), .A2(n5382), .Y(n5388) );
  NAND2X0_LVT U6766 ( .A1(n5385), .A2(n5384), .Y(n5386) );
  NAND3X0_LVT U6767 ( .A1(n5386), .A2(n_T_1187[13]), .A3(n2572), .Y(n5387) );
  NAND2X0_LVT U6768 ( .A1(n5388), .A2(n5387), .Y(N759) );
  AO21X1_LVT U6769 ( .A1(n5390), .A2(n5389), .A3(n3129), .Y(n5391) );
  OAI22X1_LVT U6770 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n3185), .Y(N756)
         );
  NOR3X0_LVT U6771 ( .A1(io_fpu_inst[23]), .A2(n5394), .A3(io_fpu_inst[22]), 
        .Y(n5395) );
  INVX1_LVT U6772 ( .A(io_dmem_perf_release), .Y(n5399) );
  OR3X1_LVT U6773 ( .A1(csr_io_time[0]), .A2(csr_io_time[4]), .A3(
        csr_io_time[3]), .Y(n5397) );
  OR3X1_LVT U6774 ( .A1(csr_io_time[1]), .A2(csr_io_time[2]), .A3(n5397), .Y(
        n5398) );
  AND3X1_LVT U6775 ( .A1(n9418), .A2(n5399), .A3(n5398), .Y(n5400) );
  OA21X1_LVT U6776 ( .A1(id_reg_pause), .A2(n5401), .A3(n5400), .Y(n1820) );
  NAND3X0_LVT U6777 ( .A1(io_imem_bht_update_valid), .A2(n3251), .A3(n5404), 
        .Y(io_fpu_killm) );
  AND2X1_LVT U6778 ( .A1(io_fpu_killm), .A2(n_T_1057), .Y(div_io_kill) );
  NAND2X0_LVT U6779 ( .A1(n5419), .A2(n5421), .Y(n5480) );
  OR2X1_LVT U6780 ( .A1(n5420), .A2(n5480), .Y(do_bypass_1) );
  INVX1_LVT U6781 ( .A(n5409), .Y(n5407) );
  AND2X1_LVT U6782 ( .A1(mem_ctrl_wxd), .A2(n2492), .Y(n5408) );
  AO222X1_LVT U6783 ( .A1(n6249), .A2(io_imem_btb_update_bits_br_pc[0]), .A3(
        n6855), .A4(n_T_918[0]), .A5(io_fpu_toint_data[0]), .A6(n6856), .Y(
        N598) );
  AND2X1_LVT U6784 ( .A1(n5414), .A2(n5413), .Y(n5416) );
  AO22X1_LVT U6785 ( .A1(n6860), .A2(io_dmem_resp_bits_data[0]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[0]), .Y(n5417) );
  AO21X1_LVT U6786 ( .A1(n3854), .A2(div_io_resp_bits_data[0]), .A3(n5417), 
        .Y(n5418) );
  AO21X1_LVT U6787 ( .A1(n3841), .A2(csr_io_rw_rdata[0]), .A3(n5418), .Y(
        n_T_427__T_1136_data[0]) );
  NAND3X0_LVT U6788 ( .A1(n5420), .A2(n572), .A3(n5419), .Y(n5422) );
  AND2X1_LVT U6789 ( .A1(n5422), .A2(n5421), .Y(n5468) );
  AND2X1_LVT U6790 ( .A1(n5425), .A2(n5424), .Y(n5433) );
  NAND2X0_LVT U6791 ( .A1(n9398), .A2(n9403), .Y(n9386) );
  AND2X1_LVT U6792 ( .A1(n5429), .A2(n9388), .Y(n5430) );
  AND2X1_LVT U6793 ( .A1(n5451), .A2(n2878), .Y(n6795) );
  AND2X1_LVT U6794 ( .A1(n5456), .A2(n2878), .Y(n6869) );
  AND2X1_LVT U6795 ( .A1(n5454), .A2(n2878), .Y(n6715) );
  AO22X1_LVT U6796 ( .A1(n3811), .A2(n_T_427[895]), .A3(n_T_427[640]), .A4(
        n3861), .Y(n5442) );
  AO22X1_LVT U6797 ( .A1(n_T_427[704]), .A2(n3804), .A3(n3860), .A4(
        n_T_427[192]), .Y(n5441) );
  AO22X1_LVT U6798 ( .A1(n_T_427[831]), .A2(n6871), .A3(n3872), .A4(
        n_T_427[256]), .Y(n5440) );
  AO22X1_LVT U6799 ( .A1(n3815), .A2(n_T_427[128]), .A3(n3839), .A4(n_T_427[0]), .Y(n5439) );
  NOR4X1_LVT U6800 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .Y(n5443)
         );
  NAND2X0_LVT U6801 ( .A1(n4318), .A2(n3959), .Y(n5444) );
  AND2X1_LVT U6802 ( .A1(n5446), .A2(n5456), .Y(n6880) );
  AND2X1_LVT U6803 ( .A1(n5446), .A2(n5455), .Y(n6891) );
  INVX1_LVT U6804 ( .A(n5447), .Y(n5448) );
  AND2X1_LVT U6805 ( .A1(n5457), .A2(n5450), .Y(n6893) );
  AO22X1_LVT U6806 ( .A1(n3934), .A2(n_T_427[1407]), .A3(n_T_427[1279]), .A4(
        n3929), .Y(n5461) );
  AND2X1_LVT U6807 ( .A1(n5457), .A2(n5452), .Y(n6895) );
  AO22X1_LVT U6808 ( .A1(n3944), .A2(n_T_427[1151]), .A3(n_T_427[1215]), .A4(
        n3939), .Y(n5460) );
  AND2X1_LVT U6809 ( .A1(n5457), .A2(n5454), .Y(n6897) );
  AO22X1_LVT U6810 ( .A1(n3954), .A2(n_T_427[1087]), .A3(n_T_427[959]), .A4(
        n3949), .Y(n5459) );
  AND2X1_LVT U6811 ( .A1(n5457), .A2(n5456), .Y(n6883) );
  AO22X1_LVT U6812 ( .A1(n3900), .A2(n_T_427[1023]), .A3(n_T_427[64]), .A4(
        n3831), .Y(n5458) );
  NOR4X1_LVT U6813 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .Y(n5462)
         );
  NAND3X0_LVT U6814 ( .A1(n5462), .A2(n5463), .A3(n5464), .Y(n5467) );
  INVX1_LVT U6815 ( .A(do_bypass_1), .Y(n5465) );
  AND2X1_LVT U6816 ( .A1(n5466), .A2(n5465), .Y(n9382) );
  MUX21X1_LVT U6817 ( .A1(n5468), .A2(n5467), .S0(n9382), .Y(N678) );
  AO222X1_LVT U6818 ( .A1(mem_br_target_1_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[1]), .A5(n_T_918[1]), .A6(n6855), .Y(N599) );
  NAND2X0_LVT U6819 ( .A1(csr_io_rw_rdata[1]), .A2(n3844), .Y(n5471) );
  AOI22X1_LVT U6820 ( .A1(n3852), .A2(io_dmem_resp_bits_data[1]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[1]), .Y(n5470) );
  NAND2X0_LVT U6821 ( .A1(div_io_resp_bits_data[1]), .A2(n3857), .Y(n5469) );
  NAND3X0_LVT U6822 ( .A1(n5471), .A2(n5470), .A3(n5469), .Y(
        n_T_427__T_1136_data[1]) );
  AO22X1_LVT U6823 ( .A1(n_T_427[896]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[449]), .Y(n5478) );
  AO22X1_LVT U6824 ( .A1(n3815), .A2(n_T_427[129]), .A3(n3871), .A4(
        n_T_427[257]), .Y(n5477) );
  AOI22X1_LVT U6825 ( .A1(n3797), .A2(n_T_427[577]), .A3(n3867), .A4(
        n_T_427[321]), .Y(n5475) );
  AOI22X1_LVT U6826 ( .A1(n6765), .A2(n_T_427[705]), .A3(n3859), .A4(
        n_T_427[193]), .Y(n5474) );
  AOI22X1_LVT U6827 ( .A1(n_T_427[641]), .A2(n3861), .A3(n3868), .A4(
        n_T_427[513]), .Y(n5473) );
  NAND2X0_LVT U6828 ( .A1(n3840), .A2(n_T_427[1]), .Y(n5472) );
  NAND4X0_LVT U6829 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .Y(n5476) );
  OR3X1_LVT U6830 ( .A1(n5478), .A2(n5477), .A3(n5476), .Y(n5479) );
  NAND2X0_LVT U6831 ( .A1(n_T_918[0]), .A2(n6899), .Y(n9125) );
  AND2X1_LVT U6832 ( .A1(n594), .A2(n_T_635[1]), .Y(n5484) );
  NAND2X0_LVT U6833 ( .A1(io_imem_sfence_bits_addr[0]), .A2(n6900), .Y(n9124)
         );
  OR2X1_LVT U6834 ( .A1(ex_reg_rs_bypass_1), .A2(n594), .Y(n9123) );
  INVX1_LVT U6835 ( .A(n5483), .Y(n9120) );
  NAND2X0_LVT U6836 ( .A1(n9120), .A2(io_fpu_dmem_resp_data[0]), .Y(n5482) );
  NAND4X0_LVT U6837 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n5482), .Y(
        n_T_702[0]) );
  NAND2X0_LVT U6838 ( .A1(n_T_918[1]), .A2(n6899), .Y(n9137) );
  NAND2X0_LVT U6839 ( .A1(n_T_635[1]), .A2(n3243), .Y(n9135) );
  NAND2X0_LVT U6840 ( .A1(io_imem_sfence_bits_addr[1]), .A2(n5484), .Y(n9136)
         );
  AO222X1_LVT U6841 ( .A1(mem_br_target_2_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[2]), .A5(n_T_918[2]), .A6(n6855), .Y(N600) );
  AO22X1_LVT U6842 ( .A1(n6860), .A2(io_dmem_resp_bits_data[2]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[2]), .Y(n5485) );
  AO21X1_LVT U6843 ( .A1(n3854), .A2(div_io_resp_bits_data[2]), .A3(n5485), 
        .Y(n5486) );
  NAND2X0_LVT U6844 ( .A1(n4324), .A2(n3958), .Y(n5503) );
  AO22X1_LVT U6845 ( .A1(n3899), .A2(n_T_427[1025]), .A3(n_T_427[194]), .A4(
        n2830), .Y(n5490) );
  AO22X1_LVT U6846 ( .A1(n3832), .A2(n_T_427[66]), .A3(n_T_427[897]), .A4(
        n3896), .Y(n5489) );
  AO22X1_LVT U6847 ( .A1(n2864), .A2(n_T_427[386]), .A3(n_T_427[706]), .A4(
        n3904), .Y(n5488) );
  AO22X1_LVT U6848 ( .A1(n2833), .A2(n_T_427[833]), .A3(n_T_427[2]), .A4(n3913), .Y(n5487) );
  NOR4X1_LVT U6849 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .Y(n5502)
         );
  AOI22X1_LVT U6850 ( .A1(n3838), .A2(n_T_427[450]), .A3(n3871), .A4(
        n_T_427[258]), .Y(n5494) );
  AOI22X1_LVT U6851 ( .A1(n3870), .A2(n_T_427[514]), .A3(n_T_427[578]), .A4(
        n3795), .Y(n5493) );
  OA22X1_LVT U6852 ( .A1(n3519), .A2(n6766), .A3(n3173), .A4(n3083), .Y(n5492)
         );
  AOI22X1_LVT U6853 ( .A1(n3816), .A2(n_T_427[130]), .A3(n_T_427[769]), .A4(
        n3812), .Y(n5491) );
  NAND4X0_LVT U6854 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .Y(n5495) );
  AO22X1_LVT U6855 ( .A1(n3923), .A2(n_T_427[1473]), .A3(n_T_427[1345]), .A4(
        n3917), .Y(n5499) );
  AO22X1_LVT U6856 ( .A1(n3933), .A2(n_T_427[1409]), .A3(n_T_427[1281]), .A4(
        n3927), .Y(n5498) );
  AO22X1_LVT U6857 ( .A1(n3943), .A2(n_T_427[1153]), .A3(n_T_427[1217]), .A4(
        n3937), .Y(n5497) );
  AO22X1_LVT U6858 ( .A1(n3953), .A2(n_T_427[1089]), .A3(n_T_427[961]), .A4(
        n3947), .Y(n5496) );
  NOR4X1_LVT U6859 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .Y(n5500)
         );
  NAND4X0_LVT U6860 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .Y(
        id_rs_1[2]) );
  NAND2X0_LVT U6861 ( .A1(n_T_918[2]), .A2(n6899), .Y(n9150) );
  NAND2X0_LVT U6862 ( .A1(n_T_635[2]), .A2(n6901), .Y(n9149) );
  NAND2X0_LVT U6863 ( .A1(io_imem_sfence_bits_addr[2]), .A2(n6900), .Y(n9148)
         );
  AO222X1_LVT U6864 ( .A1(mem_br_target_3_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[3]), .A5(n_T_918[3]), .A6(n6855), .Y(N601) );
  AO22X1_LVT U6865 ( .A1(n6860), .A2(io_dmem_resp_bits_data[3]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[3]), .Y(n5504) );
  AO21X1_LVT U6866 ( .A1(n3854), .A2(div_io_resp_bits_data[3]), .A3(n5504), 
        .Y(n5505) );
  AO22X1_LVT U6867 ( .A1(n3830), .A2(n_T_427[1793]), .A3(n_T_427[1666]), .A4(
        n3826), .Y(n5509) );
  AO22X1_LVT U6868 ( .A1(n3891), .A2(n_T_427[1538]), .A3(n_T_427[1602]), .A4(
        n3885), .Y(n5508) );
  AO22X1_LVT U6869 ( .A1(n3923), .A2(n_T_427[1474]), .A3(n_T_427[1346]), .A4(
        n3917), .Y(n5507) );
  AO22X1_LVT U6870 ( .A1(n3933), .A2(n_T_427[1410]), .A3(n_T_427[1282]), .A4(
        n3927), .Y(n5506) );
  NOR4X1_LVT U6871 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .Y(n5527)
         );
  AO22X1_LVT U6872 ( .A1(n3943), .A2(n_T_427[1154]), .A3(n_T_427[1218]), .A4(
        n3937), .Y(n5513) );
  AO22X1_LVT U6873 ( .A1(n3953), .A2(n_T_427[1090]), .A3(n_T_427[962]), .A4(
        n3947), .Y(n5512) );
  AO22X1_LVT U6874 ( .A1(n3899), .A2(n_T_427[1026]), .A3(n_T_427[898]), .A4(
        n2831), .Y(n5511) );
  AO22X1_LVT U6875 ( .A1(n3834), .A2(n_T_427[387]), .A3(n_T_427[67]), .A4(
        n3831), .Y(n5510) );
  NOR4X1_LVT U6876 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .Y(n5526)
         );
  AO22X1_LVT U6877 ( .A1(n3907), .A2(n_T_427[770]), .A3(n_T_427[451]), .A4(
        n2824), .Y(n5515) );
  AO22X1_LVT U6878 ( .A1(n2826), .A2(n_T_427[3]), .A3(n_T_427[643]), .A4(n3821), .Y(n5514) );
  AO22X1_LVT U6879 ( .A1(n6796), .A2(n_T_427[131]), .A3(n_T_427[834]), .A4(
        n3875), .Y(n5519) );
  AO22X1_LVT U6880 ( .A1(n6765), .A2(n_T_427[707]), .A3(n3859), .A4(
        n_T_427[195]), .Y(n5518) );
  AO22X1_LVT U6881 ( .A1(n_T_427[515]), .A2(n3868), .A3(n6868), .A4(
        n_T_427[323]), .Y(n5517) );
  AO22X1_LVT U6882 ( .A1(n_T_427[579]), .A2(n3796), .A3(n3871), .A4(
        n_T_427[259]), .Y(n5516) );
  NOR4X1_LVT U6883 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .Y(n5520)
         );
  AOI22X1_LVT U6884 ( .A1(n6764), .A2(n_T_427[1849]), .A3(n_T_427[1730]), .A4(
        n2866), .Y(n5522) );
  NAND2X0_LVT U6885 ( .A1(n4327), .A2(n3957), .Y(n5521) );
  AND3X1_LVT U6886 ( .A1(n5523), .A2(n5522), .A3(n5521), .Y(n5524) );
  NAND4X0_LVT U6887 ( .A1(n5527), .A2(n5524), .A3(n5525), .A4(n5526), .Y(
        id_rs_1[3]) );
  NAND2X0_LVT U6888 ( .A1(n_T_918[3]), .A2(n6899), .Y(n9157) );
  NAND2X0_LVT U6889 ( .A1(n_T_635[3]), .A2(n3243), .Y(n9156) );
  NAND2X0_LVT U6890 ( .A1(io_imem_sfence_bits_addr[3]), .A2(n6900), .Y(n9155)
         );
  AO222X1_LVT U6891 ( .A1(mem_br_target_4_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[4]), .A5(n_T_918[4]), .A6(n6855), .Y(N602) );
  AO22X1_LVT U6892 ( .A1(n6860), .A2(io_dmem_resp_bits_data[4]), .A3(n3847), 
        .A4(io_imem_sfence_bits_addr[4]), .Y(n5528) );
  AO21X1_LVT U6893 ( .A1(n3854), .A2(div_io_resp_bits_data[4]), .A3(n5528), 
        .Y(n5529) );
  AOI22X1_LVT U6894 ( .A1(n6765), .A2(n_T_427[708]), .A3(n3859), .A4(
        n_T_427[196]), .Y(n5533) );
  AOI22X1_LVT U6895 ( .A1(n6871), .A2(n_T_427[835]), .A3(n3871), .A4(
        n_T_427[260]), .Y(n5532) );
  OA22X1_LVT U6896 ( .A1(n3520), .A2(n6766), .A3(n3174), .A4(n3083), .Y(n5531)
         );
  AOI22X1_LVT U6897 ( .A1(n_T_427[899]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[580]), .Y(n5530) );
  NAND4X0_LVT U6898 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .Y(n5534) );
  NAND2X0_LVT U6899 ( .A1(n_T_918[4]), .A2(n6899), .Y(n9161) );
  NAND2X0_LVT U6900 ( .A1(n_T_635[4]), .A2(n6901), .Y(n9160) );
  NAND2X0_LVT U6901 ( .A1(io_imem_sfence_bits_addr[4]), .A2(n6900), .Y(n9159)
         );
  AO222X1_LVT U6902 ( .A1(mem_br_target_5_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[5]), .A5(n_T_918[5]), .A6(n6855), .Y(N603) );
  AO22X1_LVT U6903 ( .A1(n6860), .A2(io_dmem_resp_bits_data[5]), .A3(n3847), 
        .A4(io_imem_sfence_bits_addr[5]), .Y(n5535) );
  AO21X1_LVT U6904 ( .A1(n3854), .A2(div_io_resp_bits_data[5]), .A3(n5535), 
        .Y(n5536) );
  NAND2X0_LVT U6905 ( .A1(n4333), .A2(n3958), .Y(n5554) );
  AO22X1_LVT U6906 ( .A1(n3923), .A2(n_T_427[1476]), .A3(n_T_427[1348]), .A4(
        n3917), .Y(n5540) );
  AO22X1_LVT U6907 ( .A1(n3933), .A2(n_T_427[1412]), .A3(n_T_427[1284]), .A4(
        n3927), .Y(n5539) );
  AO22X1_LVT U6908 ( .A1(n3943), .A2(n_T_427[1156]), .A3(n_T_427[1220]), .A4(
        n3937), .Y(n5538) );
  AO22X1_LVT U6909 ( .A1(n3953), .A2(n_T_427[1092]), .A3(n_T_427[964]), .A4(
        n3947), .Y(n5537) );
  NOR4X1_LVT U6910 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .Y(n5553)
         );
  AOI22X1_LVT U6911 ( .A1(n3797), .A2(n_T_427[581]), .A3(n3867), .A4(
        n_T_427[325]), .Y(n5544) );
  AOI22X1_LVT U6912 ( .A1(n6765), .A2(n_T_427[709]), .A3(n3864), .A4(
        n_T_427[69]), .Y(n5543) );
  AOI22X1_LVT U6913 ( .A1(n3838), .A2(n_T_427[453]), .A3(n_T_427[836]), .A4(
        n3875), .Y(n5542) );
  AOI22X1_LVT U6914 ( .A1(n3863), .A2(n_T_427[645]), .A3(n3865), .A4(
        n_T_427[389]), .Y(n5541) );
  NAND4X0_LVT U6915 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .Y(n5545) );
  AO22X1_LVT U6916 ( .A1(n3899), .A2(n_T_427[1028]), .A3(n_T_427[197]), .A4(
        n2830), .Y(n5550) );
  AO22X1_LVT U6917 ( .A1(n2861), .A2(n_T_427[772]), .A3(n_T_427[900]), .A4(
        n3896), .Y(n5549) );
  AO22X1_LVT U6918 ( .A1(n2826), .A2(n_T_427[5]), .A3(n_T_427[133]), .A4(n3908), .Y(n5548) );
  AO22X1_LVT U6919 ( .A1(n3819), .A2(n_T_427[517]), .A3(n_T_427[261]), .A4(
        n2828), .Y(n5547) );
  NOR4X1_LVT U6920 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .Y(n5551)
         );
  NAND4X0_LVT U6921 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .Y(
        id_rs_1[5]) );
  NAND2X0_LVT U6922 ( .A1(io_fpu_dmem_resp_data[5]), .A2(n9165), .Y(n5558) );
  NAND2X0_LVT U6923 ( .A1(n_T_918[5]), .A2(n6899), .Y(n5557) );
  NAND2X0_LVT U6924 ( .A1(io_imem_sfence_bits_addr[5]), .A2(n6900), .Y(n5556)
         );
  NAND2X0_LVT U6925 ( .A1(n_T_635[5]), .A2(n3243), .Y(n5555) );
  NAND4X0_LVT U6926 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .Y(
        n_T_702[5]) );
  AO222X1_LVT U6927 ( .A1(mem_br_target_6_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[6]), .A5(n6855), .A6(n_T_918[6]), .Y(N604) );
  AO22X1_LVT U6928 ( .A1(n6860), .A2(io_dmem_resp_bits_data[6]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[6]), .Y(n5559) );
  AO21X1_LVT U6929 ( .A1(n3854), .A2(div_io_resp_bits_data[6]), .A3(n5559), 
        .Y(n5560) );
  AO22X1_LVT U6930 ( .A1(n3933), .A2(n_T_427[1413]), .A3(n_T_427[1285]), .A4(
        n3927), .Y(n5564) );
  AO22X1_LVT U6931 ( .A1(n3943), .A2(n_T_427[1157]), .A3(n_T_427[1221]), .A4(
        n3937), .Y(n5563) );
  AO22X1_LVT U6932 ( .A1(n3953), .A2(n_T_427[1093]), .A3(n_T_427[965]), .A4(
        n3947), .Y(n5562) );
  AO22X1_LVT U6933 ( .A1(n3900), .A2(n_T_427[1029]), .A3(n_T_427[70]), .A4(
        n3832), .Y(n5561) );
  NOR4X1_LVT U6934 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .Y(n5577)
         );
  AO22X1_LVT U6935 ( .A1(n3906), .A2(n_T_427[773]), .A3(n_T_427[710]), .A4(
        n2827), .Y(n5566) );
  AO22X1_LVT U6936 ( .A1(n1919), .A2(n_T_427[326]), .A3(n_T_427[6]), .A4(n3914), .Y(n5565) );
  AO22X1_LVT U6937 ( .A1(n6867), .A2(n_T_427[390]), .A3(n3859), .A4(
        n_T_427[198]), .Y(n5570) );
  AO22X1_LVT U6938 ( .A1(n3870), .A2(n_T_427[518]), .A3(n_T_427[454]), .A4(
        n3836), .Y(n5569) );
  AO22X1_LVT U6939 ( .A1(n_T_427[901]), .A2(n3811), .A3(n3871), .A4(
        n_T_427[262]), .Y(n5568) );
  AO22X1_LVT U6940 ( .A1(n3816), .A2(n_T_427[134]), .A3(n_T_427[837]), .A4(
        n3874), .Y(n5567) );
  NOR4X1_LVT U6941 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .Y(n5571)
         );
  AOI22X1_LVT U6942 ( .A1(n3915), .A2(n_T_427[582]), .A3(n_T_427[646]), .A4(
        n6812), .Y(n5573) );
  NAND2X0_LVT U6943 ( .A1(n4336), .A2(n3958), .Y(n5572) );
  AND3X1_LVT U6944 ( .A1(n5574), .A2(n5573), .A3(n5572), .Y(n5575) );
  NAND4X0_LVT U6945 ( .A1(n5577), .A2(n5578), .A3(n5576), .A4(n5575), .Y(
        id_rs_1[6]) );
  NAND2X0_LVT U6946 ( .A1(io_fpu_dmem_resp_data[6]), .A2(n9165), .Y(n5582) );
  NAND2X0_LVT U6947 ( .A1(n_T_918[6]), .A2(n6899), .Y(n5581) );
  NAND2X0_LVT U6948 ( .A1(io_imem_sfence_bits_addr[6]), .A2(n6900), .Y(n5580)
         );
  NAND2X0_LVT U6949 ( .A1(n_T_635[6]), .A2(n3243), .Y(n5579) );
  NAND4X0_LVT U6950 ( .A1(n5582), .A2(n5581), .A3(n5580), .A4(n5579), .Y(
        n_T_702[6]) );
  AO222X1_LVT U6951 ( .A1(mem_br_target_7_), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[7]), .A5(n6855), .A6(n_T_918[7]), .Y(N605) );
  AO22X1_LVT U6952 ( .A1(n6860), .A2(io_dmem_resp_bits_data[7]), .A3(n3847), 
        .A4(io_imem_sfence_bits_addr[7]), .Y(n5583) );
  AO21X1_LVT U6953 ( .A1(n3854), .A2(div_io_resp_bits_data[7]), .A3(n5583), 
        .Y(n5584) );
  AO22X1_LVT U6954 ( .A1(n3829), .A2(n_T_427[1797]), .A3(n_T_427[1670]), .A4(
        n3825), .Y(n5588) );
  AO22X1_LVT U6955 ( .A1(n3891), .A2(n_T_427[1542]), .A3(n_T_427[1606]), .A4(
        n3885), .Y(n5587) );
  AO22X1_LVT U6956 ( .A1(n3923), .A2(n_T_427[1478]), .A3(n_T_427[1350]), .A4(
        n3917), .Y(n5586) );
  AO22X1_LVT U6957 ( .A1(n3933), .A2(n_T_427[1414]), .A3(n_T_427[1286]), .A4(
        n3927), .Y(n5585) );
  NOR4X1_LVT U6958 ( .A1(n5588), .A2(n5587), .A3(n5586), .A4(n5585), .Y(n5602)
         );
  AO22X1_LVT U6959 ( .A1(n2860), .A2(n_T_427[774]), .A3(n_T_427[391]), .A4(
        n2865), .Y(n5590) );
  AO22X1_LVT U6960 ( .A1(n1918), .A2(n_T_427[327]), .A3(n_T_427[583]), .A4(
        n2870), .Y(n5589) );
  NOR2X0_LVT U6961 ( .A1(n5590), .A2(n5589), .Y(n5600) );
  AO22X1_LVT U6962 ( .A1(n_T_427[647]), .A2(n3863), .A3(n3804), .A4(
        n_T_427[711]), .Y(n5594) );
  AO22X1_LVT U6963 ( .A1(n3870), .A2(n_T_427[519]), .A3(n_T_427[455]), .A4(
        n3836), .Y(n5593) );
  AO22X1_LVT U6964 ( .A1(n_T_427[838]), .A2(n6871), .A3(n3871), .A4(
        n_T_427[263]), .Y(n5592) );
  AO22X1_LVT U6965 ( .A1(n3816), .A2(n_T_427[135]), .A3(n6838), .A4(n_T_427[7]), .Y(n5591) );
  NOR4X1_LVT U6966 ( .A1(n5594), .A2(n5593), .A3(n5592), .A4(n5591), .Y(n5595)
         );
  AOI22X1_LVT U6967 ( .A1(n3801), .A2(n_T_427[1853]), .A3(n_T_427[1734]), .A4(
        n2866), .Y(n5597) );
  NAND2X0_LVT U6968 ( .A1(n4339), .A2(n3958), .Y(n5596) );
  AND3X1_LVT U6969 ( .A1(n5598), .A2(n5597), .A3(n5596), .Y(n5599) );
  NAND4X0_LVT U6970 ( .A1(n5602), .A2(n5601), .A3(n5600), .A4(n5599), .Y(
        id_rs_1[7]) );
  AO22X1_LVT U6971 ( .A1(n6860), .A2(io_dmem_resp_bits_data[8]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[8]), .Y(n5603) );
  AO21X1_LVT U6972 ( .A1(n3854), .A2(div_io_resp_bits_data[8]), .A3(n5603), 
        .Y(n5604) );
  AO22X1_LVT U6973 ( .A1(n3933), .A2(n_T_427[1415]), .A3(n_T_427[1287]), .A4(
        n3927), .Y(n5608) );
  AO22X1_LVT U6974 ( .A1(n3943), .A2(n_T_427[1159]), .A3(n_T_427[1223]), .A4(
        n3937), .Y(n5607) );
  AO22X1_LVT U6975 ( .A1(n3953), .A2(n_T_427[1095]), .A3(n_T_427[967]), .A4(
        n3947), .Y(n5606) );
  AO22X1_LVT U6976 ( .A1(n3900), .A2(n_T_427[1031]), .A3(n_T_427[903]), .A4(
        n2831), .Y(n5605) );
  NOR4X1_LVT U6977 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .Y(n5621)
         );
  AO22X1_LVT U6978 ( .A1(n3907), .A2(n_T_427[775]), .A3(n_T_427[72]), .A4(
        n2871), .Y(n5610) );
  AO22X1_LVT U6979 ( .A1(n3911), .A2(n_T_427[456]), .A3(n_T_427[8]), .A4(n3913), .Y(n5609) );
  NOR2X0_LVT U6980 ( .A1(n5610), .A2(n5609), .Y(n5620) );
  AO22X1_LVT U6981 ( .A1(n6765), .A2(n_T_427[712]), .A3(n3865), .A4(
        n_T_427[392]), .Y(n5614) );
  AO22X1_LVT U6982 ( .A1(n_T_427[648]), .A2(n3863), .A3(n3859), .A4(
        n_T_427[200]), .Y(n5613) );
  AO22X1_LVT U6983 ( .A1(n3870), .A2(n_T_427[520]), .A3(n_T_427[584]), .A4(
        n3795), .Y(n5612) );
  AO22X1_LVT U6984 ( .A1(n6796), .A2(n_T_427[136]), .A3(n_T_427[839]), .A4(
        n3875), .Y(n5611) );
  NOR4X1_LVT U6985 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .Y(n5615)
         );
  AOI22X1_LVT U6986 ( .A1(n3817), .A2(n_T_427[328]), .A3(n_T_427[264]), .A4(
        n3810), .Y(n5617) );
  NAND2X0_LVT U6987 ( .A1(n4342), .A2(n3959), .Y(n5616) );
  AND3X1_LVT U6988 ( .A1(n5618), .A2(n5617), .A3(n5616), .Y(n5619) );
  NAND4X0_LVT U6989 ( .A1(n5621), .A2(n5622), .A3(n5620), .A4(n5619), .Y(
        id_rs_1[8]) );
  NAND2X0_LVT U6990 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[8]), .Y(n5626) );
  NAND2X0_LVT U6991 ( .A1(n6899), .A2(n_T_918[8]), .Y(n5625) );
  NAND2X0_LVT U6992 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[8]), .Y(n5624)
         );
  NAND2X0_LVT U6993 ( .A1(n6901), .A2(n_T_635[8]), .Y(n5623) );
  NAND4X0_LVT U6994 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .Y(
        n_T_702[8]) );
  AO22X1_LVT U6995 ( .A1(n6860), .A2(io_dmem_resp_bits_data[9]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[9]), .Y(n5627) );
  AO21X1_LVT U6996 ( .A1(n3854), .A2(div_io_resp_bits_data[9]), .A3(n5627), 
        .Y(n5628) );
  AO22X1_LVT U6997 ( .A1(n3934), .A2(n_T_427[1416]), .A3(n_T_427[1288]), .A4(
        n3927), .Y(n5632) );
  AO22X1_LVT U6998 ( .A1(n3944), .A2(n_T_427[1160]), .A3(n_T_427[1224]), .A4(
        n3937), .Y(n5631) );
  AO22X1_LVT U6999 ( .A1(n3954), .A2(n_T_427[1096]), .A3(n_T_427[968]), .A4(
        n3947), .Y(n5630) );
  AO22X1_LVT U7000 ( .A1(n3899), .A2(n_T_427[1032]), .A3(n_T_427[201]), .A4(
        n3806), .Y(n5629) );
  NOR4X1_LVT U7001 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .Y(n5645)
         );
  AO22X1_LVT U7002 ( .A1(n3834), .A2(n_T_427[393]), .A3(n_T_427[73]), .A4(
        n3833), .Y(n5634) );
  AO22X1_LVT U7003 ( .A1(n3817), .A2(n_T_427[329]), .A3(n_T_427[713]), .A4(
        n3903), .Y(n5633) );
  NOR2X0_LVT U7004 ( .A1(n5634), .A2(n5633), .Y(n5644) );
  AO22X1_LVT U7005 ( .A1(n3797), .A2(n_T_427[585]), .A3(n_T_427[457]), .A4(
        n3836), .Y(n5638) );
  AO22X1_LVT U7006 ( .A1(n_T_427[904]), .A2(n3811), .A3(n3871), .A4(
        n_T_427[265]), .Y(n5637) );
  AO22X1_LVT U7007 ( .A1(n3814), .A2(n_T_427[776]), .A3(n_T_427[840]), .A4(
        n3874), .Y(n5636) );
  AO22X1_LVT U7008 ( .A1(n3816), .A2(n_T_427[137]), .A3(n6838), .A4(n_T_427[9]), .Y(n5635) );
  NOR4X1_LVT U7009 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .Y(n5639)
         );
  AOI22X1_LVT U7010 ( .A1(n2851), .A2(n_T_427[521]), .A3(n_T_427[649]), .A4(
        n3821), .Y(n5641) );
  NAND2X0_LVT U7011 ( .A1(n4345), .A2(n3958), .Y(n5640) );
  AND3X1_LVT U7012 ( .A1(n5642), .A2(n5641), .A3(n5640), .Y(n5643) );
  NAND4X0_LVT U7013 ( .A1(n5645), .A2(n5646), .A3(n5644), .A4(n5643), .Y(
        id_rs_1[9]) );
  NAND2X0_LVT U7014 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[9]), .Y(n5650) );
  NAND2X0_LVT U7015 ( .A1(n6899), .A2(n_T_918[9]), .Y(n5649) );
  NAND2X0_LVT U7016 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[9]), .Y(n5648)
         );
  NAND2X0_LVT U7017 ( .A1(n3243), .A2(n_T_635[9]), .Y(n5647) );
  NAND4X0_LVT U7018 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .Y(
        n_T_702[9]) );
  AO22X1_LVT U7019 ( .A1(n3851), .A2(io_dmem_resp_bits_data[10]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[10]), .Y(n5651) );
  AO21X1_LVT U7020 ( .A1(n3854), .A2(div_io_resp_bits_data[10]), .A3(n5651), 
        .Y(n5652) );
  AO22X1_LVT U7021 ( .A1(n3933), .A2(n_T_427[1417]), .A3(n_T_427[1289]), .A4(
        n3927), .Y(n5656) );
  AO22X1_LVT U7022 ( .A1(n3943), .A2(n_T_427[1161]), .A3(n_T_427[1225]), .A4(
        n3937), .Y(n5655) );
  AO22X1_LVT U7023 ( .A1(n3953), .A2(n_T_427[1097]), .A3(n_T_427[969]), .A4(
        n3947), .Y(n5654) );
  AO22X1_LVT U7024 ( .A1(n3900), .A2(n_T_427[1033]), .A3(n3806), .A4(
        n_T_427[202]), .Y(n5653) );
  NOR4X1_LVT U7025 ( .A1(n5656), .A2(n5655), .A3(n5654), .A4(n5653), .Y(n5669)
         );
  AO22X1_LVT U7026 ( .A1(n2864), .A2(n_T_427[394]), .A3(n_T_427[458]), .A4(
        n3912), .Y(n5658) );
  AO22X1_LVT U7027 ( .A1(n3833), .A2(n_T_427[74]), .A3(n_T_427[905]), .A4(
        n3897), .Y(n5657) );
  AO22X1_LVT U7028 ( .A1(n_T_427[650]), .A2(n3863), .A3(n3804), .A4(
        n_T_427[714]), .Y(n5662) );
  AO22X1_LVT U7029 ( .A1(n3814), .A2(n_T_427[777]), .A3(n_T_427[841]), .A4(
        n3874), .Y(n5661) );
  AO22X1_LVT U7030 ( .A1(n_T_427[522]), .A2(n3868), .A3(n3872), .A4(
        n_T_427[266]), .Y(n5660) );
  AO22X1_LVT U7031 ( .A1(n6796), .A2(n_T_427[138]), .A3(n3839), .A4(
        n_T_427[10]), .Y(n5659) );
  NOR4X1_LVT U7032 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .Y(n5663)
         );
  AOI22X1_LVT U7033 ( .A1(n2857), .A2(n_T_427[330]), .A3(n_T_427[586]), .A4(
        n2869), .Y(n5665) );
  NAND2X0_LVT U7034 ( .A1(n4348), .A2(n3958), .Y(n5664) );
  AND3X1_LVT U7035 ( .A1(n5666), .A2(n5665), .A3(n5664), .Y(n5667) );
  NAND4X0_LVT U7036 ( .A1(n5669), .A2(n5670), .A3(n5668), .A4(n5667), .Y(
        id_rs_1[10]) );
  NAND2X0_LVT U7037 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[10]), .Y(n5674) );
  NAND2X0_LVT U7038 ( .A1(n6899), .A2(n_T_918[10]), .Y(n5673) );
  NAND2X0_LVT U7039 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[10]), .Y(n5672)
         );
  NAND2X0_LVT U7040 ( .A1(n3243), .A2(n_T_635[10]), .Y(n5671) );
  NAND4X0_LVT U7041 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .Y(
        n_T_702[10]) );
  AO22X1_LVT U7042 ( .A1(n2861), .A2(n_T_427[778]), .A3(n_T_427[587]), .A4(
        n3915), .Y(n5676) );
  AO22X1_LVT U7043 ( .A1(n3896), .A2(n_T_427[906]), .A3(n_T_427[139]), .A4(
        n3908), .Y(n5675) );
  AO22X1_LVT U7044 ( .A1(n6867), .A2(n_T_427[395]), .A3(n3859), .A4(
        n_T_427[203]), .Y(n5680) );
  AO22X1_LVT U7045 ( .A1(n_T_427[715]), .A2(n3804), .A3(n3864), .A4(
        n_T_427[75]), .Y(n5679) );
  AO22X1_LVT U7046 ( .A1(n_T_427[651]), .A2(n3863), .A3(n3867), .A4(
        n_T_427[331]), .Y(n5678) );
  AO22X1_LVT U7047 ( .A1(n3837), .A2(n_T_427[459]), .A3(n3872), .A4(
        n_T_427[267]), .Y(n5677) );
  NOR4X1_LVT U7048 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .Y(n5681)
         );
  AO22X1_LVT U7049 ( .A1(n3851), .A2(io_dmem_resp_bits_data[12]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[12]), .Y(n5682) );
  AO21X1_LVT U7050 ( .A1(n3854), .A2(div_io_resp_bits_data[12]), .A3(n5682), 
        .Y(n5683) );
  AO22X1_LVT U7051 ( .A1(n3933), .A2(n_T_427[1419]), .A3(n_T_427[1291]), .A4(
        n3927), .Y(n5687) );
  AO22X1_LVT U7052 ( .A1(n3943), .A2(n_T_427[1163]), .A3(n_T_427[1227]), .A4(
        n3937), .Y(n5686) );
  AO22X1_LVT U7053 ( .A1(n3953), .A2(n_T_427[1099]), .A3(n_T_427[971]), .A4(
        n3947), .Y(n5685) );
  AO22X1_LVT U7054 ( .A1(n3900), .A2(n_T_427[1035]), .A3(n_T_427[76]), .A4(
        n2871), .Y(n5684) );
  NOR4X1_LVT U7055 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .Y(n5700)
         );
  AO22X1_LVT U7056 ( .A1(n2856), .A2(n_T_427[332]), .A3(n_T_427[588]), .A4(
        n3916), .Y(n5689) );
  AO22X1_LVT U7057 ( .A1(n3907), .A2(n_T_427[779]), .A3(n_T_427[716]), .A4(
        n3903), .Y(n5688) );
  AO22X1_LVT U7058 ( .A1(n6867), .A2(n_T_427[396]), .A3(n3859), .A4(
        n_T_427[204]), .Y(n5693) );
  AO22X1_LVT U7059 ( .A1(n3870), .A2(n_T_427[524]), .A3(n_T_427[460]), .A4(
        n3836), .Y(n5692) );
  AO22X1_LVT U7060 ( .A1(n_T_427[907]), .A2(n3811), .A3(n3872), .A4(
        n_T_427[268]), .Y(n5691) );
  AO22X1_LVT U7061 ( .A1(n3816), .A2(n_T_427[140]), .A3(n6838), .A4(
        n_T_427[12]), .Y(n5690) );
  NOR4X1_LVT U7062 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .Y(n5694)
         );
  AOI22X1_LVT U7063 ( .A1(n2833), .A2(n_T_427[843]), .A3(n_T_427[652]), .A4(
        n2829), .Y(n5696) );
  NAND2X0_LVT U7064 ( .A1(n4354), .A2(n3958), .Y(n5695) );
  AND3X1_LVT U7065 ( .A1(n5697), .A2(n5696), .A3(n5695), .Y(n5698) );
  NAND4X0_LVT U7066 ( .A1(n5700), .A2(n5701), .A3(n5699), .A4(n5698), .Y(
        id_rs_1[12]) );
  NAND2X0_LVT U7067 ( .A1(io_fpu_dmem_resp_data[12]), .A2(n9165), .Y(n5705) );
  NAND2X0_LVT U7068 ( .A1(n_T_918[12]), .A2(n6899), .Y(n5704) );
  NAND2X0_LVT U7069 ( .A1(io_imem_sfence_bits_addr[12]), .A2(n6900), .Y(n5703)
         );
  NAND2X0_LVT U7070 ( .A1(n_T_635[12]), .A2(n6901), .Y(n5702) );
  NAND4X0_LVT U7071 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .Y(
        n_T_702[12]) );
  AO22X1_LVT U7072 ( .A1(n3851), .A2(io_dmem_resp_bits_data[13]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[13]), .Y(n5706) );
  AO21X1_LVT U7073 ( .A1(n3855), .A2(div_io_resp_bits_data[13]), .A3(n5706), 
        .Y(n5707) );
  AO22X1_LVT U7074 ( .A1(n3832), .A2(n_T_427[77]), .A3(n_T_427[717]), .A4(
        n3905), .Y(n5718) );
  AO22X1_LVT U7075 ( .A1(n2826), .A2(n_T_427[13]), .A3(n_T_427[141]), .A4(
        n3908), .Y(n5717) );
  AO22X1_LVT U7076 ( .A1(n2857), .A2(n_T_427[333]), .A3(n_T_427[525]), .A4(
        n3818), .Y(n5716) );
  AO22X1_LVT U7077 ( .A1(n_T_427[653]), .A2(n3863), .A3(n3796), .A4(
        n_T_427[589]), .Y(n5711) );
  AO22X1_LVT U7078 ( .A1(n6867), .A2(n_T_427[397]), .A3(n3859), .A4(
        n_T_427[205]), .Y(n5710) );
  AO22X1_LVT U7079 ( .A1(n_T_427[461]), .A2(n3837), .A3(n3872), .A4(
        n_T_427[269]), .Y(n5709) );
  AO22X1_LVT U7080 ( .A1(n3814), .A2(n_T_427[780]), .A3(n_T_427[844]), .A4(
        n3875), .Y(n5708) );
  NOR4X1_LVT U7081 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .Y(n5712)
         );
  NAND2X0_LVT U7082 ( .A1(n4356), .A2(n3958), .Y(n5713) );
  NAND2X0_LVT U7083 ( .A1(n5714), .A2(n5713), .Y(n5715) );
  NOR4X1_LVT U7084 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), .Y(n5725)
         );
  AO22X1_LVT U7085 ( .A1(n3933), .A2(n_T_427[1420]), .A3(n_T_427[1292]), .A4(
        n3927), .Y(n5722) );
  AO22X1_LVT U7086 ( .A1(n3943), .A2(n_T_427[1164]), .A3(n_T_427[1228]), .A4(
        n3938), .Y(n5721) );
  AO22X1_LVT U7087 ( .A1(n3953), .A2(n_T_427[1100]), .A3(n_T_427[972]), .A4(
        n3948), .Y(n5720) );
  AO22X1_LVT U7088 ( .A1(n3899), .A2(n_T_427[1036]), .A3(n_T_427[908]), .A4(
        n3897), .Y(n5719) );
  NOR4X1_LVT U7089 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .Y(n5723)
         );
  NAND3X0_LVT U7090 ( .A1(n5725), .A2(n5724), .A3(n5723), .Y(id_rs_1[13]) );
  NAND2X0_LVT U7091 ( .A1(io_fpu_dmem_resp_data[13]), .A2(n9165), .Y(n5729) );
  NAND2X0_LVT U7092 ( .A1(n_T_918[13]), .A2(n6899), .Y(n5728) );
  NAND2X0_LVT U7093 ( .A1(io_imem_sfence_bits_addr[13]), .A2(n6900), .Y(n5727)
         );
  NAND2X0_LVT U7094 ( .A1(n_T_635[13]), .A2(n6901), .Y(n5726) );
  NAND4X0_LVT U7095 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .Y(
        n_T_702[13]) );
  AO22X1_LVT U7096 ( .A1(n3851), .A2(io_dmem_resp_bits_data[14]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[14]), .Y(n5730) );
  AO21X1_LVT U7097 ( .A1(n3855), .A2(div_io_resp_bits_data[14]), .A3(n5730), 
        .Y(n5731) );
  AO22X1_LVT U7098 ( .A1(n_T_427[909]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[462]), .Y(n5735) );
  AO22X1_LVT U7099 ( .A1(n_T_427[654]), .A2(n3863), .A3(n3859), .A4(
        n_T_427[206]), .Y(n5734) );
  AO22X1_LVT U7100 ( .A1(n_T_427[718]), .A2(n3804), .A3(n3864), .A4(
        n_T_427[78]), .Y(n5733) );
  AO22X1_LVT U7101 ( .A1(n3816), .A2(n_T_427[142]), .A3(n3872), .A4(
        n_T_427[270]), .Y(n5732) );
  OR4X1_LVT U7102 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .Y(n5736)
         );
  AO22X1_LVT U7103 ( .A1(n3835), .A2(n_T_427[398]), .A3(n_T_427[1037]), .A4(
        n3898), .Y(n5740) );
  AO22X1_LVT U7104 ( .A1(n3906), .A2(n_T_427[781]), .A3(n_T_427[14]), .A4(
        n2826), .Y(n5739) );
  AO22X1_LVT U7105 ( .A1(n2856), .A2(n_T_427[334]), .A3(n_T_427[590]), .A4(
        n2870), .Y(n5738) );
  AO22X1_LVT U7106 ( .A1(n2850), .A2(n_T_427[526]), .A3(n_T_427[845]), .A4(
        n6813), .Y(n5737) );
  NAND2X0_LVT U7107 ( .A1(io_fpu_dmem_resp_data[14]), .A2(n9165), .Y(n5744) );
  NAND2X0_LVT U7108 ( .A1(n_T_918[14]), .A2(n6899), .Y(n5743) );
  NAND2X0_LVT U7109 ( .A1(io_imem_sfence_bits_addr[14]), .A2(n6900), .Y(n5742)
         );
  NAND2X0_LVT U7110 ( .A1(n_T_635[14]), .A2(n6901), .Y(n5741) );
  NAND4X0_LVT U7111 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .Y(
        n_T_702[14]) );
  AO22X1_LVT U7112 ( .A1(n3851), .A2(io_dmem_resp_bits_data[15]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[15]), .Y(n5745) );
  AO21X1_LVT U7113 ( .A1(n3855), .A2(div_io_resp_bits_data[15]), .A3(n5745), 
        .Y(n5746) );
  AO22X1_LVT U7114 ( .A1(n3835), .A2(n_T_427[399]), .A3(n_T_427[79]), .A4(
        n3833), .Y(n5757) );
  AO22X1_LVT U7115 ( .A1(n2860), .A2(n_T_427[782]), .A3(n_T_427[463]), .A4(
        n3911), .Y(n5756) );
  AO22X1_LVT U7116 ( .A1(n1919), .A2(n_T_427[335]), .A3(n_T_427[591]), .A4(
        n3916), .Y(n5755) );
  AO22X1_LVT U7117 ( .A1(n_T_427[655]), .A2(n3863), .A3(n3804), .A4(
        n_T_427[719]), .Y(n5750) );
  AO22X1_LVT U7118 ( .A1(n_T_427[910]), .A2(n3811), .A3(n3868), .A4(
        n_T_427[527]), .Y(n5749) );
  AO22X1_LVT U7119 ( .A1(n_T_427[846]), .A2(n3874), .A3(n3872), .A4(
        n_T_427[271]), .Y(n5748) );
  AO22X1_LVT U7120 ( .A1(n3816), .A2(n_T_427[143]), .A3(n3840), .A4(
        n_T_427[15]), .Y(n5747) );
  NOR4X1_LVT U7121 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .Y(n5751)
         );
  NAND2X0_LVT U7122 ( .A1(n4361), .A2(n3958), .Y(n5752) );
  NAND2X0_LVT U7123 ( .A1(n5753), .A2(n5752), .Y(n5754) );
  NOR4X1_LVT U7124 ( .A1(n5757), .A2(n5756), .A3(n5755), .A4(n5754), .Y(n5764)
         );
  AO22X1_LVT U7125 ( .A1(n3934), .A2(n_T_427[1422]), .A3(n_T_427[1294]), .A4(
        n3928), .Y(n5761) );
  AO22X1_LVT U7126 ( .A1(n3944), .A2(n_T_427[1166]), .A3(n_T_427[1230]), .A4(
        n3938), .Y(n5760) );
  AO22X1_LVT U7127 ( .A1(n3954), .A2(n_T_427[1102]), .A3(n_T_427[974]), .A4(
        n3948), .Y(n5759) );
  AO22X1_LVT U7128 ( .A1(n3899), .A2(n_T_427[1038]), .A3(n_T_427[207]), .A4(
        n3806), .Y(n5758) );
  NOR4X1_LVT U7129 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .Y(n5762)
         );
  NAND3X0_LVT U7130 ( .A1(n5764), .A2(n5763), .A3(n5762), .Y(id_rs_1[15]) );
  NAND2X0_LVT U7131 ( .A1(io_fpu_dmem_resp_data[15]), .A2(n9165), .Y(n5768) );
  NAND2X0_LVT U7132 ( .A1(n_T_918[15]), .A2(n6899), .Y(n5767) );
  NAND2X0_LVT U7133 ( .A1(io_imem_sfence_bits_addr[15]), .A2(n6900), .Y(n5766)
         );
  NAND2X0_LVT U7134 ( .A1(n_T_635[15]), .A2(n6901), .Y(n5765) );
  NAND4X0_LVT U7135 ( .A1(n5768), .A2(n5767), .A3(n5766), .A4(n5765), .Y(
        n_T_702[15]) );
  NAND2X0_LVT U7136 ( .A1(csr_io_rw_rdata[16]), .A2(n3844), .Y(n5771) );
  AOI22X1_LVT U7137 ( .A1(n3852), .A2(io_dmem_resp_bits_data[16]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[16]), .Y(n5770) );
  NAND2X0_LVT U7138 ( .A1(div_io_resp_bits_data[16]), .A2(n3856), .Y(n5769) );
  NAND3X0_LVT U7139 ( .A1(n5771), .A2(n5770), .A3(n5769), .Y(
        n_T_427__T_1136_data[16]) );
  AOI22X1_LVT U7140 ( .A1(n3870), .A2(n_T_427[528]), .A3(n3867), .A4(
        n_T_427[336]), .Y(n5775) );
  AOI22X1_LVT U7141 ( .A1(n3874), .A2(n_T_427[847]), .A3(n3840), .A4(
        n_T_427[16]), .Y(n5774) );
  OA22X1_LVT U7142 ( .A1(n3521), .A2(n6423), .A3(n3175), .A4(n6422), .Y(n5773)
         );
  AOI22X1_LVT U7143 ( .A1(n_T_427[911]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[592]), .Y(n5772) );
  NAND4X0_LVT U7144 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .Y(n5776) );
  NAND2X0_LVT U7145 ( .A1(csr_io_rw_rdata[17]), .A2(n3844), .Y(n5779) );
  AOI22X1_LVT U7146 ( .A1(n3852), .A2(io_dmem_resp_bits_data[17]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[17]), .Y(n5778) );
  NAND2X0_LVT U7147 ( .A1(div_io_resp_bits_data[17]), .A2(n3858), .Y(n5777) );
  NAND3X0_LVT U7148 ( .A1(n5779), .A2(n5778), .A3(n5777), .Y(
        n_T_427__T_1136_data[17]) );
  AO22X1_LVT U7149 ( .A1(n3816), .A2(n_T_427[145]), .A3(n_T_427[784]), .A4(
        n3812), .Y(n5783) );
  AO22X1_LVT U7150 ( .A1(n3797), .A2(n_T_427[593]), .A3(n_T_427[465]), .A4(
        n3836), .Y(n5782) );
  AO22X1_LVT U7151 ( .A1(n_T_427[912]), .A2(n3811), .A3(n3872), .A4(
        n_T_427[273]), .Y(n5781) );
  AO22X1_LVT U7152 ( .A1(n3859), .A2(n_T_427[209]), .A3(n3864), .A4(
        n_T_427[81]), .Y(n5780) );
  NOR4X1_LVT U7153 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .Y(n5784)
         );
  OA22X1_LVT U7154 ( .A1(n3541), .A2(n3799), .A3(n3139), .A4(n3803), .Y(n5787)
         );
  OA22X1_LVT U7155 ( .A1(n3142), .A2(n3081), .A3(n3494), .A4(n3082), .Y(n5786)
         );
  AOI22X1_LVT U7156 ( .A1(n3894), .A2(n_T_427[1552]), .A3(n_T_427[1616]), .A4(
        n3889), .Y(n5785) );
  AND4X1_LVT U7157 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .Y(n5796)
         );
  AO22X1_LVT U7158 ( .A1(n3924), .A2(n_T_427[1488]), .A3(n_T_427[1360]), .A4(
        n3918), .Y(n5792) );
  AO22X1_LVT U7159 ( .A1(n3934), .A2(n_T_427[1424]), .A3(n_T_427[1296]), .A4(
        n3928), .Y(n5791) );
  AO22X1_LVT U7160 ( .A1(n3944), .A2(n_T_427[1168]), .A3(n_T_427[1232]), .A4(
        n3938), .Y(n5790) );
  AO22X1_LVT U7161 ( .A1(n3954), .A2(n_T_427[1104]), .A3(n_T_427[976]), .A4(
        n3948), .Y(n5789) );
  NOR4X1_LVT U7162 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .Y(n5795)
         );
  NAND2X0_LVT U7163 ( .A1(n3958), .A2(n4367), .Y(n5793) );
  NAND4X0_LVT U7164 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .Y(
        id_rs_1[17]) );
  NAND2X0_LVT U7165 ( .A1(io_fpu_dmem_resp_data[17]), .A2(n9165), .Y(n5800) );
  NAND2X0_LVT U7166 ( .A1(n_T_918[17]), .A2(n6899), .Y(n5799) );
  NAND2X0_LVT U7167 ( .A1(io_imem_sfence_bits_addr[17]), .A2(n6900), .Y(n5798)
         );
  NAND2X0_LVT U7168 ( .A1(n_T_635[17]), .A2(n3243), .Y(n5797) );
  NAND4X0_LVT U7169 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .Y(
        n_T_702[17]) );
  AO22X1_LVT U7170 ( .A1(n3852), .A2(io_dmem_resp_bits_data[18]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[18]), .Y(n5801) );
  AO21X1_LVT U7171 ( .A1(n3855), .A2(div_io_resp_bits_data[18]), .A3(n5801), 
        .Y(n5802) );
  AO21X1_LVT U7172 ( .A1(n3843), .A2(csr_io_rw_rdata[18]), .A3(n5802), .Y(
        n_T_427__T_1136_data[18]) );
  AO22X1_LVT U7173 ( .A1(n3934), .A2(n_T_427[1425]), .A3(n_T_427[1297]), .A4(
        n3928), .Y(n5806) );
  AO22X1_LVT U7174 ( .A1(n3944), .A2(n_T_427[1169]), .A3(n_T_427[1233]), .A4(
        n3938), .Y(n5805) );
  AO22X1_LVT U7175 ( .A1(n3954), .A2(n_T_427[1105]), .A3(n_T_427[977]), .A4(
        n3948), .Y(n5804) );
  AO22X1_LVT U7176 ( .A1(n3900), .A2(n_T_427[1041]), .A3(n_T_427[913]), .A4(
        n2832), .Y(n5803) );
  NOR4X1_LVT U7177 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .Y(n5819)
         );
  AO22X1_LVT U7178 ( .A1(n2824), .A2(n_T_427[466]), .A3(n_T_427[722]), .A4(
        n3904), .Y(n5808) );
  AO22X1_LVT U7179 ( .A1(n2826), .A2(n_T_427[18]), .A3(n_T_427[146]), .A4(
        n3909), .Y(n5807) );
  NOR2X0_LVT U7180 ( .A1(n5808), .A2(n5807), .Y(n5818) );
  AOI22X1_LVT U7181 ( .A1(n2833), .A2(n_T_427[849]), .A3(n_T_427[274]), .A4(
        n2828), .Y(n5816) );
  NAND2X0_LVT U7182 ( .A1(n4370), .A2(n3959), .Y(n5815) );
  AO22X1_LVT U7183 ( .A1(n_T_427[658]), .A2(n3862), .A3(n3859), .A4(
        n_T_427[210]), .Y(n5812) );
  AO22X1_LVT U7184 ( .A1(n3813), .A2(n_T_427[785]), .A3(n_T_427[594]), .A4(
        n3795), .Y(n5811) );
  AO22X1_LVT U7185 ( .A1(n6867), .A2(n_T_427[402]), .A3(n3864), .A4(
        n_T_427[82]), .Y(n5810) );
  AO22X1_LVT U7186 ( .A1(n_T_427[530]), .A2(n3868), .A3(n6868), .A4(
        n_T_427[338]), .Y(n5809) );
  NOR4X1_LVT U7187 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .Y(n5813)
         );
  AND3X1_LVT U7188 ( .A1(n5816), .A2(n5815), .A3(n5814), .Y(n5817) );
  NAND4X0_LVT U7189 ( .A1(n5819), .A2(n5820), .A3(n5818), .A4(n5817), .Y(
        id_rs_1[18]) );
  NAND2X0_LVT U7190 ( .A1(io_fpu_dmem_resp_data[18]), .A2(n9165), .Y(n5824) );
  NAND2X0_LVT U7191 ( .A1(n_T_918[18]), .A2(n6899), .Y(n5823) );
  NAND2X0_LVT U7192 ( .A1(io_imem_sfence_bits_addr[18]), .A2(n6900), .Y(n5822)
         );
  NAND2X0_LVT U7193 ( .A1(n_T_635[18]), .A2(n3243), .Y(n5821) );
  NAND4X0_LVT U7194 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .Y(
        n_T_702[18]) );
  AO22X1_LVT U7195 ( .A1(n3852), .A2(io_dmem_resp_bits_data[19]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[19]), .Y(n5825) );
  AO21X1_LVT U7196 ( .A1(n3855), .A2(div_io_resp_bits_data[19]), .A3(n5825), 
        .Y(n5826) );
  AO21X1_LVT U7197 ( .A1(n3843), .A2(csr_io_rw_rdata[19]), .A3(n5826), .Y(
        n_T_427__T_1136_data[19]) );
  AO22X1_LVT U7198 ( .A1(n_T_427[659]), .A2(n3862), .A3(n3804), .A4(
        n_T_427[723]), .Y(n5830) );
  AO22X1_LVT U7199 ( .A1(n_T_427[914]), .A2(n3811), .A3(n3875), .A4(
        n_T_427[850]), .Y(n5829) );
  AO22X1_LVT U7200 ( .A1(n3869), .A2(n_T_427[531]), .A3(n_T_427[595]), .A4(
        n3795), .Y(n5828) );
  AO22X1_LVT U7201 ( .A1(n3815), .A2(n_T_427[147]), .A3(n3840), .A4(
        n_T_427[19]), .Y(n5827) );
  NOR4X1_LVT U7202 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .Y(n5831)
         );
  OA22X1_LVT U7203 ( .A1(n3543), .A2(n3881), .A3(n3878), .A4(n5831), .Y(n5833)
         );
  NAND2X0_LVT U7204 ( .A1(n4373), .A2(n3959), .Y(n5832) );
  NAND2X0_LVT U7205 ( .A1(io_fpu_dmem_resp_data[19]), .A2(n9165), .Y(n5837) );
  NAND2X0_LVT U7206 ( .A1(n_T_918[19]), .A2(n6899), .Y(n5836) );
  NAND2X0_LVT U7207 ( .A1(io_imem_sfence_bits_addr[19]), .A2(n6900), .Y(n5835)
         );
  NAND2X0_LVT U7208 ( .A1(n_T_635[19]), .A2(n3243), .Y(n5834) );
  NAND4X0_LVT U7209 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .Y(
        n_T_702[19]) );
  AO22X1_LVT U7210 ( .A1(n3852), .A2(io_dmem_resp_bits_data[20]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[20]), .Y(n5838) );
  AO21X1_LVT U7211 ( .A1(n3855), .A2(div_io_resp_bits_data[20]), .A3(n5838), 
        .Y(n5839) );
  AO21X1_LVT U7212 ( .A1(n3844), .A2(csr_io_rw_rdata[20]), .A3(n5839), .Y(
        n_T_427__T_1136_data[20]) );
  AO22X1_LVT U7213 ( .A1(n3933), .A2(n_T_427[1427]), .A3(n_T_427[1299]), .A4(
        n3928), .Y(n5843) );
  AO22X1_LVT U7214 ( .A1(n3943), .A2(n_T_427[1171]), .A3(n_T_427[1235]), .A4(
        n3938), .Y(n5842) );
  AO22X1_LVT U7215 ( .A1(n3953), .A2(n_T_427[1107]), .A3(n_T_427[979]), .A4(
        n3948), .Y(n5841) );
  AO22X1_LVT U7216 ( .A1(n3900), .A2(n_T_427[1043]), .A3(n_T_427[915]), .A4(
        n3896), .Y(n5840) );
  NOR4X1_LVT U7217 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .Y(n5856)
         );
  AO22X1_LVT U7218 ( .A1(n3835), .A2(n_T_427[404]), .A3(n_T_427[724]), .A4(
        n2827), .Y(n5845) );
  AO22X1_LVT U7219 ( .A1(n3913), .A2(n_T_427[20]), .A3(n_T_427[148]), .A4(
        n2863), .Y(n5844) );
  AO22X1_LVT U7220 ( .A1(n3869), .A2(n_T_427[532]), .A3(n_T_427[596]), .A4(
        n3795), .Y(n5849) );
  AO22X1_LVT U7221 ( .A1(n_T_427[660]), .A2(n3862), .A3(n3866), .A4(
        n_T_427[340]), .Y(n5848) );
  AO22X1_LVT U7222 ( .A1(n3813), .A2(n_T_427[787]), .A3(n_T_427[468]), .A4(
        n3836), .Y(n5847) );
  AO22X1_LVT U7223 ( .A1(n3860), .A2(n_T_427[212]), .A3(n6866), .A4(
        n_T_427[84]), .Y(n5846) );
  NOR4X1_LVT U7224 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .Y(n5850)
         );
  OA22X1_LVT U7225 ( .A1(n3544), .A2(n3881), .A3(n3878), .A4(n5850), .Y(n5853)
         );
  AOI22X1_LVT U7226 ( .A1(n3823), .A2(n_T_427[851]), .A3(n_T_427[276]), .A4(
        n3809), .Y(n5852) );
  NAND2X0_LVT U7227 ( .A1(n4376), .A2(n3959), .Y(n5851) );
  AND3X1_LVT U7228 ( .A1(n5853), .A2(n5852), .A3(n5851), .Y(n5854) );
  NAND4X0_LVT U7229 ( .A1(n5856), .A2(n5857), .A3(n5855), .A4(n5854), .Y(
        id_rs_1[20]) );
  NAND2X0_LVT U7230 ( .A1(io_fpu_dmem_resp_data[20]), .A2(n9165), .Y(n5861) );
  NAND2X0_LVT U7231 ( .A1(n_T_918[20]), .A2(n6899), .Y(n5860) );
  NAND2X0_LVT U7232 ( .A1(io_imem_sfence_bits_addr[20]), .A2(n6900), .Y(n5859)
         );
  NAND2X0_LVT U7233 ( .A1(n_T_635[20]), .A2(n6901), .Y(n5858) );
  NAND4X0_LVT U7234 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .Y(
        n_T_702[20]) );
  AO22X1_LVT U7235 ( .A1(n3852), .A2(io_dmem_resp_bits_data[21]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[21]), .Y(n5862) );
  AO21X1_LVT U7236 ( .A1(n3855), .A2(div_io_resp_bits_data[21]), .A3(n5862), 
        .Y(n5863) );
  AO22X1_LVT U7237 ( .A1(n_T_427[916]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[597]), .Y(n5867) );
  AO22X1_LVT U7238 ( .A1(n_T_427[661]), .A2(n3862), .A3(n3859), .A4(
        n_T_427[213]), .Y(n5866) );
  AO22X1_LVT U7239 ( .A1(n_T_427[725]), .A2(n6765), .A3(n3864), .A4(
        n_T_427[85]), .Y(n5865) );
  AO22X1_LVT U7240 ( .A1(n_T_427[852]), .A2(n3875), .A3(n3839), .A4(
        n_T_427[21]), .Y(n5864) );
  NOR4X1_LVT U7241 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .Y(n5868)
         );
  OA22X1_LVT U7242 ( .A1(n3095), .A2(n3596), .A3(n3878), .A4(n5868), .Y(n5870)
         );
  NAND2X0_LVT U7243 ( .A1(n_T_427[533]), .A2(n3819), .Y(n5869) );
  AO22X1_LVT U7244 ( .A1(n3921), .A2(n_T_427[1364]), .A3(n_T_427[1428]), .A4(
        n3932), .Y(n5874) );
  AO22X1_LVT U7245 ( .A1(n3928), .A2(n_T_427[1300]), .A3(n_T_427[1172]), .A4(
        n3942), .Y(n5873) );
  AO22X1_LVT U7246 ( .A1(n3941), .A2(n_T_427[1236]), .A3(n_T_427[1108]), .A4(
        n3952), .Y(n5872) );
  AO22X1_LVT U7247 ( .A1(n3951), .A2(n_T_427[980]), .A3(n_T_427[1044]), .A4(
        n3898), .Y(n5871) );
  NOR4X1_LVT U7248 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .Y(n5875)
         );
  NAND3X0_LVT U7249 ( .A1(n5877), .A2(n5876), .A3(n5875), .Y(id_rs_1[21]) );
  NAND2X0_LVT U7250 ( .A1(io_fpu_dmem_resp_data[21]), .A2(n9165), .Y(n5881) );
  NAND2X0_LVT U7251 ( .A1(n_T_918[21]), .A2(n6899), .Y(n5880) );
  NAND2X0_LVT U7252 ( .A1(io_imem_sfence_bits_addr[21]), .A2(n6900), .Y(n5879)
         );
  NAND2X0_LVT U7253 ( .A1(n_T_635[21]), .A2(n6901), .Y(n5878) );
  NAND4X0_LVT U7254 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .Y(
        n_T_702[21]) );
  AO22X1_LVT U7255 ( .A1(n3921), .A2(n_T_427[1365]), .A3(n_T_427[1429]), .A4(
        n3932), .Y(n5885) );
  AO22X1_LVT U7256 ( .A1(n3931), .A2(n_T_427[1301]), .A3(n_T_427[1173]), .A4(
        n3942), .Y(n5884) );
  AO22X1_LVT U7257 ( .A1(n3941), .A2(n_T_427[1237]), .A3(n_T_427[1109]), .A4(
        n3952), .Y(n5883) );
  AO22X1_LVT U7258 ( .A1(n3951), .A2(n_T_427[981]), .A3(n_T_427[1045]), .A4(
        n3899), .Y(n5882) );
  NOR4X1_LVT U7259 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .Y(n5896)
         );
  AO22X1_LVT U7260 ( .A1(n6765), .A2(n_T_427[726]), .A3(n3865), .A4(
        n_T_427[406]), .Y(n5889) );
  AO22X1_LVT U7261 ( .A1(n_T_427[662]), .A2(n3862), .A3(n3860), .A4(
        n_T_427[214]), .Y(n5888) );
  AO22X1_LVT U7262 ( .A1(n_T_427[853]), .A2(n6871), .A3(n3872), .A4(
        n_T_427[278]), .Y(n5887) );
  AO22X1_LVT U7263 ( .A1(n3815), .A2(n_T_427[150]), .A3(n_T_427[789]), .A4(
        n3812), .Y(n5886) );
  NOR4X1_LVT U7264 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .Y(n5890)
         );
  OA22X1_LVT U7265 ( .A1(n3094), .A2(n3596), .A3(n3878), .A4(n5890), .Y(n5893)
         );
  AOI22X1_LVT U7266 ( .A1(n2850), .A2(n_T_427[534]), .A3(n_T_427[22]), .A4(
        n3913), .Y(n5892) );
  NAND2X0_LVT U7267 ( .A1(n_T_427[598]), .A2(n2870), .Y(n5891) );
  AND3X1_LVT U7268 ( .A1(n5893), .A2(n5892), .A3(n5891), .Y(n5894) );
  NAND4X0_LVT U7269 ( .A1(n5897), .A2(n5895), .A3(n5896), .A4(n5894), .Y(
        id_rs_1[22]) );
  NAND2X0_LVT U7270 ( .A1(io_fpu_dmem_resp_data[22]), .A2(n9165), .Y(n5901) );
  NAND2X0_LVT U7271 ( .A1(n_T_918[22]), .A2(n6899), .Y(n5900) );
  NAND2X0_LVT U7272 ( .A1(io_imem_sfence_bits_addr[22]), .A2(n6900), .Y(n5899)
         );
  NAND2X0_LVT U7273 ( .A1(n_T_635[22]), .A2(n3243), .Y(n5898) );
  NAND4X0_LVT U7274 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .Y(
        n_T_702[22]) );
  NAND2X0_LVT U7275 ( .A1(csr_io_rw_rdata[23]), .A2(n3844), .Y(n5904) );
  AOI22X1_LVT U7276 ( .A1(n3852), .A2(io_dmem_resp_bits_data[23]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[23]), .Y(n5903) );
  NAND2X0_LVT U7277 ( .A1(div_io_resp_bits_data[23]), .A2(n3858), .Y(n5902) );
  NAND3X0_LVT U7278 ( .A1(n5904), .A2(n5903), .A3(n5902), .Y(
        n_T_427__T_1136_data[23]) );
  AOI22X1_LVT U7279 ( .A1(n3870), .A2(n_T_427[535]), .A3(n_T_427[599]), .A4(
        n3795), .Y(n5910) );
  AOI22X1_LVT U7280 ( .A1(n3814), .A2(n_T_427[790]), .A3(n3871), .A4(
        n_T_427[279]), .Y(n5909) );
  AOI22X1_LVT U7281 ( .A1(n6765), .A2(n_T_427[727]), .A3(n6868), .A4(
        n_T_427[343]), .Y(n5908) );
  OA22X1_LVT U7282 ( .A1(n5906), .A2(n3526), .A3(n3177), .A4(n5905), .Y(n5907)
         );
  NAND4X0_LVT U7283 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .Y(n5911) );
  AO22X1_LVT U7284 ( .A1(n3924), .A2(n_T_427[1494]), .A3(n_T_427[1366]), .A4(
        n3918), .Y(n5915) );
  AO22X1_LVT U7285 ( .A1(n3934), .A2(n_T_427[1430]), .A3(n_T_427[1302]), .A4(
        n3928), .Y(n5914) );
  AO22X1_LVT U7286 ( .A1(n3944), .A2(n_T_427[1174]), .A3(n_T_427[1238]), .A4(
        n3938), .Y(n5913) );
  AO22X1_LVT U7287 ( .A1(n3954), .A2(n_T_427[1110]), .A3(n_T_427[982]), .A4(
        n3948), .Y(n5912) );
  NOR4X1_LVT U7288 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .Y(n5922)
         );
  AO22X1_LVT U7289 ( .A1(n2865), .A2(n_T_427[407]), .A3(n_T_427[471]), .A4(
        n3911), .Y(n5919) );
  AO22X1_LVT U7290 ( .A1(n3900), .A2(n_T_427[1046]), .A3(n_T_427[215]), .A4(
        n3808), .Y(n5918) );
  AO22X1_LVT U7291 ( .A1(n2871), .A2(n_T_427[87]), .A3(n_T_427[918]), .A4(
        n3897), .Y(n5917) );
  AO22X1_LVT U7292 ( .A1(n2833), .A2(n_T_427[854]), .A3(n_T_427[663]), .A4(
        n3820), .Y(n5916) );
  NOR4X1_LVT U7293 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .Y(n5921)
         );
  NAND2X0_LVT U7294 ( .A1(n3957), .A2(n4383), .Y(n5920) );
  NAND4X0_LVT U7295 ( .A1(n5922), .A2(n5923), .A3(n5921), .A4(n5920), .Y(
        id_rs_1[23]) );
  NAND2X0_LVT U7296 ( .A1(io_fpu_dmem_resp_data[23]), .A2(n9165), .Y(n5927) );
  NAND2X0_LVT U7297 ( .A1(n_T_918[23]), .A2(n6899), .Y(n5926) );
  NAND2X0_LVT U7298 ( .A1(io_imem_sfence_bits_addr[23]), .A2(n6900), .Y(n5925)
         );
  NAND2X0_LVT U7299 ( .A1(n_T_635[23]), .A2(n3243), .Y(n5924) );
  NAND4X0_LVT U7300 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .Y(
        n_T_702[23]) );
  AO22X1_LVT U7301 ( .A1(n3852), .A2(io_dmem_resp_bits_data[24]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[24]), .Y(n5928) );
  AO21X1_LVT U7302 ( .A1(n3855), .A2(div_io_resp_bits_data[24]), .A3(n5928), 
        .Y(n5929) );
  AO21X1_LVT U7303 ( .A1(n3844), .A2(csr_io_rw_rdata[24]), .A3(n5929), .Y(
        n_T_427__T_1136_data[24]) );
  AO22X1_LVT U7304 ( .A1(n3944), .A2(n_T_427[1175]), .A3(n_T_427[1239]), .A4(
        n3938), .Y(n5933) );
  AO22X1_LVT U7305 ( .A1(n3954), .A2(n_T_427[1111]), .A3(n_T_427[983]), .A4(
        n3948), .Y(n5932) );
  AO22X1_LVT U7306 ( .A1(n3900), .A2(n_T_427[1047]), .A3(n_T_427[216]), .A4(
        n2830), .Y(n5931) );
  AO22X1_LVT U7307 ( .A1(n3907), .A2(n_T_427[791]), .A3(n_T_427[408]), .A4(
        n3834), .Y(n5930) );
  NOR4X1_LVT U7308 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .Y(n5946)
         );
  AO22X1_LVT U7309 ( .A1(n3817), .A2(n_T_427[344]), .A3(n_T_427[600]), .A4(
        n2869), .Y(n5935) );
  AO22X1_LVT U7310 ( .A1(n3912), .A2(n_T_427[472]), .A3(n_T_427[24]), .A4(
        n2879), .Y(n5934) );
  NAND2X0_LVT U7311 ( .A1(n4386), .A2(n3959), .Y(n5943) );
  AO22X1_LVT U7312 ( .A1(n_T_427[664]), .A2(n3862), .A3(n3868), .A4(
        n_T_427[536]), .Y(n5939) );
  AO22X1_LVT U7313 ( .A1(n3815), .A2(n_T_427[152]), .A3(n_T_427[855]), .A4(
        n3874), .Y(n5938) );
  AO22X1_LVT U7314 ( .A1(n_T_427[728]), .A2(n6765), .A3(n3864), .A4(
        n_T_427[88]), .Y(n5937) );
  AO22X1_LVT U7315 ( .A1(n_T_427[919]), .A2(n3811), .A3(n3872), .A4(
        n_T_427[280]), .Y(n5936) );
  NOR4X1_LVT U7316 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .Y(n5940)
         );
  OA22X1_LVT U7317 ( .A1(n3545), .A2(n3881), .A3(n3878), .A4(n5940), .Y(n5942)
         );
  OA22X1_LVT U7318 ( .A1(n3546), .A2(n3799), .A3(n3137), .A4(n3803), .Y(n5941)
         );
  AND3X1_LVT U7319 ( .A1(n5943), .A2(n5942), .A3(n5941), .Y(n5944) );
  NAND4X0_LVT U7320 ( .A1(n5946), .A2(n5947), .A3(n5945), .A4(n5944), .Y(
        id_rs_1[24]) );
  NAND2X0_LVT U7321 ( .A1(io_fpu_dmem_resp_data[24]), .A2(n9165), .Y(n5951) );
  NAND2X0_LVT U7322 ( .A1(n_T_918[24]), .A2(n6899), .Y(n5950) );
  NAND2X0_LVT U7323 ( .A1(io_imem_sfence_bits_addr[24]), .A2(n6900), .Y(n5949)
         );
  NAND2X0_LVT U7324 ( .A1(n_T_635[24]), .A2(n6901), .Y(n5948) );
  NAND4X0_LVT U7325 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .Y(
        n_T_702[24]) );
  AO22X1_LVT U7326 ( .A1(n3852), .A2(io_dmem_resp_bits_data[25]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[25]), .Y(n5952) );
  AO21X1_LVT U7327 ( .A1(n3855), .A2(div_io_resp_bits_data[25]), .A3(n5952), 
        .Y(n5953) );
  AO22X1_LVT U7328 ( .A1(n3907), .A2(n_T_427[792]), .A3(n_T_427[217]), .A4(
        n3807), .Y(n5964) );
  AO22X1_LVT U7329 ( .A1(n2872), .A2(n_T_427[89]), .A3(n_T_427[153]), .A4(
        n3909), .Y(n5963) );
  AO22X1_LVT U7330 ( .A1(n2824), .A2(n_T_427[473]), .A3(n_T_427[537]), .A4(
        n2851), .Y(n5962) );
  AO22X1_LVT U7331 ( .A1(n_T_427[920]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[601]), .Y(n5957) );
  AO22X1_LVT U7332 ( .A1(n3804), .A2(n_T_427[729]), .A3(n3865), .A4(
        n_T_427[409]), .Y(n5956) );
  AO22X1_LVT U7333 ( .A1(n_T_427[665]), .A2(n3862), .A3(n3867), .A4(
        n_T_427[345]), .Y(n5955) );
  AO22X1_LVT U7334 ( .A1(n_T_427[856]), .A2(n3875), .A3(n3872), .A4(
        n_T_427[281]), .Y(n5954) );
  NOR4X1_LVT U7335 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .Y(n5958)
         );
  OA22X1_LVT U7336 ( .A1(n3097), .A2(n3596), .A3(n3878), .A4(n5958), .Y(n5960)
         );
  NAND2X0_LVT U7337 ( .A1(n_T_427[25]), .A2(n3914), .Y(n5959) );
  NAND2X0_LVT U7338 ( .A1(n5960), .A2(n5959), .Y(n5961) );
  AO22X1_LVT U7339 ( .A1(n2866), .A2(n_T_427[1752]), .A3(n_T_427[1814]), .A4(
        n3829), .Y(n5967) );
  AO22X1_LVT U7340 ( .A1(n_T_427[1868]), .A2(n3802), .A3(n3884), .A4(
        n_T_427[1906]), .Y(n5966) );
  AO22X1_LVT U7341 ( .A1(n3826), .A2(n_T_427[1688]), .A3(n_T_427[1560]), .A4(
        n3890), .Y(n5965) );
  NAND2X0_LVT U7342 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[25]), .Y(n5971) );
  NAND2X0_LVT U7343 ( .A1(n_T_918[25]), .A2(n6899), .Y(n5970) );
  NAND2X0_LVT U7344 ( .A1(io_imem_sfence_bits_addr[25]), .A2(n6900), .Y(n5969)
         );
  NAND2X0_LVT U7345 ( .A1(n_T_635[25]), .A2(n6901), .Y(n5968) );
  NAND4X0_LVT U7346 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .Y(
        n_T_702[25]) );
  AO22X1_LVT U7347 ( .A1(n3852), .A2(io_dmem_resp_bits_data[26]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[26]), .Y(n5972) );
  AO21X1_LVT U7348 ( .A1(n3855), .A2(div_io_resp_bits_data[26]), .A3(n5972), 
        .Y(n5973) );
  AO22X1_LVT U7349 ( .A1(n3921), .A2(n_T_427[1369]), .A3(n_T_427[1433]), .A4(
        n3932), .Y(n5977) );
  AO22X1_LVT U7350 ( .A1(n3931), .A2(n_T_427[1305]), .A3(n_T_427[1177]), .A4(
        n3942), .Y(n5976) );
  AO22X1_LVT U7351 ( .A1(n3941), .A2(n_T_427[1241]), .A3(n_T_427[1113]), .A4(
        n3952), .Y(n5975) );
  AO22X1_LVT U7352 ( .A1(n3951), .A2(n_T_427[985]), .A3(n_T_427[1049]), .A4(
        n3898), .Y(n5974) );
  NOR4X1_LVT U7353 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .Y(n5990)
         );
  AO22X1_LVT U7354 ( .A1(n3831), .A2(n_T_427[90]), .A3(n_T_427[218]), .A4(
        n2830), .Y(n5979) );
  AO22X1_LVT U7355 ( .A1(n2857), .A2(n_T_427[346]), .A3(n_T_427[921]), .A4(
        n3895), .Y(n5978) );
  AO22X1_LVT U7356 ( .A1(n6765), .A2(n_T_427[730]), .A3(n_T_427[602]), .A4(
        n3795), .Y(n5983) );
  AO22X1_LVT U7357 ( .A1(n3813), .A2(n_T_427[793]), .A3(n_T_427[857]), .A4(
        n3874), .Y(n5982) );
  AO22X1_LVT U7358 ( .A1(n3837), .A2(n_T_427[474]), .A3(n3872), .A4(
        n_T_427[282]), .Y(n5981) );
  AO22X1_LVT U7359 ( .A1(n3815), .A2(n_T_427[154]), .A3(n6838), .A4(
        n_T_427[26]), .Y(n5980) );
  NOR4X1_LVT U7360 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .Y(n5984)
         );
  OA22X1_LVT U7361 ( .A1(n3096), .A2(n3596), .A3(n3878), .A4(n5984), .Y(n5987)
         );
  AOI22X1_LVT U7362 ( .A1(n3835), .A2(n_T_427[410]), .A3(n_T_427[666]), .A4(
        n3820), .Y(n5986) );
  NAND2X0_LVT U7363 ( .A1(n_T_427[538]), .A2(n3818), .Y(n5985) );
  AND3X1_LVT U7364 ( .A1(n5987), .A2(n5986), .A3(n5985), .Y(n5988) );
  NAND4X0_LVT U7365 ( .A1(n5990), .A2(n5991), .A3(n5989), .A4(n5988), .Y(
        id_rs_1[26]) );
  NAND2X0_LVT U7366 ( .A1(io_fpu_dmem_resp_data[26]), .A2(n9165), .Y(n5995) );
  NAND2X0_LVT U7367 ( .A1(n_T_918[26]), .A2(n6899), .Y(n5994) );
  NAND2X0_LVT U7368 ( .A1(io_imem_sfence_bits_addr[26]), .A2(n6900), .Y(n5993)
         );
  NAND2X0_LVT U7369 ( .A1(n_T_635[26]), .A2(n3243), .Y(n5992) );
  NAND4X0_LVT U7370 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .Y(
        n_T_702[26]) );
  AO22X1_LVT U7371 ( .A1(n3852), .A2(io_dmem_resp_bits_data[27]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[27]), .Y(n5996) );
  AO21X1_LVT U7372 ( .A1(n3856), .A2(div_io_resp_bits_data[27]), .A3(n5996), 
        .Y(n5997) );
  AO21X1_LVT U7373 ( .A1(n3843), .A2(csr_io_rw_rdata[27]), .A3(n5997), .Y(
        n_T_427__T_1136_data[27]) );
  AOI22X1_LVT U7374 ( .A1(n3797), .A2(n_T_427[603]), .A3(n3871), .A4(
        n_T_427[283]), .Y(n6001) );
  AOI22X1_LVT U7375 ( .A1(n3814), .A2(n_T_427[794]), .A3(n_T_427[858]), .A4(
        n3875), .Y(n6000) );
  AOI22X1_LVT U7376 ( .A1(n6765), .A2(n_T_427[731]), .A3(n3864), .A4(
        n_T_427[91]), .Y(n5999) );
  AOI22X1_LVT U7377 ( .A1(n3863), .A2(n_T_427[667]), .A3(n3865), .A4(
        n_T_427[411]), .Y(n5998) );
  NAND4X0_LVT U7378 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .Y(n6002) );
  NAND2X0_LVT U7379 ( .A1(n6877), .A2(n6002), .Y(n6005) );
  NAND2X0_LVT U7380 ( .A1(n3957), .A2(n4393), .Y(n6004) );
  NAND2X0_LVT U7381 ( .A1(n_T_427[1908]), .A2(n3884), .Y(n6003) );
  AO22X1_LVT U7382 ( .A1(n3934), .A2(n_T_427[1434]), .A3(n_T_427[1306]), .A4(
        n3928), .Y(n6009) );
  AO22X1_LVT U7383 ( .A1(n3944), .A2(n_T_427[1178]), .A3(n_T_427[1242]), .A4(
        n3938), .Y(n6008) );
  AO22X1_LVT U7384 ( .A1(n3954), .A2(n_T_427[1114]), .A3(n_T_427[986]), .A4(
        n3948), .Y(n6007) );
  AO22X1_LVT U7385 ( .A1(n3900), .A2(n_T_427[1050]), .A3(n_T_427[219]), .A4(
        n2830), .Y(n6006) );
  NOR4X1_LVT U7386 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .Y(n6010)
         );
  NAND3X0_LVT U7387 ( .A1(n6012), .A2(n6011), .A3(n6010), .Y(id_rs_1[27]) );
  AO22X1_LVT U7388 ( .A1(n3851), .A2(io_dmem_resp_bits_data[28]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[28]), .Y(n6013) );
  AO21X1_LVT U7389 ( .A1(n3855), .A2(div_io_resp_bits_data[28]), .A3(n6013), 
        .Y(n6014) );
  AO22X1_LVT U7390 ( .A1(n2864), .A2(n_T_427[412]), .A3(n_T_427[220]), .A4(
        n3807), .Y(n6025) );
  AO22X1_LVT U7391 ( .A1(n2871), .A2(n_T_427[92]), .A3(n_T_427[28]), .A4(n3914), .Y(n6024) );
  AO22X1_LVT U7392 ( .A1(n3910), .A2(n_T_427[476]), .A3(n3810), .A4(
        n_T_427[284]), .Y(n6023) );
  AO22X1_LVT U7393 ( .A1(n_T_427[668]), .A2(n3862), .A3(n3804), .A4(
        n_T_427[732]), .Y(n6018) );
  AO22X1_LVT U7394 ( .A1(n_T_427[923]), .A2(n3811), .A3(n3875), .A4(
        n_T_427[859]), .Y(n6017) );
  AO22X1_LVT U7395 ( .A1(n3815), .A2(n_T_427[156]), .A3(n_T_427[795]), .A4(
        n3812), .Y(n6016) );
  AO22X1_LVT U7396 ( .A1(n_T_427[540]), .A2(n3869), .A3(n3866), .A4(
        n_T_427[348]), .Y(n6015) );
  NOR4X1_LVT U7397 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .Y(n6019)
         );
  OA22X1_LVT U7398 ( .A1(n3596), .A2(n3090), .A3(n3878), .A4(n6019), .Y(n6021)
         );
  NAND2X0_LVT U7399 ( .A1(n_T_427[604]), .A2(n3915), .Y(n6020) );
  NAND2X0_LVT U7400 ( .A1(n6021), .A2(n6020), .Y(n6022) );
  NAND2X0_LVT U7401 ( .A1(io_fpu_dmem_resp_data[28]), .A2(n9165), .Y(n6029) );
  NAND2X0_LVT U7402 ( .A1(n_T_918[28]), .A2(n6899), .Y(n6028) );
  NAND2X0_LVT U7403 ( .A1(io_imem_sfence_bits_addr[28]), .A2(n6900), .Y(n6027)
         );
  NAND2X0_LVT U7404 ( .A1(n_T_635[28]), .A2(n3243), .Y(n6026) );
  NAND4X0_LVT U7405 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .Y(
        n_T_702[28]) );
  AO22X1_LVT U7406 ( .A1(n3851), .A2(io_dmem_resp_bits_data[29]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[29]), .Y(n6030) );
  AO21X1_LVT U7407 ( .A1(n3856), .A2(div_io_resp_bits_data[29]), .A3(n6030), 
        .Y(n6031) );
  AO21X1_LVT U7408 ( .A1(n3843), .A2(csr_io_rw_rdata[29]), .A3(n6031), .Y(
        n_T_427__T_1136_data[29]) );
  AO22X1_LVT U7409 ( .A1(n3831), .A2(n_T_427[93]), .A3(n_T_427[221]), .A4(
        n3808), .Y(n6041) );
  AO22X1_LVT U7410 ( .A1(n2832), .A2(n_T_427[924]), .A3(n_T_427[29]), .A4(
        n2879), .Y(n6040) );
  AO22X1_LVT U7411 ( .A1(n2865), .A2(n_T_427[413]), .A3(n_T_427[860]), .A4(
        n3823), .Y(n6039) );
  AOI22X1_LVT U7412 ( .A1(n3797), .A2(n_T_427[605]), .A3(n3867), .A4(
        n_T_427[349]), .Y(n6035) );
  AOI22X1_LVT U7413 ( .A1(n_T_427[477]), .A2(n3837), .A3(n3871), .A4(
        n_T_427[285]), .Y(n6034) );
  AOI22X1_LVT U7414 ( .A1(n3816), .A2(n_T_427[157]), .A3(n_T_427[796]), .A4(
        n3812), .Y(n6033) );
  AOI22X1_LVT U7415 ( .A1(n3863), .A2(n_T_427[669]), .A3(n3804), .A4(
        n_T_427[733]), .Y(n6032) );
  NAND4X0_LVT U7416 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .Y(n6036) );
  AO22X1_LVT U7417 ( .A1(n3957), .A2(n4398), .A3(n6036), .A4(n6877), .Y(n6037)
         );
  AO21X1_LVT U7418 ( .A1(n_T_427[541]), .A2(n3819), .A3(n6037), .Y(n6038) );
  NOR4X1_LVT U7419 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .Y(n6048)
         );
  AO22X1_LVT U7420 ( .A1(n3921), .A2(n_T_427[1372]), .A3(n_T_427[1436]), .A4(
        n3932), .Y(n6045) );
  AO22X1_LVT U7421 ( .A1(n3931), .A2(n_T_427[1308]), .A3(n_T_427[1180]), .A4(
        n3942), .Y(n6044) );
  AO22X1_LVT U7422 ( .A1(n3941), .A2(n_T_427[1244]), .A3(n_T_427[1116]), .A4(
        n3952), .Y(n6043) );
  AO22X1_LVT U7423 ( .A1(n3951), .A2(n_T_427[988]), .A3(n_T_427[1052]), .A4(
        n3899), .Y(n6042) );
  NOR4X1_LVT U7424 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .Y(n6046)
         );
  NAND3X0_LVT U7425 ( .A1(n6048), .A2(n6047), .A3(n6046), .Y(id_rs_1[29]) );
  NAND2X0_LVT U7426 ( .A1(io_fpu_dmem_resp_data[29]), .A2(n9165), .Y(n6052) );
  NAND2X0_LVT U7427 ( .A1(n_T_918[29]), .A2(n6899), .Y(n6051) );
  NAND2X0_LVT U7428 ( .A1(io_imem_sfence_bits_addr[29]), .A2(n6900), .Y(n6050)
         );
  NAND2X0_LVT U7429 ( .A1(n_T_635[29]), .A2(n3243), .Y(n6049) );
  NAND4X0_LVT U7430 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .Y(
        n_T_702[29]) );
  AO22X1_LVT U7431 ( .A1(n3851), .A2(io_dmem_resp_bits_data[30]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[30]), .Y(n6053) );
  AO21X1_LVT U7432 ( .A1(n3856), .A2(div_io_resp_bits_data[30]), .A3(n6053), 
        .Y(n6054) );
  AO21X1_LVT U7433 ( .A1(n3843), .A2(csr_io_rw_rdata[30]), .A3(n6054), .Y(
        n_T_427__T_1136_data[30]) );
  AO22X1_LVT U7434 ( .A1(n3830), .A2(n_T_427[1819]), .A3(n_T_427[1693]), .A4(
        n3827), .Y(n6058) );
  AO22X1_LVT U7435 ( .A1(n3892), .A2(n_T_427[1565]), .A3(n_T_427[1629]), .A4(
        n3886), .Y(n6057) );
  AO22X1_LVT U7436 ( .A1(n3924), .A2(n_T_427[1501]), .A3(n_T_427[1373]), .A4(
        n3918), .Y(n6056) );
  AO22X1_LVT U7437 ( .A1(n3934), .A2(n_T_427[1437]), .A3(n_T_427[1309]), .A4(
        n3928), .Y(n6055) );
  NOR4X1_LVT U7438 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .Y(n6076)
         );
  AO22X1_LVT U7439 ( .A1(n3944), .A2(n_T_427[1181]), .A3(n_T_427[1245]), .A4(
        n3938), .Y(n6062) );
  AO22X1_LVT U7440 ( .A1(n3954), .A2(n_T_427[1117]), .A3(n_T_427[989]), .A4(
        n3948), .Y(n6061) );
  AO22X1_LVT U7441 ( .A1(n3900), .A2(n_T_427[1053]), .A3(n_T_427[222]), .A4(
        n3806), .Y(n6060) );
  AO22X1_LVT U7442 ( .A1(n2865), .A2(n_T_427[414]), .A3(n_T_427[734]), .A4(
        n3904), .Y(n6059) );
  NOR4X1_LVT U7443 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .Y(n6075)
         );
  AO22X1_LVT U7444 ( .A1(n1918), .A2(n_T_427[350]), .A3(n_T_427[478]), .A4(
        n3910), .Y(n6064) );
  AO22X1_LVT U7445 ( .A1(n2851), .A2(n_T_427[542]), .A3(n_T_427[861]), .A4(
        n3822), .Y(n6063) );
  NOR2X0_LVT U7446 ( .A1(n6064), .A2(n6063), .Y(n6074) );
  AO22X1_LVT U7447 ( .A1(n_T_427[925]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[606]), .Y(n6068) );
  AO22X1_LVT U7448 ( .A1(n_T_427[670]), .A2(n3862), .A3(n3864), .A4(
        n_T_427[94]), .Y(n6067) );
  AO22X1_LVT U7449 ( .A1(n_T_427[797]), .A2(n3812), .A3(n3872), .A4(
        n_T_427[286]), .Y(n6066) );
  AO22X1_LVT U7450 ( .A1(n3815), .A2(n_T_427[158]), .A3(n3840), .A4(
        n_T_427[30]), .Y(n6065) );
  NOR4X1_LVT U7451 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .Y(n6069)
         );
  OA22X1_LVT U7452 ( .A1(n3547), .A2(n3881), .A3(n3878), .A4(n6069), .Y(n6072)
         );
  OA22X1_LVT U7453 ( .A1(n3548), .A2(n3799), .A3(n3140), .A4(n3803), .Y(n6071)
         );
  NAND2X0_LVT U7454 ( .A1(n4401), .A2(n3959), .Y(n6070) );
  AND3X1_LVT U7455 ( .A1(n6072), .A2(n6071), .A3(n6070), .Y(n6073) );
  NAND4X0_LVT U7456 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .Y(
        id_rs_1[30]) );
  NAND2X0_LVT U7457 ( .A1(io_fpu_dmem_resp_data[30]), .A2(n9165), .Y(n6080) );
  NAND2X0_LVT U7458 ( .A1(n_T_918[30]), .A2(n6899), .Y(n6079) );
  NAND2X0_LVT U7459 ( .A1(io_imem_sfence_bits_addr[30]), .A2(n6900), .Y(n6078)
         );
  NAND2X0_LVT U7460 ( .A1(n_T_635[30]), .A2(n6901), .Y(n6077) );
  NAND4X0_LVT U7461 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .Y(
        n_T_702[30]) );
  AO22X1_LVT U7462 ( .A1(n6856), .A2(io_fpu_toint_data[31]), .A3(n6855), .A4(
        n_T_918[31]), .Y(n6081) );
  AO21X1_LVT U7463 ( .A1(mem_br_target_31_), .A2(n6249), .A3(n6081), .Y(N629)
         );
  AO22X1_LVT U7464 ( .A1(n3851), .A2(io_dmem_resp_bits_data[31]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[31]), .Y(n6082) );
  AO21X1_LVT U7465 ( .A1(n3856), .A2(div_io_resp_bits_data[31]), .A3(n6082), 
        .Y(n6083) );
  AO22X1_LVT U7466 ( .A1(n_T_427[671]), .A2(n3862), .A3(n3868), .A4(
        n_T_427[543]), .Y(n6087) );
  AO22X1_LVT U7467 ( .A1(n6867), .A2(n_T_427[415]), .A3(n3860), .A4(
        n_T_427[223]), .Y(n6086) );
  AO22X1_LVT U7468 ( .A1(n3837), .A2(n_T_427[479]), .A3(n3873), .A4(
        n_T_427[287]), .Y(n6085) );
  AO22X1_LVT U7469 ( .A1(n_T_427[798]), .A2(n3812), .A3(n3839), .A4(
        n_T_427[31]), .Y(n6084) );
  NOR4X1_LVT U7470 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .Y(n6088)
         );
  OA22X1_LVT U7471 ( .A1(n3099), .A2(n3596), .A3(n3878), .A4(n6088), .Y(n6090)
         );
  NAND2X0_LVT U7472 ( .A1(n_T_427[607]), .A2(n2869), .Y(n6089) );
  AO22X1_LVT U7473 ( .A1(n3921), .A2(n_T_427[1374]), .A3(n_T_427[1438]), .A4(
        n3932), .Y(n6094) );
  AO22X1_LVT U7474 ( .A1(n3931), .A2(n_T_427[1310]), .A3(n_T_427[1182]), .A4(
        n3942), .Y(n6093) );
  AO22X1_LVT U7475 ( .A1(n3941), .A2(n_T_427[1246]), .A3(n_T_427[1118]), .A4(
        n3952), .Y(n6092) );
  AO22X1_LVT U7476 ( .A1(n3951), .A2(n_T_427[990]), .A3(n_T_427[1054]), .A4(
        n3899), .Y(n6091) );
  NOR4X1_LVT U7477 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .Y(n6095)
         );
  NAND3X0_LVT U7478 ( .A1(n6097), .A2(n6096), .A3(n6095), .Y(id_rs_1[31]) );
  NAND2X0_LVT U7479 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[31]), .Y(n6101) );
  NAND2X0_LVT U7480 ( .A1(n_T_918[31]), .A2(n6899), .Y(n6100) );
  NAND2X0_LVT U7481 ( .A1(io_imem_sfence_bits_addr[31]), .A2(n6900), .Y(n6099)
         );
  NAND2X0_LVT U7482 ( .A1(n_T_635[31]), .A2(n6901), .Y(n6098) );
  NAND4X0_LVT U7483 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .Y(
        n_T_702[31]) );
  AO22X1_LVT U7484 ( .A1(n6856), .A2(io_fpu_toint_data[32]), .A3(n6855), .A4(
        n_T_918[32]), .Y(n6102) );
  AO21X1_LVT U7485 ( .A1(mem_br_target_32_), .A2(n6249), .A3(n6102), .Y(N630)
         );
  NAND2X0_LVT U7486 ( .A1(csr_io_rw_rdata[32]), .A2(n3844), .Y(n6105) );
  AOI22X1_LVT U7487 ( .A1(n3852), .A2(io_dmem_resp_bits_data[32]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[32]), .Y(n6104) );
  NAND2X0_LVT U7488 ( .A1(div_io_resp_bits_data[32]), .A2(n3858), .Y(n6103) );
  NAND3X0_LVT U7489 ( .A1(n6105), .A2(n6104), .A3(n6103), .Y(
        n_T_427__T_1136_data[32]) );
  AO22X1_LVT U7490 ( .A1(n_T_427[672]), .A2(n3862), .A3(n3865), .A4(
        n_T_427[416]), .Y(n6109) );
  AO22X1_LVT U7491 ( .A1(n3815), .A2(n_T_427[160]), .A3(n_T_427[799]), .A4(
        n3812), .Y(n6108) );
  AO22X1_LVT U7492 ( .A1(n3837), .A2(n_T_427[480]), .A3(n3866), .A4(
        n_T_427[352]), .Y(n6107) );
  AO22X1_LVT U7493 ( .A1(n_T_427[927]), .A2(n3811), .A3(n3873), .A4(
        n_T_427[288]), .Y(n6106) );
  NOR4X1_LVT U7494 ( .A1(n6109), .A2(n6108), .A3(n6107), .A4(n6106), .Y(n6110)
         );
  NAND2X0_LVT U7495 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[32]), .Y(n6114) );
  NAND2X0_LVT U7496 ( .A1(n6899), .A2(n_T_918[32]), .Y(n6113) );
  NAND2X0_LVT U7497 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[32]), .Y(n6112)
         );
  NAND2X0_LVT U7498 ( .A1(n3243), .A2(n_T_635[32]), .Y(n6111) );
  NAND4X0_LVT U7499 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .Y(
        n_T_702[32]) );
  AO22X1_LVT U7500 ( .A1(n6856), .A2(io_fpu_toint_data[33]), .A3(n6855), .A4(
        n_T_918[33]), .Y(n6115) );
  AO21X1_LVT U7501 ( .A1(mem_br_target_33_), .A2(n6249), .A3(n6115), .Y(N631)
         );
  NAND2X0_LVT U7502 ( .A1(csr_io_rw_rdata[33]), .A2(n3844), .Y(n6118) );
  AOI22X1_LVT U7503 ( .A1(n3853), .A2(io_dmem_resp_bits_data[33]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[33]), .Y(n6117) );
  NAND2X0_LVT U7504 ( .A1(div_io_resp_bits_data[33]), .A2(n3858), .Y(n6116) );
  AO22X1_LVT U7505 ( .A1(n3918), .A2(n_T_427[1376]), .A3(n_T_427[1440]), .A4(
        n3932), .Y(n6122) );
  AO22X1_LVT U7506 ( .A1(n3930), .A2(n_T_427[1312]), .A3(n_T_427[1184]), .A4(
        n3942), .Y(n6121) );
  AO22X1_LVT U7507 ( .A1(n3940), .A2(n_T_427[1248]), .A3(n_T_427[1120]), .A4(
        n3952), .Y(n6120) );
  AO22X1_LVT U7508 ( .A1(n3950), .A2(n_T_427[992]), .A3(n_T_427[1056]), .A4(
        n3899), .Y(n6119) );
  NOR4X1_LVT U7509 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .Y(n6133)
         );
  AO22X1_LVT U7510 ( .A1(n6765), .A2(n_T_427[737]), .A3(n3865), .A4(
        n_T_427[417]), .Y(n6126) );
  AO22X1_LVT U7511 ( .A1(n3869), .A2(n_T_427[545]), .A3(n_T_427[609]), .A4(
        n3795), .Y(n6125) );
  AO22X1_LVT U7512 ( .A1(n_T_427[673]), .A2(n3862), .A3(n3866), .A4(
        n_T_427[353]), .Y(n6124) );
  AO22X1_LVT U7513 ( .A1(n3813), .A2(n_T_427[800]), .A3(n_T_427[864]), .A4(
        n3874), .Y(n6123) );
  NOR4X1_LVT U7514 ( .A1(n6126), .A2(n6125), .A3(n6124), .A4(n6123), .Y(n6127)
         );
  OA22X1_LVT U7515 ( .A1(n3091), .A2(n3596), .A3(n3878), .A4(n6127), .Y(n6130)
         );
  AOI22X1_LVT U7516 ( .A1(n3911), .A2(n_T_427[481]), .A3(n_T_427[289]), .A4(
        n6774), .Y(n6129) );
  NAND2X0_LVT U7517 ( .A1(n_T_427[33]), .A2(n2879), .Y(n6128) );
  AND3X1_LVT U7518 ( .A1(n6130), .A2(n6129), .A3(n6128), .Y(n6131) );
  NAND4X0_LVT U7519 ( .A1(n6133), .A2(n6134), .A3(n6132), .A4(n6131), .Y(
        id_rs_1[33]) );
  NAND2X0_LVT U7520 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[33]), .Y(n6138) );
  NAND2X0_LVT U7521 ( .A1(n6899), .A2(n_T_918[33]), .Y(n6137) );
  NAND2X0_LVT U7522 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[33]), .Y(n6136)
         );
  NAND2X0_LVT U7523 ( .A1(n6901), .A2(n_T_635[33]), .Y(n6135) );
  NAND4X0_LVT U7524 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .Y(
        n_T_702[33]) );
  NAND2X0_LVT U7525 ( .A1(csr_io_rw_rdata[34]), .A2(n3844), .Y(n6141) );
  AOI22X1_LVT U7526 ( .A1(n3853), .A2(io_dmem_resp_bits_data[34]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[34]), .Y(n6140) );
  NAND2X0_LVT U7527 ( .A1(div_io_resp_bits_data[34]), .A2(n3858), .Y(n6139) );
  NAND3X0_LVT U7528 ( .A1(n6141), .A2(n6140), .A3(n6139), .Y(
        n_T_427__T_1136_data[34]) );
  AOI22X1_LVT U7529 ( .A1(n3816), .A2(n_T_427[162]), .A3(n_T_427[801]), .A4(
        n3812), .Y(n6145) );
  OA22X1_LVT U7530 ( .A1(n6767), .A2(n3527), .A3(n3141), .A4(n3805), .Y(n6144)
         );
  AOI22X1_LVT U7531 ( .A1(n_T_427[674]), .A2(n3861), .A3(n3868), .A4(
        n_T_427[546]), .Y(n6143) );
  AOI22X1_LVT U7532 ( .A1(n_T_427[929]), .A2(n6794), .A3(n3875), .A4(
        n_T_427[865]), .Y(n6142) );
  NAND4X0_LVT U7533 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .Y(n6146) );
  AO22X1_LVT U7534 ( .A1(n3924), .A2(n_T_427[1505]), .A3(n_T_427[1377]), .A4(
        n3919), .Y(n6150) );
  AO22X1_LVT U7535 ( .A1(n3934), .A2(n_T_427[1441]), .A3(n_T_427[1313]), .A4(
        n3929), .Y(n6149) );
  AO22X1_LVT U7536 ( .A1(n3944), .A2(n_T_427[1185]), .A3(n_T_427[1249]), .A4(
        n3939), .Y(n6148) );
  AO22X1_LVT U7537 ( .A1(n3954), .A2(n_T_427[1121]), .A3(n_T_427[993]), .A4(
        n3949), .Y(n6147) );
  NOR4X1_LVT U7538 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .Y(n6157)
         );
  AO22X1_LVT U7539 ( .A1(n2824), .A2(n_T_427[482]), .A3(n_T_427[98]), .A4(
        n2871), .Y(n6154) );
  AO22X1_LVT U7540 ( .A1(n3901), .A2(n_T_427[1057]), .A3(n_T_427[226]), .A4(
        n3807), .Y(n6153) );
  AO22X1_LVT U7541 ( .A1(n1919), .A2(n_T_427[354]), .A3(n_T_427[34]), .A4(
        n3913), .Y(n6152) );
  AO22X1_LVT U7542 ( .A1(n3916), .A2(n_T_427[610]), .A3(n_T_427[290]), .A4(
        n3810), .Y(n6151) );
  NOR4X1_LVT U7543 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .Y(n6156)
         );
  NAND2X0_LVT U7544 ( .A1(n3957), .A2(n4411), .Y(n6155) );
  NAND4X0_LVT U7545 ( .A1(n6157), .A2(n6158), .A3(n6156), .A4(n6155), .Y(
        id_rs_1[34]) );
  NAND2X0_LVT U7546 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[34]), .Y(n6162) );
  NAND2X0_LVT U7547 ( .A1(n6899), .A2(n_T_918[34]), .Y(n6161) );
  NAND2X0_LVT U7548 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[34]), .Y(n6160)
         );
  NAND2X0_LVT U7549 ( .A1(n3243), .A2(n_T_635[34]), .Y(n6159) );
  NAND4X0_LVT U7550 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .Y(
        n_T_702[34]) );
  AO22X1_LVT U7551 ( .A1(n6856), .A2(io_fpu_toint_data[35]), .A3(n6855), .A4(
        n_T_918[35]), .Y(n6163) );
  AO21X1_LVT U7552 ( .A1(mem_br_target_35_), .A2(n6249), .A3(n6163), .Y(N633)
         );
  NAND2X0_LVT U7553 ( .A1(csr_io_rw_rdata[35]), .A2(n3845), .Y(n6166) );
  AOI22X1_LVT U7554 ( .A1(n3853), .A2(io_dmem_resp_bits_data[35]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[35]), .Y(n6165) );
  NAND2X0_LVT U7555 ( .A1(div_io_resp_bits_data[35]), .A2(n3858), .Y(n6164) );
  AO22X1_LVT U7556 ( .A1(n3920), .A2(n_T_427[1378]), .A3(n_T_427[1442]), .A4(
        n3932), .Y(n6170) );
  AO22X1_LVT U7557 ( .A1(n3931), .A2(n_T_427[1314]), .A3(n_T_427[1186]), .A4(
        n3942), .Y(n6169) );
  AO22X1_LVT U7558 ( .A1(n3938), .A2(n_T_427[1250]), .A3(n_T_427[1122]), .A4(
        n3952), .Y(n6168) );
  AO22X1_LVT U7559 ( .A1(n3948), .A2(n_T_427[994]), .A3(n_T_427[1058]), .A4(
        n3899), .Y(n6167) );
  NOR4X1_LVT U7560 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .Y(n6183)
         );
  AO22X1_LVT U7561 ( .A1(n3835), .A2(n_T_427[419]), .A3(n_T_427[611]), .A4(
        n2870), .Y(n6172) );
  AO22X1_LVT U7562 ( .A1(n3806), .A2(n_T_427[227]), .A3(n_T_427[738]), .A4(
        n3903), .Y(n6171) );
  AOI22X1_LVT U7563 ( .A1(n6886), .A2(n_T_427[163]), .A3(n_T_427[675]), .A4(
        n2829), .Y(n6180) );
  NAND2X0_LVT U7564 ( .A1(n_T_427[291]), .A2(n3809), .Y(n6179) );
  AO22X1_LVT U7565 ( .A1(n_T_427[930]), .A2(n3811), .A3(n3875), .A4(
        n_T_427[866]), .Y(n6176) );
  AO22X1_LVT U7566 ( .A1(n3870), .A2(n_T_427[547]), .A3(n_T_427[483]), .A4(
        n3836), .Y(n6175) );
  AO22X1_LVT U7567 ( .A1(n_T_427[802]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[35]), .Y(n6174) );
  AO22X1_LVT U7568 ( .A1(n6866), .A2(n_T_427[99]), .A3(n3866), .A4(
        n_T_427[355]), .Y(n6173) );
  NOR4X1_LVT U7569 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .Y(n6177)
         );
  OA22X1_LVT U7570 ( .A1(n3183), .A2(n3596), .A3(n3878), .A4(n6177), .Y(n6178)
         );
  AND3X1_LVT U7571 ( .A1(n6180), .A2(n6179), .A3(n6178), .Y(n6181) );
  NAND4X0_LVT U7572 ( .A1(n6183), .A2(n6184), .A3(n6182), .A4(n6181), .Y(
        id_rs_1[35]) );
  NAND2X0_LVT U7573 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[35]), .Y(n6188) );
  NAND2X0_LVT U7574 ( .A1(n6899), .A2(n_T_918[35]), .Y(n6187) );
  NAND2X0_LVT U7575 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[35]), .Y(n6186)
         );
  NAND2X0_LVT U7576 ( .A1(n3243), .A2(n_T_635[35]), .Y(n6185) );
  NAND4X0_LVT U7577 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .Y(
        n_T_702[35]) );
  AO22X1_LVT U7578 ( .A1(n3851), .A2(io_dmem_resp_bits_data[36]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[36]), .Y(n6189) );
  AO21X1_LVT U7579 ( .A1(n3856), .A2(div_io_resp_bits_data[36]), .A3(n6189), 
        .Y(n6190) );
  AO21X1_LVT U7580 ( .A1(n3843), .A2(csr_io_rw_rdata[36]), .A3(n6190), .Y(
        n_T_427__T_1136_data[36]) );
  AO22X1_LVT U7581 ( .A1(n3916), .A2(n_T_427[612]), .A3(n_T_427[164]), .A4(
        n3909), .Y(n6192) );
  AO22X1_LVT U7582 ( .A1(n2828), .A2(n_T_427[292]), .A3(n_T_427[676]), .A4(
        n6812), .Y(n6191) );
  NOR2X0_LVT U7583 ( .A1(n6192), .A2(n6191), .Y(n6202) );
  AO22X1_LVT U7584 ( .A1(n3869), .A2(n_T_427[548]), .A3(n_T_427[867]), .A4(
        n3874), .Y(n6196) );
  AO22X1_LVT U7585 ( .A1(n6867), .A2(n_T_427[420]), .A3(n6866), .A4(
        n_T_427[100]), .Y(n6195) );
  AO22X1_LVT U7586 ( .A1(n3860), .A2(n_T_427[228]), .A3(n3866), .A4(
        n_T_427[356]), .Y(n6194) );
  AO22X1_LVT U7587 ( .A1(n_T_427[803]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[36]), .Y(n6193) );
  NOR4X1_LVT U7588 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .Y(n6197)
         );
  OA22X1_LVT U7589 ( .A1(n3549), .A2(n3881), .A3(n3878), .A4(n6197), .Y(n6200)
         );
  OA22X1_LVT U7590 ( .A1(n3145), .A2(n3803), .A3(n3497), .A4(n3800), .Y(n6199)
         );
  NAND2X0_LVT U7591 ( .A1(n4416), .A2(n3959), .Y(n6198) );
  AND3X1_LVT U7592 ( .A1(n6200), .A2(n6199), .A3(n6198), .Y(n6201) );
  NAND4X0_LVT U7593 ( .A1(n6203), .A2(n6204), .A3(n6202), .A4(n6201), .Y(
        id_rs_1[36]) );
  NAND2X0_LVT U7594 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[36]), .Y(n6208) );
  NAND2X0_LVT U7595 ( .A1(n6899), .A2(n_T_918[36]), .Y(n6207) );
  NAND2X0_LVT U7596 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[36]), .Y(n6206)
         );
  NAND2X0_LVT U7597 ( .A1(n3243), .A2(n_T_635[36]), .Y(n6205) );
  NAND4X0_LVT U7598 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .Y(
        n_T_702[36]) );
  NAND2X0_LVT U7599 ( .A1(csr_io_rw_rdata[37]), .A2(n3845), .Y(n6211) );
  AOI22X1_LVT U7600 ( .A1(n3853), .A2(io_dmem_resp_bits_data[37]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[37]), .Y(n6210) );
  NAND2X0_LVT U7601 ( .A1(div_io_resp_bits_data[37]), .A2(n3858), .Y(n6209) );
  NAND3X0_LVT U7602 ( .A1(n6211), .A2(n6210), .A3(n6209), .Y(
        n_T_427__T_1136_data[37]) );
  AO22X1_LVT U7603 ( .A1(n3910), .A2(n_T_427[485]), .A3(n_T_427[165]), .A4(
        n2862), .Y(n6213) );
  AO22X1_LVT U7604 ( .A1(n3818), .A2(n_T_427[549]), .A3(n_T_427[868]), .A4(
        n3823), .Y(n6212) );
  NOR2X0_LVT U7605 ( .A1(n6213), .A2(n6212), .Y(n6223) );
  AO22X1_LVT U7606 ( .A1(n_T_427[677]), .A2(n3861), .A3(n3865), .A4(
        n_T_427[421]), .Y(n6217) );
  AO22X1_LVT U7607 ( .A1(n_T_427[613]), .A2(n3797), .A3(n3866), .A4(
        n_T_427[357]), .Y(n6216) );
  AO22X1_LVT U7608 ( .A1(n_T_427[932]), .A2(n3811), .A3(n3873), .A4(
        n_T_427[293]), .Y(n6215) );
  AO22X1_LVT U7609 ( .A1(n_T_427[804]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[37]), .Y(n6214) );
  NOR4X1_LVT U7610 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .Y(n6218)
         );
  OA22X1_LVT U7611 ( .A1(n3550), .A2(n3881), .A3(n3878), .A4(n6218), .Y(n6221)
         );
  OA22X1_LVT U7612 ( .A1(n3146), .A2(n3803), .A3(n3498), .A4(n3800), .Y(n6220)
         );
  NAND2X0_LVT U7613 ( .A1(n3957), .A2(n4419), .Y(n6219) );
  AND3X1_LVT U7614 ( .A1(n6221), .A2(n6220), .A3(n6219), .Y(n6222) );
  NAND4X0_LVT U7615 ( .A1(n6224), .A2(n6225), .A3(n6223), .A4(n6222), .Y(
        id_rs_1[37]) );
  NAND2X0_LVT U7616 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[37]), .Y(n6229) );
  NAND2X0_LVT U7617 ( .A1(n6899), .A2(n_T_918[37]), .Y(n6228) );
  NAND2X0_LVT U7618 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[37]), .Y(n6227)
         );
  NAND2X0_LVT U7619 ( .A1(n6901), .A2(n_T_635[37]), .Y(n6226) );
  NAND4X0_LVT U7620 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .Y(
        n_T_702[37]) );
  AO22X1_LVT U7621 ( .A1(n6856), .A2(io_fpu_toint_data[38]), .A3(n6855), .A4(
        n_T_918[38]), .Y(n6230) );
  AO21X1_LVT U7622 ( .A1(mem_br_target_38_), .A2(n6249), .A3(n6230), .Y(N636)
         );
  AO22X1_LVT U7623 ( .A1(n3851), .A2(io_dmem_resp_bits_data[38]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[38]), .Y(n6231) );
  AO21X1_LVT U7624 ( .A1(n3856), .A2(div_io_resp_bits_data[38]), .A3(n6231), 
        .Y(n6232) );
  AO22X1_LVT U7625 ( .A1(n3806), .A2(n_T_427[230]), .A3(n_T_427[166]), .A4(
        n2862), .Y(n6244) );
  AO22X1_LVT U7626 ( .A1(n2869), .A2(n_T_427[614]), .A3(n_T_427[102]), .A4(
        n3832), .Y(n6243) );
  AO22X1_LVT U7627 ( .A1(n3913), .A2(n_T_427[38]), .A3(n_T_427[294]), .A4(
        n3809), .Y(n6242) );
  AO22X1_LVT U7628 ( .A1(n_T_427[933]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[486]), .Y(n6236) );
  AO22X1_LVT U7629 ( .A1(n6765), .A2(n_T_427[741]), .A3(n3865), .A4(
        n_T_427[422]), .Y(n6235) );
  AO22X1_LVT U7630 ( .A1(n_T_427[678]), .A2(n3861), .A3(n3866), .A4(
        n_T_427[358]), .Y(n6234) );
  AO22X1_LVT U7631 ( .A1(n3813), .A2(n_T_427[805]), .A3(n_T_427[869]), .A4(
        n3874), .Y(n6233) );
  NOR4X1_LVT U7632 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .Y(n6237)
         );
  OA22X1_LVT U7633 ( .A1(n3098), .A2(n3596), .A3(n3877), .A4(n6237), .Y(n6240)
         );
  NAND2X0_LVT U7634 ( .A1(n_T_427[550]), .A2(n2850), .Y(n6239) );
  NAND2X0_LVT U7635 ( .A1(n6240), .A2(n6239), .Y(n6241) );
  NAND2X0_LVT U7636 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[38]), .Y(n6248) );
  NAND2X0_LVT U7637 ( .A1(n6899), .A2(n_T_918[38]), .Y(n6247) );
  NAND2X0_LVT U7638 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[38]), .Y(n6246)
         );
  NAND2X0_LVT U7639 ( .A1(n3243), .A2(n_T_635[38]), .Y(n6245) );
  NAND4X0_LVT U7640 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .Y(
        n_T_702[38]) );
  AOI22X1_LVT U7641 ( .A1(n6856), .A2(io_fpu_toint_data[39]), .A3(n6855), .A4(
        n_T_918[39]), .Y(n6250) );
  NAND2X0_LVT U7642 ( .A1(n6857), .A2(n6250), .Y(N637) );
  NAND2X0_LVT U7643 ( .A1(csr_io_rw_rdata[39]), .A2(n3845), .Y(n6253) );
  AOI22X1_LVT U7644 ( .A1(n3853), .A2(io_dmem_resp_bits_data[39]), .A3(n3846), 
        .A4(n_T_1165[39]), .Y(n6252) );
  NAND2X0_LVT U7645 ( .A1(div_io_resp_bits_data[39]), .A2(n3858), .Y(n6251) );
  NAND3X0_LVT U7646 ( .A1(n6253), .A2(n6252), .A3(n6251), .Y(
        n_T_427__T_1136_data[39]) );
  AOI22X1_LVT U7647 ( .A1(n3870), .A2(n_T_427[551]), .A3(n_T_427[615]), .A4(
        n3795), .Y(n6257) );
  AOI22X1_LVT U7648 ( .A1(n6871), .A2(n_T_427[870]), .A3(n6838), .A4(
        n_T_427[39]), .Y(n6256) );
  AOI22X1_LVT U7649 ( .A1(n3865), .A2(n_T_427[423]), .A3(n_T_427[742]), .A4(
        n3804), .Y(n6255) );
  OA22X1_LVT U7650 ( .A1(n3523), .A2(n6423), .A3(n3179), .A4(n3083), .Y(n6254)
         );
  NAND4X0_LVT U7651 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .Y(n6258) );
  AO22X1_LVT U7652 ( .A1(n3925), .A2(n_T_427[1510]), .A3(n_T_427[1382]), .A4(
        n3919), .Y(n6262) );
  AO22X1_LVT U7653 ( .A1(n3935), .A2(n_T_427[1446]), .A3(n_T_427[1318]), .A4(
        n3929), .Y(n6261) );
  AO22X1_LVT U7654 ( .A1(n3945), .A2(n_T_427[1190]), .A3(n_T_427[1254]), .A4(
        n3939), .Y(n6260) );
  AO22X1_LVT U7655 ( .A1(n3955), .A2(n_T_427[1126]), .A3(n_T_427[998]), .A4(
        n3949), .Y(n6259) );
  NOR4X1_LVT U7656 ( .A1(n6262), .A2(n6261), .A3(n6260), .A4(n6259), .Y(n6269)
         );
  AO22X1_LVT U7657 ( .A1(n2860), .A2(n_T_427[806]), .A3(n_T_427[103]), .A4(
        n3832), .Y(n6266) );
  AO22X1_LVT U7658 ( .A1(n3901), .A2(n_T_427[1062]), .A3(n_T_427[934]), .A4(
        n3895), .Y(n6265) );
  AO22X1_LVT U7659 ( .A1(n3910), .A2(n_T_427[487]), .A3(n_T_427[167]), .A4(
        n2863), .Y(n6264) );
  AO22X1_LVT U7660 ( .A1(n2857), .A2(n_T_427[359]), .A3(n_T_427[295]), .A4(
        n3809), .Y(n6263) );
  NOR4X1_LVT U7661 ( .A1(n6266), .A2(n6265), .A3(n6264), .A4(n6263), .Y(n6268)
         );
  NAND2X0_LVT U7662 ( .A1(n3957), .A2(n4424), .Y(n6267) );
  NAND4X0_LVT U7663 ( .A1(n6269), .A2(n6270), .A3(n6268), .A4(n6267), .Y(
        id_rs_1[39]) );
  NAND2X0_LVT U7664 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[39]), .Y(n6274) );
  NAND2X0_LVT U7665 ( .A1(n6899), .A2(n_T_918[39]), .Y(n6273) );
  NAND2X0_LVT U7666 ( .A1(n6900), .A2(n_T_1165[39]), .Y(n6272) );
  NAND2X0_LVT U7667 ( .A1(n6901), .A2(n_T_635[39]), .Y(n6271) );
  NAND4X0_LVT U7668 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6271), .Y(
        n_T_702[39]) );
  AOI22X1_LVT U7669 ( .A1(n6856), .A2(io_fpu_toint_data[40]), .A3(n6855), .A4(
        n_T_918[40]), .Y(n6275) );
  NAND2X0_LVT U7670 ( .A1(n6857), .A2(n6275), .Y(N638) );
  NAND2X0_LVT U7671 ( .A1(csr_io_rw_rdata[40]), .A2(n3845), .Y(n6278) );
  AOI22X1_LVT U7672 ( .A1(n3853), .A2(io_dmem_resp_bits_data[40]), .A3(n3846), 
        .A4(n_T_1165[40]), .Y(n6277) );
  NAND2X0_LVT U7673 ( .A1(div_io_resp_bits_data[40]), .A2(n3858), .Y(n6276) );
  NAND3X0_LVT U7674 ( .A1(n6278), .A2(n6277), .A3(n6276), .Y(
        n_T_427__T_1136_data[40]) );
  AO22X1_LVT U7675 ( .A1(n2861), .A2(n_T_427[807]), .A3(n_T_427[168]), .A4(
        n2863), .Y(n6280) );
  AO22X1_LVT U7676 ( .A1(n3817), .A2(n_T_427[360]), .A3(n_T_427[680]), .A4(
        n6812), .Y(n6279) );
  AO22X1_LVT U7677 ( .A1(n6765), .A2(n_T_427[743]), .A3(n3865), .A4(
        n_T_427[424]), .Y(n6284) );
  AO22X1_LVT U7678 ( .A1(n3869), .A2(n_T_427[552]), .A3(n_T_427[616]), .A4(
        n3795), .Y(n6283) );
  AO22X1_LVT U7679 ( .A1(n3837), .A2(n_T_427[488]), .A3(n3873), .A4(
        n_T_427[296]), .Y(n6282) );
  AO22X1_LVT U7680 ( .A1(n_T_427[871]), .A2(n6871), .A3(n3839), .A4(
        n_T_427[40]), .Y(n6281) );
  NOR4X1_LVT U7681 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .Y(n6285)
         );
  OA22X1_LVT U7682 ( .A1(n3551), .A2(n3881), .A3(n3877), .A4(n6285), .Y(n6288)
         );
  NAND2X0_LVT U7683 ( .A1(n3958), .A2(n4427), .Y(n6287) );
  OA22X1_LVT U7684 ( .A1(n3147), .A2(n3803), .A3(n3499), .A4(n3800), .Y(n6286)
         );
  AND3X1_LVT U7685 ( .A1(n6288), .A2(n6287), .A3(n6286), .Y(n6289) );
  NAND4X0_LVT U7686 ( .A1(n6291), .A2(n6292), .A3(n6290), .A4(n6289), .Y(
        id_rs_1[40]) );
  NAND2X0_LVT U7687 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[40]), .Y(n6296) );
  NAND2X0_LVT U7688 ( .A1(n6899), .A2(n_T_918[40]), .Y(n6295) );
  NAND2X0_LVT U7689 ( .A1(n6900), .A2(n_T_1165[40]), .Y(n6294) );
  NAND2X0_LVT U7690 ( .A1(n3243), .A2(n_T_635[40]), .Y(n6293) );
  NAND4X0_LVT U7691 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .Y(
        n_T_702[40]) );
  AOI22X1_LVT U7692 ( .A1(n6856), .A2(io_fpu_toint_data[41]), .A3(n6855), .A4(
        n_T_918[41]), .Y(n6297) );
  NAND2X0_LVT U7693 ( .A1(n6857), .A2(n6297), .Y(N639) );
  AO22X1_LVT U7694 ( .A1(n3851), .A2(io_dmem_resp_bits_data[41]), .A3(n3848), 
        .A4(n_T_1165[41]), .Y(n6298) );
  AO21X1_LVT U7695 ( .A1(n3856), .A2(div_io_resp_bits_data[41]), .A3(n6298), 
        .Y(n6299) );
  AO21X1_LVT U7696 ( .A1(n3842), .A2(csr_io_rw_rdata[41]), .A3(n6299), .Y(
        n_T_427__T_1136_data[41]) );
  AO22X1_LVT U7697 ( .A1(n3945), .A2(n_T_427[1192]), .A3(n_T_427[1256]), .A4(
        n3939), .Y(n6303) );
  AO22X1_LVT U7698 ( .A1(n3955), .A2(n_T_427[1128]), .A3(n_T_427[1000]), .A4(
        n3949), .Y(n6302) );
  AO22X1_LVT U7699 ( .A1(n3901), .A2(n_T_427[1064]), .A3(n_T_427[233]), .A4(
        n6773), .Y(n6301) );
  AO22X1_LVT U7700 ( .A1(n2861), .A2(n_T_427[808]), .A3(n_T_427[489]), .A4(
        n3911), .Y(n6300) );
  NOR4X1_LVT U7701 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .Y(n6316)
         );
  AO22X1_LVT U7702 ( .A1(n2833), .A2(n_T_427[872]), .A3(n_T_427[169]), .A4(
        n2862), .Y(n6305) );
  AO22X1_LVT U7703 ( .A1(n3809), .A2(n_T_427[297]), .A3(n_T_427[681]), .A4(
        n3821), .Y(n6304) );
  NOR2X0_LVT U7704 ( .A1(n6305), .A2(n6304), .Y(n6315) );
  AO22X1_LVT U7705 ( .A1(n3869), .A2(n_T_427[553]), .A3(n_T_427[617]), .A4(
        n3795), .Y(n6309) );
  AO22X1_LVT U7706 ( .A1(n_T_427[744]), .A2(n3804), .A3(n6866), .A4(
        n_T_427[105]), .Y(n6308) );
  AO22X1_LVT U7707 ( .A1(n6867), .A2(n_T_427[425]), .A3(n3866), .A4(
        n_T_427[361]), .Y(n6307) );
  AO22X1_LVT U7708 ( .A1(n_T_427[936]), .A2(n6794), .A3(n3839), .A4(
        n_T_427[41]), .Y(n6306) );
  NOR4X1_LVT U7709 ( .A1(n6309), .A2(n6308), .A3(n6307), .A4(n6306), .Y(n6310)
         );
  OA22X1_LVT U7710 ( .A1(n3552), .A2(n3881), .A3(n1993), .A4(n6310), .Y(n6313)
         );
  OA22X1_LVT U7711 ( .A1(n3148), .A2(n3803), .A3(n3500), .A4(n3799), .Y(n6312)
         );
  NAND2X0_LVT U7712 ( .A1(n4430), .A2(n3959), .Y(n6311) );
  AND3X1_LVT U7713 ( .A1(n6313), .A2(n6312), .A3(n6311), .Y(n6314) );
  NAND4X0_LVT U7714 ( .A1(n6316), .A2(n6317), .A3(n6315), .A4(n6314), .Y(
        id_rs_1[41]) );
  NAND2X0_LVT U7715 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[41]), .Y(n6321) );
  NAND2X0_LVT U7716 ( .A1(n6899), .A2(n_T_918[41]), .Y(n6320) );
  NAND2X0_LVT U7717 ( .A1(n6900), .A2(n_T_1165[41]), .Y(n6319) );
  NAND2X0_LVT U7718 ( .A1(n6901), .A2(n_T_635[41]), .Y(n6318) );
  NAND4X0_LVT U7719 ( .A1(n6321), .A2(n6320), .A3(n6319), .A4(n6318), .Y(
        n_T_702[41]) );
  AOI22X1_LVT U7720 ( .A1(n6856), .A2(io_fpu_toint_data[42]), .A3(n6855), .A4(
        n_T_918[42]), .Y(n6322) );
  NAND2X0_LVT U7721 ( .A1(n6857), .A2(n6322), .Y(N640) );
  AO22X1_LVT U7722 ( .A1(n3851), .A2(io_dmem_resp_bits_data[42]), .A3(n3848), 
        .A4(n_T_1165[42]), .Y(n6323) );
  AO21X1_LVT U7723 ( .A1(n3857), .A2(div_io_resp_bits_data[42]), .A3(n6323), 
        .Y(n6324) );
  AO21X1_LVT U7724 ( .A1(n3842), .A2(csr_io_rw_rdata[42]), .A3(n6324), .Y(
        n_T_427__T_1136_data[42]) );
  AO22X1_LVT U7725 ( .A1(n3945), .A2(n_T_427[1193]), .A3(n_T_427[1257]), .A4(
        n3940), .Y(n6328) );
  AO22X1_LVT U7726 ( .A1(n3955), .A2(n_T_427[1129]), .A3(n_T_427[1001]), .A4(
        n3950), .Y(n6327) );
  AO22X1_LVT U7727 ( .A1(n3901), .A2(n_T_427[1065]), .A3(n_T_427[234]), .A4(
        n6773), .Y(n6326) );
  AO22X1_LVT U7728 ( .A1(n2865), .A2(n_T_427[426]), .A3(n_T_427[745]), .A4(
        n3904), .Y(n6325) );
  NOR4X1_LVT U7729 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .Y(n6341)
         );
  AO22X1_LVT U7730 ( .A1(n3912), .A2(n_T_427[490]), .A3(n_T_427[170]), .A4(
        n3908), .Y(n6330) );
  AO22X1_LVT U7731 ( .A1(n2833), .A2(n_T_427[873]), .A3(n_T_427[298]), .A4(
        n3809), .Y(n6329) );
  AO22X1_LVT U7732 ( .A1(n_T_427[937]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[618]), .Y(n6334) );
  AO22X1_LVT U7733 ( .A1(n_T_427[682]), .A2(n3861), .A3(n6866), .A4(
        n_T_427[106]), .Y(n6333) );
  AO22X1_LVT U7734 ( .A1(n_T_427[554]), .A2(n3869), .A3(n3866), .A4(
        n_T_427[362]), .Y(n6332) );
  AO22X1_LVT U7735 ( .A1(n_T_427[809]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[42]), .Y(n6331) );
  NOR4X1_LVT U7736 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .Y(n6335)
         );
  OA22X1_LVT U7737 ( .A1(n3553), .A2(n3881), .A3(n1993), .A4(n6335), .Y(n6338)
         );
  OA22X1_LVT U7738 ( .A1(n3149), .A2(n3803), .A3(n3501), .A4(n3799), .Y(n6337)
         );
  NAND2X0_LVT U7739 ( .A1(n4433), .A2(n3959), .Y(n6336) );
  AND3X1_LVT U7740 ( .A1(n6338), .A2(n6337), .A3(n6336), .Y(n6339) );
  NAND4X0_LVT U7741 ( .A1(n6341), .A2(n6342), .A3(n6340), .A4(n6339), .Y(
        id_rs_1[42]) );
  NAND2X0_LVT U7742 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[42]), .Y(n6346) );
  NAND2X0_LVT U7743 ( .A1(n6899), .A2(n_T_918[42]), .Y(n6345) );
  NAND2X0_LVT U7744 ( .A1(n6900), .A2(n_T_1165[42]), .Y(n6344) );
  NAND2X0_LVT U7745 ( .A1(n3243), .A2(n_T_635[42]), .Y(n6343) );
  NAND4X0_LVT U7746 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .Y(
        n_T_702[42]) );
  AOI22X1_LVT U7747 ( .A1(n6856), .A2(io_fpu_toint_data[43]), .A3(n6855), .A4(
        n_T_918[43]), .Y(n6347) );
  NAND2X0_LVT U7748 ( .A1(n6857), .A2(n6347), .Y(N641) );
  AO22X1_LVT U7749 ( .A1(n3851), .A2(io_dmem_resp_bits_data[43]), .A3(n3848), 
        .A4(n_T_1165[43]), .Y(n6348) );
  AO21X1_LVT U7750 ( .A1(n3857), .A2(div_io_resp_bits_data[43]), .A3(n6348), 
        .Y(n6349) );
  AO21X1_LVT U7751 ( .A1(n3842), .A2(csr_io_rw_rdata[43]), .A3(n6349), .Y(
        n_T_427__T_1136_data[43]) );
  AO22X1_LVT U7752 ( .A1(n3915), .A2(n_T_427[619]), .A3(n_T_427[171]), .A4(
        n3909), .Y(n6351) );
  AO22X1_LVT U7753 ( .A1(n3810), .A2(n_T_427[299]), .A3(n_T_427[683]), .A4(
        n2829), .Y(n6350) );
  NOR2X0_LVT U7754 ( .A1(n6351), .A2(n6350), .Y(n6361) );
  AO22X1_LVT U7755 ( .A1(n3869), .A2(n_T_427[555]), .A3(n_T_427[491]), .A4(
        n3836), .Y(n6355) );
  AO22X1_LVT U7756 ( .A1(n6867), .A2(n_T_427[427]), .A3(n6866), .A4(
        n_T_427[107]), .Y(n6354) );
  AO22X1_LVT U7757 ( .A1(n3860), .A2(n_T_427[235]), .A3(n3866), .A4(
        n_T_427[363]), .Y(n6353) );
  AO22X1_LVT U7758 ( .A1(n_T_427[874]), .A2(n6871), .A3(n3839), .A4(
        n_T_427[43]), .Y(n6352) );
  NOR4X1_LVT U7759 ( .A1(n6355), .A2(n6354), .A3(n6353), .A4(n6352), .Y(n6356)
         );
  OA22X1_LVT U7760 ( .A1(n3554), .A2(n3881), .A3(n3877), .A4(n6356), .Y(n6359)
         );
  OA22X1_LVT U7761 ( .A1(n3150), .A2(n3803), .A3(n3502), .A4(n3799), .Y(n6358)
         );
  NAND2X0_LVT U7762 ( .A1(n4436), .A2(n3959), .Y(n6357) );
  AND3X1_LVT U7763 ( .A1(n6359), .A2(n6358), .A3(n6357), .Y(n6360) );
  NAND4X0_LVT U7764 ( .A1(n6362), .A2(n6363), .A3(n6361), .A4(n6360), .Y(
        id_rs_1[43]) );
  NAND2X0_LVT U7765 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[43]), .Y(n6367) );
  NAND2X0_LVT U7766 ( .A1(n6899), .A2(n_T_918[43]), .Y(n6366) );
  NAND2X0_LVT U7767 ( .A1(n6900), .A2(n_T_1165[43]), .Y(n6365) );
  NAND2X0_LVT U7768 ( .A1(n3243), .A2(n_T_635[43]), .Y(n6364) );
  NAND4X0_LVT U7769 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .Y(
        n_T_702[43]) );
  AOI22X1_LVT U7770 ( .A1(n6856), .A2(io_fpu_toint_data[44]), .A3(n6855), .A4(
        n_T_918[44]), .Y(n6368) );
  NAND2X0_LVT U7771 ( .A1(n6857), .A2(n6368), .Y(N642) );
  NAND2X0_LVT U7772 ( .A1(csr_io_rw_rdata[44]), .A2(n3845), .Y(n6371) );
  AOI22X1_LVT U7773 ( .A1(n3853), .A2(io_dmem_resp_bits_data[44]), .A3(n3846), 
        .A4(n_T_1165[44]), .Y(n6370) );
  NAND2X0_LVT U7774 ( .A1(div_io_resp_bits_data[44]), .A2(n3858), .Y(n6369) );
  NAND3X0_LVT U7775 ( .A1(n6371), .A2(n6370), .A3(n6369), .Y(
        n_T_427__T_1136_data[44]) );
  AOI22X1_LVT U7776 ( .A1(n3797), .A2(n_T_427[620]), .A3(n3867), .A4(
        n_T_427[364]), .Y(n6375) );
  AOI22X1_LVT U7777 ( .A1(n6871), .A2(n_T_427[875]), .A3(n3871), .A4(
        n_T_427[300]), .Y(n6374) );
  AOI22X1_LVT U7778 ( .A1(n6765), .A2(n_T_427[747]), .A3(n3864), .A4(
        n_T_427[108]), .Y(n6373) );
  AOI22X1_LVT U7779 ( .A1(n3863), .A2(n_T_427[684]), .A3(n3865), .A4(
        n_T_427[428]), .Y(n6372) );
  NAND4X0_LVT U7780 ( .A1(n6375), .A2(n6374), .A3(n6373), .A4(n6372), .Y(n6376) );
  AO22X1_LVT U7781 ( .A1(n3901), .A2(n_T_427[1067]), .A3(n_T_427[236]), .A4(
        n3807), .Y(n6380) );
  AO22X1_LVT U7782 ( .A1(n2860), .A2(n_T_427[811]), .A3(n_T_427[939]), .A4(
        n3895), .Y(n6379) );
  AO22X1_LVT U7783 ( .A1(n3912), .A2(n_T_427[492]), .A3(n_T_427[172]), .A4(
        n3909), .Y(n6378) );
  AO22X1_LVT U7784 ( .A1(n3818), .A2(n_T_427[556]), .A3(n_T_427[44]), .A4(
        n3914), .Y(n6377) );
  NOR4X1_LVT U7785 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .Y(n6387)
         );
  AO22X1_LVT U7786 ( .A1(n3925), .A2(n_T_427[1515]), .A3(n_T_427[1387]), .A4(
        n3920), .Y(n6384) );
  AO22X1_LVT U7787 ( .A1(n3935), .A2(n_T_427[1451]), .A3(n_T_427[1323]), .A4(
        n3930), .Y(n6383) );
  AO22X1_LVT U7788 ( .A1(n3945), .A2(n_T_427[1195]), .A3(n_T_427[1259]), .A4(
        n3940), .Y(n6382) );
  AO22X1_LVT U7789 ( .A1(n3955), .A2(n_T_427[1131]), .A3(n_T_427[1003]), .A4(
        n3950), .Y(n6381) );
  NOR4X1_LVT U7790 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .Y(n6386)
         );
  NAND2X0_LVT U7791 ( .A1(n3957), .A2(n4439), .Y(n6385) );
  NAND4X0_LVT U7792 ( .A1(n6387), .A2(n6388), .A3(n6386), .A4(n6385), .Y(
        id_rs_1[44]) );
  NAND2X0_LVT U7793 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[44]), .Y(n6392) );
  NAND2X0_LVT U7794 ( .A1(n6899), .A2(n_T_918[44]), .Y(n6391) );
  NAND2X0_LVT U7795 ( .A1(n6900), .A2(n_T_1165[44]), .Y(n6390) );
  NAND2X0_LVT U7796 ( .A1(n6901), .A2(n_T_635[44]), .Y(n6389) );
  NAND4X0_LVT U7797 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .Y(
        n_T_702[44]) );
  AOI22X1_LVT U7798 ( .A1(n6856), .A2(io_fpu_toint_data[45]), .A3(n6855), .A4(
        n_T_918[45]), .Y(n6393) );
  NAND2X0_LVT U7799 ( .A1(n6857), .A2(n6393), .Y(N643) );
  AO22X1_LVT U7800 ( .A1(n3851), .A2(io_dmem_resp_bits_data[45]), .A3(n3848), 
        .A4(n_T_1165[45]), .Y(n6394) );
  AO21X1_LVT U7801 ( .A1(n3857), .A2(div_io_resp_bits_data[45]), .A3(n6394), 
        .Y(n6395) );
  AO21X1_LVT U7802 ( .A1(n3842), .A2(csr_io_rw_rdata[45]), .A3(n6395), .Y(
        n_T_427__T_1136_data[45]) );
  AO22X1_LVT U7803 ( .A1(n3818), .A2(n_T_427[557]), .A3(n_T_427[45]), .A4(
        n2826), .Y(n6397) );
  AO22X1_LVT U7804 ( .A1(n3822), .A2(n_T_427[876]), .A3(n_T_427[685]), .A4(
        n3820), .Y(n6396) );
  NOR2X0_LVT U7805 ( .A1(n6397), .A2(n6396), .Y(n6407) );
  AO22X1_LVT U7806 ( .A1(n3815), .A2(n_T_427[173]), .A3(n_T_427[812]), .A4(
        n3812), .Y(n6401) );
  AO22X1_LVT U7807 ( .A1(n6765), .A2(n_T_427[748]), .A3(n3860), .A4(
        n_T_427[237]), .Y(n6400) );
  AO22X1_LVT U7808 ( .A1(n_T_427[621]), .A2(n3796), .A3(n3866), .A4(
        n_T_427[365]), .Y(n6399) );
  AO22X1_LVT U7809 ( .A1(n3838), .A2(n_T_427[493]), .A3(n3873), .A4(
        n_T_427[301]), .Y(n6398) );
  NOR4X1_LVT U7810 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .Y(n6402)
         );
  OA22X1_LVT U7811 ( .A1(n3151), .A2(n3803), .A3(n3503), .A4(n3800), .Y(n6404)
         );
  NAND2X0_LVT U7812 ( .A1(n4442), .A2(n3959), .Y(n6403) );
  AND3X1_LVT U7813 ( .A1(n6405), .A2(n6404), .A3(n6403), .Y(n6406) );
  NAND4X0_LVT U7814 ( .A1(n6408), .A2(n6409), .A3(n6407), .A4(n6406), .Y(
        id_rs_1[45]) );
  NAND2X0_LVT U7815 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[45]), .Y(n6413) );
  NAND2X0_LVT U7816 ( .A1(n6899), .A2(n_T_918[45]), .Y(n6412) );
  NAND2X0_LVT U7817 ( .A1(n6900), .A2(n_T_1165[45]), .Y(n6411) );
  NAND2X0_LVT U7818 ( .A1(n3243), .A2(n_T_635[45]), .Y(n6410) );
  NAND4X0_LVT U7819 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .Y(
        n_T_702[45]) );
  AOI22X1_LVT U7820 ( .A1(n6856), .A2(io_fpu_toint_data[46]), .A3(n6855), .A4(
        n_T_918[46]), .Y(n6414) );
  NAND2X0_LVT U7821 ( .A1(n6857), .A2(n6414), .Y(N644) );
  NAND2X0_LVT U7822 ( .A1(csr_io_rw_rdata[46]), .A2(n3845), .Y(n6417) );
  AOI22X1_LVT U7823 ( .A1(n3853), .A2(io_dmem_resp_bits_data[46]), .A3(n3847), 
        .A4(n_T_1165[46]), .Y(n6416) );
  NAND2X0_LVT U7824 ( .A1(div_io_resp_bits_data[46]), .A2(n3858), .Y(n6415) );
  NAND3X0_LVT U7825 ( .A1(n6417), .A2(n6416), .A3(n6415), .Y(
        n_T_427__T_1136_data[46]) );
  AO22X1_LVT U7826 ( .A1(n3925), .A2(n_T_427[1517]), .A3(n_T_427[1389]), .A4(
        n3920), .Y(n6421) );
  AO22X1_LVT U7827 ( .A1(n3935), .A2(n_T_427[1453]), .A3(n_T_427[1325]), .A4(
        n3930), .Y(n6420) );
  AO22X1_LVT U7828 ( .A1(n3945), .A2(n_T_427[1197]), .A3(n_T_427[1261]), .A4(
        n3940), .Y(n6419) );
  AO22X1_LVT U7829 ( .A1(n3955), .A2(n_T_427[1133]), .A3(n_T_427[1005]), .A4(
        n3950), .Y(n6418) );
  NOR4X1_LVT U7830 ( .A1(n6421), .A2(n6420), .A3(n6419), .A4(n6418), .Y(n6436)
         );
  AOI22X1_LVT U7831 ( .A1(n3870), .A2(n_T_427[558]), .A3(n6868), .A4(
        n_T_427[366]), .Y(n6427) );
  AOI22X1_LVT U7832 ( .A1(n3814), .A2(n_T_427[813]), .A3(n_T_427[877]), .A4(
        n3875), .Y(n6426) );
  OA22X1_LVT U7833 ( .A1(n3522), .A2(n6423), .A3(n3176), .A4(n6422), .Y(n6425)
         );
  AOI22X1_LVT U7834 ( .A1(n_T_427[941]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[622]), .Y(n6424) );
  NAND4X0_LVT U7835 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .Y(n6428) );
  AO22X1_LVT U7836 ( .A1(n2864), .A2(n_T_427[430]), .A3(n_T_427[1069]), .A4(
        n3898), .Y(n6432) );
  AO22X1_LVT U7837 ( .A1(n3911), .A2(n_T_427[494]), .A3(n_T_427[749]), .A4(
        n3905), .Y(n6431) );
  AO22X1_LVT U7838 ( .A1(n2879), .A2(n_T_427[46]), .A3(n_T_427[174]), .A4(
        n2862), .Y(n6430) );
  AO22X1_LVT U7839 ( .A1(n3810), .A2(n_T_427[302]), .A3(n_T_427[686]), .A4(
        n2829), .Y(n6429) );
  NOR4X1_LVT U7840 ( .A1(n6432), .A2(n6431), .A3(n6430), .A4(n6429), .Y(n6434)
         );
  NAND2X0_LVT U7841 ( .A1(n3957), .A2(n4445), .Y(n6433) );
  NAND4X0_LVT U7842 ( .A1(n6436), .A2(n6435), .A3(n6434), .A4(n6433), .Y(
        id_rs_1[46]) );
  NAND2X0_LVT U7843 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[46]), .Y(n6440) );
  NAND2X0_LVT U7844 ( .A1(n6899), .A2(n_T_918[46]), .Y(n6439) );
  NAND2X0_LVT U7845 ( .A1(n6900), .A2(n_T_1165[46]), .Y(n6438) );
  NAND2X0_LVT U7846 ( .A1(n6901), .A2(n_T_635[46]), .Y(n6437) );
  NAND4X0_LVT U7847 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .Y(
        n_T_702[46]) );
  AOI22X1_LVT U7848 ( .A1(n6856), .A2(io_fpu_toint_data[47]), .A3(n6855), .A4(
        n_T_918[47]), .Y(n6441) );
  NAND2X0_LVT U7849 ( .A1(n6857), .A2(n6441), .Y(N645) );
  NAND2X0_LVT U7850 ( .A1(csr_io_rw_rdata[47]), .A2(n3845), .Y(n6444) );
  AOI22X1_LVT U7851 ( .A1(n3853), .A2(io_dmem_resp_bits_data[47]), .A3(n3847), 
        .A4(n_T_1165[47]), .Y(n6443) );
  NAND2X0_LVT U7852 ( .A1(div_io_resp_bits_data[47]), .A2(n3858), .Y(n6442) );
  NAND3X0_LVT U7853 ( .A1(n6444), .A2(n6443), .A3(n6442), .Y(
        n_T_427__T_1136_data[47]) );
  AO22X1_LVT U7854 ( .A1(n3817), .A2(n_T_427[367]), .A3(n_T_427[495]), .A4(
        n3912), .Y(n6446) );
  AO22X1_LVT U7855 ( .A1(n3916), .A2(n_T_427[623]), .A3(n_T_427[878]), .A4(
        n3822), .Y(n6445) );
  NOR2X0_LVT U7856 ( .A1(n6446), .A2(n6445), .Y(n6456) );
  AO22X1_LVT U7857 ( .A1(n_T_427[942]), .A2(n6794), .A3(n3868), .A4(
        n_T_427[559]), .Y(n6450) );
  AO22X1_LVT U7858 ( .A1(n_T_427[687]), .A2(n3861), .A3(n6866), .A4(
        n_T_427[111]), .Y(n6449) );
  AO22X1_LVT U7859 ( .A1(n_T_427[814]), .A2(n3813), .A3(n3873), .A4(
        n_T_427[303]), .Y(n6448) );
  AO22X1_LVT U7860 ( .A1(n3815), .A2(n_T_427[175]), .A3(n3839), .A4(
        n_T_427[47]), .Y(n6447) );
  NOR4X1_LVT U7861 ( .A1(n6450), .A2(n6449), .A3(n6448), .A4(n6447), .Y(n6451)
         );
  OA22X1_LVT U7862 ( .A1(n3556), .A2(n3882), .A3(n3877), .A4(n6451), .Y(n6454)
         );
  NAND2X0_LVT U7863 ( .A1(n3957), .A2(n4448), .Y(n6453) );
  OA22X1_LVT U7864 ( .A1(n3152), .A2(n3803), .A3(n3504), .A4(n3800), .Y(n6452)
         );
  AND3X1_LVT U7865 ( .A1(n6454), .A2(n6453), .A3(n6452), .Y(n6455) );
  NAND4X0_LVT U7866 ( .A1(n6457), .A2(n6458), .A3(n6456), .A4(n6455), .Y(
        id_rs_1[47]) );
  NAND2X0_LVT U7867 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[47]), .Y(n6462) );
  NAND2X0_LVT U7868 ( .A1(n6899), .A2(n_T_918[47]), .Y(n6461) );
  NAND2X0_LVT U7869 ( .A1(n6900), .A2(n_T_1165[47]), .Y(n6460) );
  NAND2X0_LVT U7870 ( .A1(n3243), .A2(n_T_635[47]), .Y(n6459) );
  NAND4X0_LVT U7871 ( .A1(n6462), .A2(n6461), .A3(n6460), .A4(n6459), .Y(
        n_T_702[47]) );
  NAND2X0_LVT U7872 ( .A1(csr_io_rw_rdata[48]), .A2(n3845), .Y(n6465) );
  AOI22X1_LVT U7873 ( .A1(n3853), .A2(io_dmem_resp_bits_data[48]), .A3(n3847), 
        .A4(n_T_1165[48]), .Y(n6464) );
  NAND2X0_LVT U7874 ( .A1(div_io_resp_bits_data[48]), .A2(n3858), .Y(n6463) );
  NAND3X0_LVT U7875 ( .A1(n6465), .A2(n6464), .A3(n6463), .Y(
        n_T_427__T_1136_data[48]) );
  AO22X1_LVT U7876 ( .A1(n3828), .A2(n_T_427[1836]), .A3(n_T_427[1711]), .A4(
        n3824), .Y(n6469) );
  AO22X1_LVT U7877 ( .A1(n3893), .A2(n_T_427[1583]), .A3(n_T_427[1647]), .A4(
        n3888), .Y(n6468) );
  AO22X1_LVT U7878 ( .A1(n3925), .A2(n_T_427[1519]), .A3(n_T_427[1391]), .A4(
        n3920), .Y(n6467) );
  AO22X1_LVT U7879 ( .A1(n3935), .A2(n_T_427[1455]), .A3(n_T_427[1327]), .A4(
        n3930), .Y(n6466) );
  NOR4X1_LVT U7880 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .Y(n6483)
         );
  AO22X1_LVT U7881 ( .A1(n3911), .A2(n_T_427[496]), .A3(n_T_427[751]), .A4(
        n3903), .Y(n6471) );
  AO22X1_LVT U7882 ( .A1(n3915), .A2(n_T_427[624]), .A3(n_T_427[688]), .A4(
        n2829), .Y(n6470) );
  NOR2X0_LVT U7883 ( .A1(n6471), .A2(n6470), .Y(n6481) );
  AO22X1_LVT U7884 ( .A1(n3813), .A2(n_T_427[815]), .A3(n_T_427[879]), .A4(
        n3874), .Y(n6475) );
  AO22X1_LVT U7885 ( .A1(n_T_427[560]), .A2(n3869), .A3(n3873), .A4(
        n_T_427[304]), .Y(n6474) );
  AO22X1_LVT U7886 ( .A1(n3815), .A2(n_T_427[176]), .A3(n3839), .A4(
        n_T_427[48]), .Y(n6473) );
  AO22X1_LVT U7887 ( .A1(n6866), .A2(n_T_427[112]), .A3(n3867), .A4(
        n_T_427[368]), .Y(n6472) );
  NOR4X1_LVT U7888 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .Y(n6476)
         );
  OA22X1_LVT U7889 ( .A1(n3557), .A2(n3882), .A3(n1993), .A4(n6476), .Y(n6479)
         );
  NAND2X0_LVT U7890 ( .A1(n3957), .A2(n4451), .Y(n6478) );
  OA22X1_LVT U7891 ( .A1(n3153), .A2(n3803), .A3(n3505), .A4(n3800), .Y(n6477)
         );
  AND3X1_LVT U7892 ( .A1(n6479), .A2(n6478), .A3(n6477), .Y(n6480) );
  NAND4X0_LVT U7893 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .Y(
        id_rs_1[48]) );
  NAND2X0_LVT U7894 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[48]), .Y(n6487) );
  NAND2X0_LVT U7895 ( .A1(n6899), .A2(n_T_918[48]), .Y(n6486) );
  NAND2X0_LVT U7896 ( .A1(n6900), .A2(n_T_1165[48]), .Y(n6485) );
  NAND2X0_LVT U7897 ( .A1(n3243), .A2(n_T_635[48]), .Y(n6484) );
  NAND4X0_LVT U7898 ( .A1(n6487), .A2(n6486), .A3(n6485), .A4(n6484), .Y(
        n_T_702[48]) );
  AO22X1_LVT U7899 ( .A1(n6860), .A2(io_dmem_resp_bits_data[49]), .A3(n3848), 
        .A4(n_T_1165[49]), .Y(n6488) );
  AO21X1_LVT U7900 ( .A1(n3856), .A2(div_io_resp_bits_data[49]), .A3(n6488), 
        .Y(n6489) );
  AO21X1_LVT U7901 ( .A1(n3842), .A2(csr_io_rw_rdata[49]), .A3(n6489), .Y(
        n_T_427__T_1136_data[49]) );
  AO22X1_LVT U7902 ( .A1(n3830), .A2(n_T_427[1837]), .A3(n_T_427[1712]), .A4(
        n3824), .Y(n6493) );
  AO22X1_LVT U7903 ( .A1(n3893), .A2(n_T_427[1584]), .A3(n_T_427[1648]), .A4(
        n3887), .Y(n6492) );
  AO22X1_LVT U7904 ( .A1(n3925), .A2(n_T_427[1520]), .A3(n_T_427[1392]), .A4(
        n3919), .Y(n6491) );
  AO22X1_LVT U7905 ( .A1(n3935), .A2(n_T_427[1456]), .A3(n_T_427[1328]), .A4(
        n3930), .Y(n6490) );
  NOR4X1_LVT U7906 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .Y(n6507)
         );
  AO22X1_LVT U7907 ( .A1(n2857), .A2(n_T_427[369]), .A3(n_T_427[561]), .A4(
        n2850), .Y(n6495) );
  AO22X1_LVT U7908 ( .A1(n3822), .A2(n_T_427[880]), .A3(n_T_427[305]), .A4(
        n2828), .Y(n6494) );
  NAND2X0_LVT U7909 ( .A1(n4454), .A2(n3959), .Y(n6503) );
  AO22X1_LVT U7910 ( .A1(n_T_427[689]), .A2(n3861), .A3(n3796), .A4(
        n_T_427[625]), .Y(n6499) );
  AO22X1_LVT U7911 ( .A1(n_T_427[944]), .A2(n6794), .A3(n3812), .A4(
        n_T_427[816]), .Y(n6498) );
  AO22X1_LVT U7912 ( .A1(n6867), .A2(n_T_427[433]), .A3(n3860), .A4(
        n_T_427[241]), .Y(n6497) );
  AO22X1_LVT U7913 ( .A1(n3816), .A2(n_T_427[177]), .A3(n3839), .A4(
        n_T_427[49]), .Y(n6496) );
  NOR4X1_LVT U7914 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .Y(n6500)
         );
  OA22X1_LVT U7915 ( .A1(n3154), .A2(n3803), .A3(n3506), .A4(n3800), .Y(n6501)
         );
  AND3X1_LVT U7916 ( .A1(n6503), .A2(n6502), .A3(n6501), .Y(n6504) );
  NAND4X0_LVT U7917 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .Y(
        id_rs_1[49]) );
  NAND2X0_LVT U7918 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[49]), .Y(n6511) );
  NAND2X0_LVT U7919 ( .A1(n6899), .A2(n_T_918[49]), .Y(n6510) );
  NAND2X0_LVT U7920 ( .A1(n6900), .A2(n_T_1165[49]), .Y(n6509) );
  NAND2X0_LVT U7921 ( .A1(n6901), .A2(n_T_635[49]), .Y(n6508) );
  NAND4X0_LVT U7922 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .Y(
        n_T_702[49]) );
  NAND2X0_LVT U7923 ( .A1(csr_io_rw_rdata[50]), .A2(n3845), .Y(n6514) );
  AOI22X1_LVT U7924 ( .A1(n3853), .A2(io_dmem_resp_bits_data[50]), .A3(n3847), 
        .A4(n_T_1165[50]), .Y(n6513) );
  NAND2X0_LVT U7925 ( .A1(div_io_resp_bits_data[50]), .A2(n3857), .Y(n6512) );
  NAND3X0_LVT U7926 ( .A1(n6514), .A2(n6513), .A3(n6512), .Y(
        n_T_427__T_1136_data[50]) );
  AO22X1_LVT U7927 ( .A1(n3945), .A2(n_T_427[1201]), .A3(n_T_427[1265]), .A4(
        n3940), .Y(n6518) );
  AO22X1_LVT U7928 ( .A1(n3955), .A2(n_T_427[1137]), .A3(n_T_427[1009]), .A4(
        n3950), .Y(n6517) );
  AO22X1_LVT U7929 ( .A1(n3901), .A2(n_T_427[1073]), .A3(n_T_427[242]), .A4(
        n2830), .Y(n6516) );
  AO22X1_LVT U7930 ( .A1(n2864), .A2(n_T_427[434]), .A3(n_T_427[114]), .A4(
        n3831), .Y(n6515) );
  NOR4X1_LVT U7931 ( .A1(n6518), .A2(n6517), .A3(n6516), .A4(n6515), .Y(n6531)
         );
  AO22X1_LVT U7932 ( .A1(n3906), .A2(n_T_427[817]), .A3(n_T_427[753]), .A4(
        n3905), .Y(n6520) );
  AO22X1_LVT U7933 ( .A1(n2856), .A2(n_T_427[370]), .A3(n_T_427[306]), .A4(
        n2828), .Y(n6519) );
  NOR2X0_LVT U7934 ( .A1(n6520), .A2(n6519), .Y(n6530) );
  NAND2X0_LVT U7935 ( .A1(n3958), .A2(n4457), .Y(n6528) );
  AO22X1_LVT U7936 ( .A1(n_T_427[690]), .A2(n3861), .A3(n3868), .A4(
        n_T_427[562]), .Y(n6524) );
  AO22X1_LVT U7937 ( .A1(n_T_427[945]), .A2(n6794), .A3(n3875), .A4(
        n_T_427[881]), .Y(n6523) );
  AO22X1_LVT U7938 ( .A1(n3797), .A2(n_T_427[626]), .A3(n_T_427[498]), .A4(
        n3836), .Y(n6522) );
  AO22X1_LVT U7939 ( .A1(n3816), .A2(n_T_427[178]), .A3(n3840), .A4(
        n_T_427[50]), .Y(n6521) );
  NOR4X1_LVT U7940 ( .A1(n6524), .A2(n6523), .A3(n6522), .A4(n6521), .Y(n6525)
         );
  OA22X1_LVT U7941 ( .A1(n3155), .A2(n2027), .A3(n3507), .A4(n3800), .Y(n6526)
         );
  AND3X1_LVT U7942 ( .A1(n6528), .A2(n6527), .A3(n6526), .Y(n6529) );
  NAND4X0_LVT U7943 ( .A1(n6531), .A2(n6532), .A3(n6530), .A4(n6529), .Y(
        id_rs_1[50]) );
  NAND2X0_LVT U7944 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[50]), .Y(n6536) );
  NAND2X0_LVT U7945 ( .A1(n6899), .A2(n_T_918[50]), .Y(n6535) );
  NAND2X0_LVT U7946 ( .A1(n6900), .A2(n_T_1165[50]), .Y(n6534) );
  NAND2X0_LVT U7947 ( .A1(n3243), .A2(n_T_635[50]), .Y(n6533) );
  NAND4X0_LVT U7948 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .Y(
        n_T_702[50]) );
  AO22X1_LVT U7949 ( .A1(n6860), .A2(io_dmem_resp_bits_data[51]), .A3(n3848), 
        .A4(n_T_1165[51]), .Y(n6537) );
  AO21X1_LVT U7950 ( .A1(n3857), .A2(div_io_resp_bits_data[51]), .A3(n6537), 
        .Y(n6538) );
  AO21X1_LVT U7951 ( .A1(n3841), .A2(csr_io_rw_rdata[51]), .A3(n6538), .Y(
        n_T_427__T_1136_data[51]) );
  AO22X1_LVT U7952 ( .A1(n3828), .A2(n_T_427[1839]), .A3(n_T_427[1714]), .A4(
        n3824), .Y(n6542) );
  AO22X1_LVT U7953 ( .A1(n3893), .A2(n_T_427[1586]), .A3(n_T_427[1650]), .A4(
        n3888), .Y(n6541) );
  AO22X1_LVT U7954 ( .A1(n3925), .A2(n_T_427[1522]), .A3(n_T_427[1394]), .A4(
        n3920), .Y(n6540) );
  AO22X1_LVT U7955 ( .A1(n3935), .A2(n_T_427[1458]), .A3(n_T_427[1330]), .A4(
        n3930), .Y(n6539) );
  NOR4X1_LVT U7956 ( .A1(n6542), .A2(n6541), .A3(n6540), .A4(n6539), .Y(n6556)
         );
  AO22X1_LVT U7957 ( .A1(n2851), .A2(n_T_427[563]), .A3(n_T_427[51]), .A4(
        n2879), .Y(n6544) );
  AO22X1_LVT U7958 ( .A1(n3822), .A2(n_T_427[882]), .A3(n_T_427[691]), .A4(
        n3821), .Y(n6543) );
  NOR2X0_LVT U7959 ( .A1(n6544), .A2(n6543), .Y(n6554) );
  AO22X1_LVT U7960 ( .A1(n3815), .A2(n_T_427[179]), .A3(n_T_427[818]), .A4(
        n3812), .Y(n6548) );
  AO22X1_LVT U7961 ( .A1(n6867), .A2(n_T_427[435]), .A3(n6866), .A4(
        n_T_427[115]), .Y(n6547) );
  AO22X1_LVT U7962 ( .A1(n_T_427[627]), .A2(n3797), .A3(n3867), .A4(
        n_T_427[371]), .Y(n6546) );
  AO22X1_LVT U7963 ( .A1(n3838), .A2(n_T_427[499]), .A3(n3873), .A4(
        n_T_427[307]), .Y(n6545) );
  NOR4X1_LVT U7964 ( .A1(n6548), .A2(n6547), .A3(n6546), .A4(n6545), .Y(n6549)
         );
  OA22X1_LVT U7965 ( .A1(n3156), .A2(n3080), .A3(n3508), .A4(n3800), .Y(n6551)
         );
  NAND2X0_LVT U7966 ( .A1(n4460), .A2(n6898), .Y(n6550) );
  AND3X1_LVT U7967 ( .A1(n6552), .A2(n6551), .A3(n6550), .Y(n6553) );
  NAND4X0_LVT U7968 ( .A1(n6556), .A2(n6555), .A3(n6554), .A4(n6553), .Y(
        id_rs_1[51]) );
  NAND2X0_LVT U7969 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[51]), .Y(n6560) );
  NAND2X0_LVT U7970 ( .A1(n6899), .A2(n_T_918[51]), .Y(n6559) );
  NAND2X0_LVT U7971 ( .A1(n6900), .A2(n_T_1165[51]), .Y(n6558) );
  NAND2X0_LVT U7972 ( .A1(n6901), .A2(n_T_635[51]), .Y(n6557) );
  NAND4X0_LVT U7973 ( .A1(n6560), .A2(n6559), .A3(n6558), .A4(n6557), .Y(
        n_T_702[51]) );
  AO22X1_LVT U7974 ( .A1(n6860), .A2(io_dmem_resp_bits_data[52]), .A3(n3848), 
        .A4(n_T_1165[52]), .Y(n6561) );
  AO21X1_LVT U7975 ( .A1(n3856), .A2(div_io_resp_bits_data[52]), .A3(n6561), 
        .Y(n6562) );
  AO21X1_LVT U7976 ( .A1(n3841), .A2(csr_io_rw_rdata[52]), .A3(n6562), .Y(
        n_T_427__T_1136_data[52]) );
  AO22X1_LVT U7977 ( .A1(n3829), .A2(n_T_427[1840]), .A3(n_T_427[1715]), .A4(
        n3824), .Y(n6566) );
  AO22X1_LVT U7978 ( .A1(n3893), .A2(n_T_427[1587]), .A3(n_T_427[1651]), .A4(
        n3888), .Y(n6565) );
  AO22X1_LVT U7979 ( .A1(n3925), .A2(n_T_427[1523]), .A3(n_T_427[1395]), .A4(
        n3920), .Y(n6564) );
  AO22X1_LVT U7980 ( .A1(n3935), .A2(n_T_427[1459]), .A3(n_T_427[1331]), .A4(
        n3930), .Y(n6563) );
  NOR4X1_LVT U7981 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .Y(n6584)
         );
  AO22X1_LVT U7982 ( .A1(n3945), .A2(n_T_427[1203]), .A3(n_T_427[1267]), .A4(
        n3940), .Y(n6570) );
  AO22X1_LVT U7983 ( .A1(n3955), .A2(n_T_427[1139]), .A3(n_T_427[1011]), .A4(
        n3950), .Y(n6569) );
  AO22X1_LVT U7984 ( .A1(n3902), .A2(n_T_427[1075]), .A3(n_T_427[244]), .A4(
        n3806), .Y(n6568) );
  AO22X1_LVT U7985 ( .A1(n2871), .A2(n_T_427[116]), .A3(n_T_427[947]), .A4(
        n3895), .Y(n6567) );
  NOR4X1_LVT U7986 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .Y(n6583)
         );
  AO22X1_LVT U7987 ( .A1(n2860), .A2(n_T_427[819]), .A3(n_T_427[755]), .A4(
        n3904), .Y(n6572) );
  AO22X1_LVT U7988 ( .A1(n2879), .A2(n_T_427[52]), .A3(n_T_427[692]), .A4(
        n3820), .Y(n6571) );
  NOR2X0_LVT U7989 ( .A1(n6572), .A2(n6571), .Y(n6582) );
  AO22X1_LVT U7990 ( .A1(n3816), .A2(n_T_427[180]), .A3(n_T_427[883]), .A4(
        n3874), .Y(n6576) );
  AO22X1_LVT U7991 ( .A1(n3870), .A2(n_T_427[564]), .A3(n_T_427[628]), .A4(
        n3795), .Y(n6575) );
  AO22X1_LVT U7992 ( .A1(n6867), .A2(n_T_427[436]), .A3(n3867), .A4(
        n_T_427[372]), .Y(n6574) );
  AO22X1_LVT U7993 ( .A1(n3838), .A2(n_T_427[500]), .A3(n3873), .A4(
        n_T_427[308]), .Y(n6573) );
  NOR4X1_LVT U7994 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .Y(n6577)
         );
  OA22X1_LVT U7995 ( .A1(n3157), .A2(n1994), .A3(n3509), .A4(n3800), .Y(n6579)
         );
  NAND2X0_LVT U7996 ( .A1(n4463), .A2(n6898), .Y(n6578) );
  AND3X1_LVT U7997 ( .A1(n6580), .A2(n6579), .A3(n6578), .Y(n6581) );
  NAND4X0_LVT U7998 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .Y(
        id_rs_1[52]) );
  NAND2X0_LVT U7999 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[52]), .Y(n6588) );
  NAND2X0_LVT U8000 ( .A1(n6899), .A2(n_T_918[52]), .Y(n6587) );
  NAND2X0_LVT U8001 ( .A1(n6900), .A2(n_T_1165[52]), .Y(n6586) );
  NAND2X0_LVT U8002 ( .A1(n6901), .A2(n_T_635[52]), .Y(n6585) );
  NAND4X0_LVT U8003 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .Y(
        n_T_702[52]) );
  NAND2X0_LVT U8004 ( .A1(csr_io_rw_rdata[53]), .A2(n3845), .Y(n6591) );
  AOI22X1_LVT U8005 ( .A1(n3853), .A2(io_dmem_resp_bits_data[53]), .A3(n3847), 
        .A4(n_T_1165[53]), .Y(n6590) );
  NAND2X0_LVT U8006 ( .A1(div_io_resp_bits_data[53]), .A2(n3857), .Y(n6589) );
  NAND3X0_LVT U8007 ( .A1(n6591), .A2(n6590), .A3(n6589), .Y(
        n_T_427__T_1136_data[53]) );
  AO22X1_LVT U8008 ( .A1(n3946), .A2(n_T_427[1204]), .A3(n_T_427[1268]), .A4(
        n3940), .Y(n6595) );
  AO22X1_LVT U8009 ( .A1(n3956), .A2(n_T_427[1140]), .A3(n_T_427[1012]), .A4(
        n3950), .Y(n6594) );
  AO22X1_LVT U8010 ( .A1(n3902), .A2(n_T_427[1076]), .A3(n_T_427[245]), .A4(
        n3808), .Y(n6593) );
  AO22X1_LVT U8011 ( .A1(n2832), .A2(n_T_427[948]), .A3(n_T_427[756]), .A4(
        n2827), .Y(n6592) );
  NOR4X1_LVT U8012 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .Y(n6608)
         );
  AO22X1_LVT U8013 ( .A1(n3906), .A2(n_T_427[820]), .A3(n_T_427[373]), .A4(
        n1918), .Y(n6597) );
  AO22X1_LVT U8014 ( .A1(n2850), .A2(n_T_427[565]), .A3(n_T_427[693]), .A4(
        n3820), .Y(n6596) );
  NOR2X0_LVT U8015 ( .A1(n6597), .A2(n6596), .Y(n6607) );
  AO22X1_LVT U8016 ( .A1(n3797), .A2(n_T_427[629]), .A3(n_T_427[501]), .A4(
        n3836), .Y(n6601) );
  AO22X1_LVT U8017 ( .A1(n6867), .A2(n_T_427[437]), .A3(n3864), .A4(
        n_T_427[117]), .Y(n6600) );
  AO22X1_LVT U8018 ( .A1(n_T_427[884]), .A2(n6871), .A3(n3873), .A4(
        n_T_427[309]), .Y(n6599) );
  AO22X1_LVT U8019 ( .A1(n3816), .A2(n_T_427[181]), .A3(n3840), .A4(
        n_T_427[53]), .Y(n6598) );
  NOR4X1_LVT U8020 ( .A1(n6601), .A2(n6600), .A3(n6599), .A4(n6598), .Y(n6602)
         );
  OA22X1_LVT U8021 ( .A1(n3561), .A2(n3882), .A3(n1993), .A4(n6602), .Y(n6605)
         );
  NAND2X0_LVT U8022 ( .A1(n3958), .A2(n4466), .Y(n6604) );
  OA22X1_LVT U8023 ( .A1(n3158), .A2(n2027), .A3(n3510), .A4(n3800), .Y(n6603)
         );
  AND3X1_LVT U8024 ( .A1(n6605), .A2(n6604), .A3(n6603), .Y(n6606) );
  NAND4X0_LVT U8025 ( .A1(n6608), .A2(n6609), .A3(n6607), .A4(n6606), .Y(
        id_rs_1[53]) );
  NAND2X0_LVT U8026 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[53]), .Y(n6613) );
  NAND2X0_LVT U8027 ( .A1(n6899), .A2(n_T_918[53]), .Y(n6612) );
  NAND2X0_LVT U8028 ( .A1(n6900), .A2(n_T_1165[53]), .Y(n6611) );
  NAND2X0_LVT U8029 ( .A1(n6901), .A2(n_T_635[53]), .Y(n6610) );
  NAND4X0_LVT U8030 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .Y(
        n_T_702[53]) );
  AO22X1_LVT U8031 ( .A1(n6860), .A2(io_dmem_resp_bits_data[54]), .A3(n3848), 
        .A4(n_T_1165[54]), .Y(n6614) );
  AO21X1_LVT U8032 ( .A1(n3856), .A2(div_io_resp_bits_data[54]), .A3(n6614), 
        .Y(n6615) );
  AO21X1_LVT U8033 ( .A1(n3841), .A2(csr_io_rw_rdata[54]), .A3(n6615), .Y(
        n_T_427__T_1136_data[54]) );
  AO22X1_LVT U8034 ( .A1(n2856), .A2(n_T_427[374]), .A3(n_T_427[182]), .A4(
        n3908), .Y(n6617) );
  AO22X1_LVT U8035 ( .A1(n3809), .A2(n_T_427[310]), .A3(n_T_427[694]), .A4(
        n2829), .Y(n6616) );
  NOR2X0_LVT U8036 ( .A1(n6617), .A2(n6616), .Y(n6627) );
  AO22X1_LVT U8037 ( .A1(n3870), .A2(n_T_427[566]), .A3(n3860), .A4(
        n_T_427[246]), .Y(n6621) );
  AO22X1_LVT U8038 ( .A1(n_T_427[757]), .A2(n3804), .A3(n6866), .A4(
        n_T_427[118]), .Y(n6620) );
  AO22X1_LVT U8039 ( .A1(n3797), .A2(n_T_427[630]), .A3(n_T_427[502]), .A4(
        n3836), .Y(n6619) );
  AO22X1_LVT U8040 ( .A1(n_T_427[885]), .A2(n6871), .A3(n3840), .A4(
        n_T_427[54]), .Y(n6618) );
  NOR4X1_LVT U8041 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .Y(n6622)
         );
  OA22X1_LVT U8042 ( .A1(n3159), .A2(n3080), .A3(n3511), .A4(n3800), .Y(n6624)
         );
  NAND2X0_LVT U8043 ( .A1(n4469), .A2(n6898), .Y(n6623) );
  AND3X1_LVT U8044 ( .A1(n6625), .A2(n6624), .A3(n6623), .Y(n6626) );
  NAND4X0_LVT U8045 ( .A1(n6628), .A2(n6629), .A3(n6627), .A4(n6626), .Y(
        id_rs_1[54]) );
  NAND2X0_LVT U8046 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[54]), .Y(n6633) );
  NAND2X0_LVT U8047 ( .A1(n6899), .A2(n_T_918[54]), .Y(n6632) );
  NAND2X0_LVT U8048 ( .A1(n6900), .A2(n_T_1165[54]), .Y(n6631) );
  NAND2X0_LVT U8049 ( .A1(n3243), .A2(n_T_635[54]), .Y(n6630) );
  NAND4X0_LVT U8050 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .Y(
        n_T_702[54]) );
  NAND2X0_LVT U8051 ( .A1(csr_io_rw_rdata[55]), .A2(n3845), .Y(n6636) );
  AOI22X1_LVT U8052 ( .A1(n3853), .A2(io_dmem_resp_bits_data[55]), .A3(n3847), 
        .A4(n_T_1165[55]), .Y(n6635) );
  NAND2X0_LVT U8053 ( .A1(div_io_resp_bits_data[55]), .A2(n3857), .Y(n6634) );
  NAND3X0_LVT U8054 ( .A1(n6636), .A2(n6635), .A3(n6634), .Y(
        n_T_427__T_1136_data[55]) );
  AO22X1_LVT U8055 ( .A1(n_T_427[695]), .A2(n3862), .A3(n3860), .A4(
        n_T_427[247]), .Y(n6640) );
  AO22X1_LVT U8056 ( .A1(n3816), .A2(n_T_427[183]), .A3(n_T_427[886]), .A4(
        n3874), .Y(n6639) );
  AO22X1_LVT U8057 ( .A1(n6867), .A2(n_T_427[439]), .A3(n6866), .A4(
        n_T_427[119]), .Y(n6638) );
  AO22X1_LVT U8058 ( .A1(n3838), .A2(n_T_427[503]), .A3(n3867), .A4(
        n_T_427[375]), .Y(n6637) );
  NOR4X1_LVT U8059 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .Y(n6641)
         );
  OA22X1_LVT U8060 ( .A1(n3563), .A2(n3882), .A3(n3877), .A4(n6641), .Y(n6645)
         );
  OA22X1_LVT U8061 ( .A1(n3160), .A2(n3080), .A3(n3512), .A4(n3800), .Y(n6644)
         );
  AOI22X1_LVT U8062 ( .A1(n3894), .A2(n_T_427[1590]), .A3(n_T_427[1654]), .A4(
        n3889), .Y(n6643) );
  OA22X1_LVT U8063 ( .A1(n3161), .A2(n3081), .A3(n3513), .A4(n3082), .Y(n6642)
         );
  AND4X1_LVT U8064 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .Y(n6657)
         );
  AO22X1_LVT U8065 ( .A1(n3902), .A2(n_T_427[1078]), .A3(n_T_427[950]), .A4(
        n2832), .Y(n6649) );
  AO22X1_LVT U8066 ( .A1(n2861), .A2(n_T_427[822]), .A3(n_T_427[758]), .A4(
        n2827), .Y(n6648) );
  AO22X1_LVT U8067 ( .A1(n2869), .A2(n_T_427[631]), .A3(n_T_427[55]), .A4(
        n2826), .Y(n6647) );
  AO22X1_LVT U8068 ( .A1(n2850), .A2(n_T_427[567]), .A3(n_T_427[311]), .A4(
        n6774), .Y(n6646) );
  NOR4X1_LVT U8069 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .Y(n6656)
         );
  AO22X1_LVT U8070 ( .A1(n3926), .A2(n_T_427[1526]), .A3(n_T_427[1398]), .A4(
        n3919), .Y(n6653) );
  AO22X1_LVT U8071 ( .A1(n3936), .A2(n_T_427[1462]), .A3(n_T_427[1334]), .A4(
        n3930), .Y(n6652) );
  AO22X1_LVT U8072 ( .A1(n3946), .A2(n_T_427[1206]), .A3(n_T_427[1270]), .A4(
        n3939), .Y(n6651) );
  AO22X1_LVT U8073 ( .A1(n3956), .A2(n_T_427[1142]), .A3(n_T_427[1014]), .A4(
        n3949), .Y(n6650) );
  NOR4X1_LVT U8074 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .Y(n6655)
         );
  NAND2X0_LVT U8075 ( .A1(n3957), .A2(n4472), .Y(n6654) );
  NAND4X0_LVT U8076 ( .A1(n6656), .A2(n6657), .A3(n6655), .A4(n6654), .Y(
        id_rs_1[55]) );
  NAND2X0_LVT U8077 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[55]), .Y(n6661) );
  NAND2X0_LVT U8078 ( .A1(n6899), .A2(n_T_918[55]), .Y(n6660) );
  NAND2X0_LVT U8079 ( .A1(n6900), .A2(n_T_1165[55]), .Y(n6659) );
  NAND2X0_LVT U8080 ( .A1(n6901), .A2(n_T_635[55]), .Y(n6658) );
  NAND4X0_LVT U8081 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .Y(
        n_T_702[55]) );
  AO22X1_LVT U8082 ( .A1(n6860), .A2(io_dmem_resp_bits_data[56]), .A3(n3848), 
        .A4(n_T_1165[56]), .Y(n6662) );
  AO21X1_LVT U8083 ( .A1(n3856), .A2(div_io_resp_bits_data[56]), .A3(n6662), 
        .Y(n6663) );
  AO21X1_LVT U8084 ( .A1(n3841), .A2(csr_io_rw_rdata[56]), .A3(n6663), .Y(
        n_T_427__T_1136_data[56]) );
  AO22X1_LVT U8085 ( .A1(n3830), .A2(n_T_427[1843]), .A3(n_T_427[1719]), .A4(
        n3824), .Y(n6667) );
  AO22X1_LVT U8086 ( .A1(n3894), .A2(n_T_427[1591]), .A3(n_T_427[1655]), .A4(
        n3887), .Y(n6666) );
  AO22X1_LVT U8087 ( .A1(n3926), .A2(n_T_427[1527]), .A3(n_T_427[1399]), .A4(
        n3920), .Y(n6665) );
  AO22X1_LVT U8088 ( .A1(n3936), .A2(n_T_427[1463]), .A3(n_T_427[1335]), .A4(
        n3929), .Y(n6664) );
  NOR4X1_LVT U8089 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .Y(n6681)
         );
  AO22X1_LVT U8090 ( .A1(n1919), .A2(n_T_427[376]), .A3(n_T_427[632]), .A4(
        n2870), .Y(n6669) );
  AO22X1_LVT U8091 ( .A1(n3822), .A2(n_T_427[887]), .A3(n_T_427[696]), .A4(
        n2829), .Y(n6668) );
  NOR2X0_LVT U8092 ( .A1(n6669), .A2(n6668), .Y(n6679) );
  AO22X1_LVT U8093 ( .A1(n3870), .A2(n_T_427[568]), .A3(n3860), .A4(
        n_T_427[248]), .Y(n6673) );
  AO22X1_LVT U8094 ( .A1(n_T_427[759]), .A2(n3804), .A3(n6866), .A4(
        n_T_427[120]), .Y(n6672) );
  AO22X1_LVT U8095 ( .A1(n3838), .A2(n_T_427[504]), .A3(n3873), .A4(
        n_T_427[312]), .Y(n6671) );
  AO22X1_LVT U8096 ( .A1(n_T_427[823]), .A2(n3813), .A3(n3840), .A4(
        n_T_427[56]), .Y(n6670) );
  NOR4X1_LVT U8097 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .Y(n6674)
         );
  NAND2X0_LVT U8098 ( .A1(n4475), .A2(n6898), .Y(n6675) );
  AND3X1_LVT U8099 ( .A1(n6677), .A2(n6676), .A3(n6675), .Y(n6678) );
  NAND4X0_LVT U8100 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .Y(
        id_rs_1[56]) );
  NAND2X0_LVT U8101 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[56]), .Y(n6685) );
  NAND2X0_LVT U8102 ( .A1(n6899), .A2(n_T_918[56]), .Y(n6684) );
  NAND2X0_LVT U8103 ( .A1(n6900), .A2(n_T_1165[56]), .Y(n6683) );
  NAND2X0_LVT U8104 ( .A1(n6901), .A2(n_T_635[56]), .Y(n6682) );
  NAND4X0_LVT U8105 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .Y(
        n_T_702[56]) );
  NAND2X0_LVT U8106 ( .A1(csr_io_rw_rdata[57]), .A2(n3845), .Y(n6688) );
  AOI22X1_LVT U8107 ( .A1(n3853), .A2(io_dmem_resp_bits_data[57]), .A3(n3847), 
        .A4(n_T_1165[57]), .Y(n6687) );
  NAND2X0_LVT U8108 ( .A1(div_io_resp_bits_data[57]), .A2(n3857), .Y(n6686) );
  NAND3X0_LVT U8109 ( .A1(n6688), .A2(n6687), .A3(n6686), .Y(
        n_T_427__T_1136_data[57]) );
  AO22X1_LVT U8110 ( .A1(n3907), .A2(n_T_427[824]), .A3(n_T_427[185]), .A4(
        n3908), .Y(n6690) );
  AO22X1_LVT U8111 ( .A1(n2870), .A2(n_T_427[633]), .A3(n_T_427[888]), .A4(
        n3822), .Y(n6689) );
  NOR2X0_LVT U8112 ( .A1(n6690), .A2(n6689), .Y(n6700) );
  AO22X1_LVT U8113 ( .A1(n_T_427[697]), .A2(n3861), .A3(n3865), .A4(
        n_T_427[441]), .Y(n6694) );
  AO22X1_LVT U8114 ( .A1(n_T_427[952]), .A2(n6794), .A3(n3837), .A4(
        n_T_427[505]), .Y(n6693) );
  AO22X1_LVT U8115 ( .A1(n_T_427[569]), .A2(n3869), .A3(n3867), .A4(
        n_T_427[377]), .Y(n6692) );
  AO22X1_LVT U8116 ( .A1(n3871), .A2(n_T_427[313]), .A3(n3840), .A4(
        n_T_427[57]), .Y(n6691) );
  NOR4X1_LVT U8117 ( .A1(n6694), .A2(n6693), .A3(n6692), .A4(n6691), .Y(n6695)
         );
  NAND2X0_LVT U8118 ( .A1(n3958), .A2(n4478), .Y(n6697) );
  OA22X1_LVT U8119 ( .A1(n3163), .A2(n3080), .A3(n3515), .A4(n3800), .Y(n6696)
         );
  AND3X1_LVT U8120 ( .A1(n6698), .A2(n6697), .A3(n6696), .Y(n6699) );
  NAND4X0_LVT U8121 ( .A1(n6701), .A2(n6702), .A3(n6700), .A4(n6699), .Y(
        id_rs_1[57]) );
  NAND2X0_LVT U8122 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[57]), .Y(n6706) );
  NAND2X0_LVT U8123 ( .A1(n6899), .A2(n_T_918[57]), .Y(n6705) );
  NAND2X0_LVT U8124 ( .A1(n6900), .A2(n_T_1165[57]), .Y(n6704) );
  NAND2X0_LVT U8125 ( .A1(n3243), .A2(n_T_635[57]), .Y(n6703) );
  NAND4X0_LVT U8126 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .Y(
        n_T_702[57]) );
  AO22X1_LVT U8127 ( .A1(n6860), .A2(io_dmem_resp_bits_data[58]), .A3(n3849), 
        .A4(n_T_1165[58]), .Y(n6707) );
  AO21X1_LVT U8128 ( .A1(n3856), .A2(div_io_resp_bits_data[58]), .A3(n6707), 
        .Y(n6708) );
  AO21X1_LVT U8129 ( .A1(n3841), .A2(csr_io_rw_rdata[58]), .A3(n6708), .Y(
        n_T_427__T_1136_data[58]) );
  AO22X1_LVT U8130 ( .A1(n3828), .A2(n_T_427[1845]), .A3(n_T_427[1721]), .A4(
        n3824), .Y(n6712) );
  AO22X1_LVT U8131 ( .A1(n3894), .A2(n_T_427[1593]), .A3(n_T_427[1657]), .A4(
        n3888), .Y(n6711) );
  AO22X1_LVT U8132 ( .A1(n3926), .A2(n_T_427[1529]), .A3(n_T_427[1401]), .A4(
        n3921), .Y(n6710) );
  AO22X1_LVT U8133 ( .A1(n3936), .A2(n_T_427[1465]), .A3(n_T_427[1337]), .A4(
        n3931), .Y(n6709) );
  NOR4X1_LVT U8134 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .Y(n6727)
         );
  AO22X1_LVT U8135 ( .A1(n3912), .A2(n_T_427[506]), .A3(n_T_427[889]), .A4(
        n2833), .Y(n6714) );
  AO22X1_LVT U8136 ( .A1(n3810), .A2(n_T_427[314]), .A3(n_T_427[698]), .A4(
        n3820), .Y(n6713) );
  NOR2X0_LVT U8137 ( .A1(n6714), .A2(n6713), .Y(n6725) );
  AO22X1_LVT U8138 ( .A1(n_T_427[953]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[634]), .Y(n6719) );
  AO22X1_LVT U8139 ( .A1(n6867), .A2(n_T_427[442]), .A3(n6866), .A4(
        n_T_427[122]), .Y(n6718) );
  AO22X1_LVT U8140 ( .A1(n_T_427[570]), .A2(n3869), .A3(n3867), .A4(
        n_T_427[378]), .Y(n6717) );
  AO22X1_LVT U8141 ( .A1(n3816), .A2(n_T_427[186]), .A3(n3840), .A4(
        n_T_427[58]), .Y(n6716) );
  NOR4X1_LVT U8142 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .Y(n6720)
         );
  OA22X1_LVT U8143 ( .A1(n3164), .A2(n3080), .A3(n3516), .A4(n3800), .Y(n6722)
         );
  NAND2X0_LVT U8144 ( .A1(n4481), .A2(n3958), .Y(n6721) );
  AND3X1_LVT U8145 ( .A1(n6723), .A2(n6722), .A3(n6721), .Y(n6724) );
  NAND4X0_LVT U8146 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .Y(
        id_rs_1[58]) );
  NAND2X0_LVT U8147 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[58]), .Y(n6731) );
  NAND2X0_LVT U8148 ( .A1(n6899), .A2(n_T_918[58]), .Y(n6730) );
  NAND2X0_LVT U8149 ( .A1(n6900), .A2(n_T_1165[58]), .Y(n6729) );
  NAND2X0_LVT U8150 ( .A1(n3243), .A2(n_T_635[58]), .Y(n6728) );
  NAND4X0_LVT U8151 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .Y(
        n_T_702[58]) );
  NAND2X0_LVT U8152 ( .A1(csr_io_rw_rdata[59]), .A2(n3845), .Y(n6734) );
  AOI22X1_LVT U8153 ( .A1(n3853), .A2(io_dmem_resp_bits_data[59]), .A3(n3847), 
        .A4(n_T_1165[59]), .Y(n6733) );
  NAND2X0_LVT U8154 ( .A1(div_io_resp_bits_data[59]), .A2(n3857), .Y(n6732) );
  NAND3X0_LVT U8155 ( .A1(n6734), .A2(n6733), .A3(n6732), .Y(
        n_T_427__T_1136_data[59]) );
  AO22X1_LVT U8156 ( .A1(n3814), .A2(n_T_427[826]), .A3(n_T_427[890]), .A4(
        n3874), .Y(n6738) );
  AO22X1_LVT U8157 ( .A1(n_T_427[699]), .A2(n3861), .A3(n6866), .A4(
        n_T_427[123]), .Y(n6737) );
  AO22X1_LVT U8158 ( .A1(n3838), .A2(n_T_427[507]), .A3(n3867), .A4(
        n_T_427[379]), .Y(n6736) );
  AO22X1_LVT U8159 ( .A1(n3816), .A2(n_T_427[187]), .A3(n3840), .A4(
        n_T_427[59]), .Y(n6735) );
  NOR4X1_LVT U8160 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .Y(n6739)
         );
  OA22X1_LVT U8161 ( .A1(n3165), .A2(n2027), .A3(n3517), .A4(n3800), .Y(n6742)
         );
  OA22X1_LVT U8162 ( .A1(n3166), .A2(n3081), .A3(n3518), .A4(n3082), .Y(n6741)
         );
  AOI22X1_LVT U8163 ( .A1(n3894), .A2(n_T_427[1594]), .A3(n_T_427[1658]), .A4(
        n3889), .Y(n6740) );
  AND4X1_LVT U8164 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .Y(n6755)
         );
  AO22X1_LVT U8165 ( .A1(n3902), .A2(n_T_427[1082]), .A3(n_T_427[251]), .A4(
        n3808), .Y(n6747) );
  AO22X1_LVT U8166 ( .A1(n2864), .A2(n_T_427[443]), .A3(n_T_427[954]), .A4(
        n3897), .Y(n6746) );
  AO22X1_LVT U8167 ( .A1(n3915), .A2(n_T_427[635]), .A3(n_T_427[762]), .A4(
        n2827), .Y(n6745) );
  AO22X1_LVT U8168 ( .A1(n2851), .A2(n_T_427[571]), .A3(n_T_427[315]), .A4(
        n2828), .Y(n6744) );
  NOR4X1_LVT U8169 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .Y(n6754)
         );
  AO22X1_LVT U8170 ( .A1(n3926), .A2(n_T_427[1530]), .A3(n_T_427[1402]), .A4(
        n3920), .Y(n6751) );
  AO22X1_LVT U8171 ( .A1(n3936), .A2(n_T_427[1466]), .A3(n_T_427[1338]), .A4(
        n3931), .Y(n6750) );
  AO22X1_LVT U8172 ( .A1(n3946), .A2(n_T_427[1210]), .A3(n_T_427[1274]), .A4(
        n3940), .Y(n6749) );
  AO22X1_LVT U8173 ( .A1(n3956), .A2(n_T_427[1146]), .A3(n_T_427[1018]), .A4(
        n3950), .Y(n6748) );
  NOR4X1_LVT U8174 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .Y(n6753)
         );
  NAND2X0_LVT U8175 ( .A1(n3957), .A2(n4484), .Y(n6752) );
  NAND4X0_LVT U8176 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .Y(
        id_rs_1[59]) );
  NAND2X0_LVT U8177 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[59]), .Y(n6759) );
  NAND2X0_LVT U8178 ( .A1(n6899), .A2(n_T_918[59]), .Y(n6758) );
  NAND2X0_LVT U8179 ( .A1(n6900), .A2(n_T_1165[59]), .Y(n6757) );
  NAND2X0_LVT U8180 ( .A1(n6901), .A2(n_T_635[59]), .Y(n6756) );
  NAND4X0_LVT U8181 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .Y(
        n_T_702[59]) );
  NAND2X0_LVT U8182 ( .A1(csr_io_rw_rdata[60]), .A2(n3845), .Y(n6762) );
  AOI22X1_LVT U8183 ( .A1(n3853), .A2(io_dmem_resp_bits_data[60]), .A3(n3847), 
        .A4(n_T_1165[60]), .Y(n6761) );
  NAND2X0_LVT U8184 ( .A1(div_io_resp_bits_data[60]), .A2(n3857), .Y(n6760) );
  NAND3X0_LVT U8185 ( .A1(n6762), .A2(n6761), .A3(n6760), .Y(
        n_T_427__T_1136_data[60]) );
  AOI22X1_LVT U8186 ( .A1(n6765), .A2(n_T_427[763]), .A3(n3864), .A4(
        n_T_427[124]), .Y(n6771) );
  AOI22X1_LVT U8187 ( .A1(n3814), .A2(n_T_427[827]), .A3(n6838), .A4(
        n_T_427[60]), .Y(n6770) );
  AOI22X1_LVT U8188 ( .A1(n3838), .A2(n_T_427[508]), .A3(n_T_427[572]), .A4(
        n3868), .Y(n6769) );
  OA22X1_LVT U8189 ( .A1(n6767), .A2(n3525), .A3(n3172), .A4(n6766), .Y(n6768)
         );
  NAND4X0_LVT U8190 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .Y(n6772) );
  AO22X1_LVT U8191 ( .A1(n3902), .A2(n_T_427[1083]), .A3(n_T_427[252]), .A4(
        n3807), .Y(n6778) );
  AO22X1_LVT U8192 ( .A1(n3915), .A2(n_T_427[636]), .A3(n_T_427[891]), .A4(
        n6813), .Y(n6777) );
  AO22X1_LVT U8193 ( .A1(n2831), .A2(n_T_427[955]), .A3(n_T_427[188]), .A4(
        n2862), .Y(n6776) );
  AO22X1_LVT U8194 ( .A1(n3810), .A2(n_T_427[316]), .A3(n_T_427[700]), .A4(
        n3821), .Y(n6775) );
  NOR4X1_LVT U8195 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .Y(n6785)
         );
  AO22X1_LVT U8196 ( .A1(n3926), .A2(n_T_427[1531]), .A3(n_T_427[1403]), .A4(
        n3921), .Y(n6782) );
  AO22X1_LVT U8197 ( .A1(n3936), .A2(n_T_427[1467]), .A3(n_T_427[1339]), .A4(
        n3931), .Y(n6781) );
  AO22X1_LVT U8198 ( .A1(n3946), .A2(n_T_427[1211]), .A3(n_T_427[1275]), .A4(
        n3941), .Y(n6780) );
  AO22X1_LVT U8199 ( .A1(n3956), .A2(n_T_427[1147]), .A3(n_T_427[1019]), .A4(
        n3951), .Y(n6779) );
  NOR4X1_LVT U8200 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .Y(n6784)
         );
  NAND2X0_LVT U8201 ( .A1(n3957), .A2(n4487), .Y(n6783) );
  NAND4X0_LVT U8202 ( .A1(n6785), .A2(n6786), .A3(n6784), .A4(n6783), .Y(
        id_rs_1[60]) );
  NAND2X0_LVT U8203 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[60]), .Y(n6790) );
  NAND2X0_LVT U8204 ( .A1(n6899), .A2(n_T_918[60]), .Y(n6789) );
  NAND2X0_LVT U8205 ( .A1(n6900), .A2(n_T_1165[60]), .Y(n6788) );
  NAND2X0_LVT U8206 ( .A1(n6901), .A2(n_T_635[60]), .Y(n6787) );
  NAND4X0_LVT U8207 ( .A1(n6790), .A2(n6789), .A3(n6788), .A4(n6787), .Y(
        n_T_702[60]) );
  NAND2X0_LVT U8208 ( .A1(csr_io_rw_rdata[61]), .A2(n3842), .Y(n6793) );
  AOI22X1_LVT U8209 ( .A1(n3853), .A2(io_dmem_resp_bits_data[61]), .A3(n3847), 
        .A4(n_T_1165[61]), .Y(n6792) );
  NAND2X0_LVT U8210 ( .A1(div_io_resp_bits_data[61]), .A2(n3857), .Y(n6791) );
  NAND3X0_LVT U8211 ( .A1(n6793), .A2(n6792), .A3(n6791), .Y(
        n_T_427__T_1136_data[61]) );
  AO22X1_LVT U8212 ( .A1(n_T_427[956]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[509]), .Y(n6800) );
  AO22X1_LVT U8213 ( .A1(n_T_427[828]), .A2(n3813), .A3(n3873), .A4(
        n_T_427[317]), .Y(n6799) );
  AO22X1_LVT U8214 ( .A1(n3816), .A2(n_T_427[189]), .A3(n3840), .A4(
        n_T_427[61]), .Y(n6798) );
  AO22X1_LVT U8215 ( .A1(n3860), .A2(n_T_427[253]), .A3(n6866), .A4(
        n_T_427[125]), .Y(n6797) );
  NOR4X1_LVT U8216 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .Y(n6801)
         );
  OA22X1_LVT U8217 ( .A1(n3167), .A2(n1994), .A3(n3485), .A4(n3800), .Y(n6804)
         );
  OA22X1_LVT U8218 ( .A1(n3168), .A2(n3081), .A3(n3486), .A4(n3082), .Y(n6803)
         );
  AOI22X1_LVT U8219 ( .A1(n3894), .A2(n_T_427[1596]), .A3(n_T_427[1660]), .A4(
        n3889), .Y(n6802) );
  AND4X1_LVT U8220 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .Y(n6821)
         );
  AO22X1_LVT U8221 ( .A1(n3926), .A2(n_T_427[1532]), .A3(n_T_427[1404]), .A4(
        n3921), .Y(n6809) );
  AO22X1_LVT U8222 ( .A1(n3936), .A2(n_T_427[1468]), .A3(n_T_427[1340]), .A4(
        n3931), .Y(n6808) );
  AO22X1_LVT U8223 ( .A1(n3946), .A2(n_T_427[1212]), .A3(n_T_427[1276]), .A4(
        n3941), .Y(n6807) );
  AO22X1_LVT U8224 ( .A1(n3956), .A2(n_T_427[1148]), .A3(n_T_427[1020]), .A4(
        n3951), .Y(n6806) );
  NOR4X1_LVT U8225 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .Y(n6820)
         );
  AO22X1_LVT U8226 ( .A1(n3834), .A2(n_T_427[445]), .A3(n_T_427[1084]), .A4(
        n3898), .Y(n6817) );
  AO22X1_LVT U8227 ( .A1(n1918), .A2(n_T_427[381]), .A3(n_T_427[764]), .A4(
        n3903), .Y(n6816) );
  AO22X1_LVT U8228 ( .A1(n3818), .A2(n_T_427[573]), .A3(n_T_427[637]), .A4(
        n2869), .Y(n6815) );
  AO22X1_LVT U8229 ( .A1(n3823), .A2(n_T_427[892]), .A3(n_T_427[701]), .A4(
        n3821), .Y(n6814) );
  NOR4X1_LVT U8230 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(n6814), .Y(n6819)
         );
  NAND2X0_LVT U8231 ( .A1(n3958), .A2(n4490), .Y(n6818) );
  NAND4X0_LVT U8232 ( .A1(n6820), .A2(n6821), .A3(n6819), .A4(n6818), .Y(
        id_rs_1[61]) );
  NAND2X0_LVT U8233 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[61]), .Y(n6825) );
  NAND2X0_LVT U8234 ( .A1(n6899), .A2(n_T_918[61]), .Y(n6824) );
  NAND2X0_LVT U8235 ( .A1(n6900), .A2(n_T_1165[61]), .Y(n6823) );
  NAND2X0_LVT U8236 ( .A1(n3243), .A2(n_T_635[61]), .Y(n6822) );
  NAND4X0_LVT U8237 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .Y(
        n_T_702[61]) );
  NAND2X0_LVT U8238 ( .A1(csr_io_rw_rdata[62]), .A2(n3844), .Y(n6828) );
  AOI22X1_LVT U8239 ( .A1(n3852), .A2(io_dmem_resp_bits_data[62]), .A3(n3847), 
        .A4(n_T_1165[62]), .Y(n6827) );
  NAND2X0_LVT U8240 ( .A1(div_io_resp_bits_data[62]), .A2(n3857), .Y(n6826) );
  NAND3X0_LVT U8241 ( .A1(n6828), .A2(n6827), .A3(n6826), .Y(
        n_T_427__T_1136_data[62]) );
  AO22X1_LVT U8242 ( .A1(n3946), .A2(n_T_427[1213]), .A3(n_T_427[1277]), .A4(
        n3940), .Y(n6834) );
  AO22X1_LVT U8243 ( .A1(n3956), .A2(n_T_427[1149]), .A3(n_T_427[1021]), .A4(
        n3950), .Y(n6833) );
  AO22X1_LVT U8244 ( .A1(n3902), .A2(n_T_427[1085]), .A3(n_T_427[957]), .A4(
        n2832), .Y(n6832) );
  AO22X1_LVT U8245 ( .A1(n2864), .A2(n_T_427[446]), .A3(n_T_427[126]), .A4(
        n2872), .Y(n6831) );
  NOR4X1_LVT U8246 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .Y(n6849)
         );
  AO22X1_LVT U8247 ( .A1(n2860), .A2(n_T_427[829]), .A3(n_T_427[765]), .A4(
        n2827), .Y(n6836) );
  AO22X1_LVT U8248 ( .A1(n2869), .A2(n_T_427[638]), .A3(n_T_427[190]), .A4(
        n2863), .Y(n6835) );
  NOR2X0_LVT U8249 ( .A1(n6836), .A2(n6835), .Y(n6848) );
  AO22X1_LVT U8250 ( .A1(n_T_427[702]), .A2(n3861), .A3(n3860), .A4(
        n_T_427[254]), .Y(n6842) );
  AO22X1_LVT U8251 ( .A1(n_T_427[574]), .A2(n3868), .A3(n6868), .A4(
        n_T_427[382]), .Y(n6841) );
  AO22X1_LVT U8252 ( .A1(n3837), .A2(n_T_427[510]), .A3(n3873), .A4(
        n_T_427[318]), .Y(n6840) );
  AO22X1_LVT U8253 ( .A1(n_T_427[893]), .A2(n6871), .A3(n6838), .A4(
        n_T_427[62]), .Y(n6839) );
  NOR4X1_LVT U8254 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .Y(n6843)
         );
  NAND2X0_LVT U8255 ( .A1(n3957), .A2(n4493), .Y(n6845) );
  OA22X1_LVT U8256 ( .A1(n3169), .A2(n2027), .A3(n3487), .A4(n3800), .Y(n6844)
         );
  AND3X1_LVT U8257 ( .A1(n6846), .A2(n6845), .A3(n6844), .Y(n6847) );
  NAND4X0_LVT U8258 ( .A1(n6849), .A2(n6850), .A3(n6848), .A4(n6847), .Y(
        id_rs_1[62]) );
  NAND2X0_LVT U8259 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[62]), .Y(n6854) );
  NAND2X0_LVT U8260 ( .A1(n6899), .A2(n_T_918[62]), .Y(n6853) );
  NAND2X0_LVT U8261 ( .A1(n6900), .A2(n_T_1165[62]), .Y(n6852) );
  NAND2X0_LVT U8262 ( .A1(n6901), .A2(n_T_635[62]), .Y(n6851) );
  NAND4X0_LVT U8263 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .Y(
        n_T_702[62]) );
  NAND2X0_LVT U8264 ( .A1(csr_io_rw_rdata[63]), .A2(n3844), .Y(n6864) );
  AOI22X1_LVT U8265 ( .A1(n3852), .A2(io_dmem_resp_bits_data[63]), .A3(n3847), 
        .A4(n_T_1165[63]), .Y(n6863) );
  NAND2X0_LVT U8266 ( .A1(div_io_resp_bits_data[63]), .A2(n3858), .Y(n6862) );
  NAND3X0_LVT U8267 ( .A1(n6864), .A2(n6863), .A3(n6862), .Y(
        n_T_427__T_1136_data[63]) );
  AO22X1_LVT U8268 ( .A1(n_T_427[703]), .A2(n3861), .A3(n3859), .A4(
        n_T_427[255]), .Y(n6875) );
  AO22X1_LVT U8269 ( .A1(n6867), .A2(n_T_427[447]), .A3(n3864), .A4(
        n_T_427[127]), .Y(n6874) );
  AO22X1_LVT U8270 ( .A1(n_T_427[575]), .A2(n3869), .A3(n3866), .A4(
        n_T_427[383]), .Y(n6873) );
  AO22X1_LVT U8271 ( .A1(n_T_427[894]), .A2(n3875), .A3(n3871), .A4(
        n_T_427[319]), .Y(n6872) );
  NOR4X1_LVT U8272 ( .A1(n6875), .A2(n6874), .A3(n6873), .A4(n6872), .Y(n6876)
         );
  OA22X1_LVT U8273 ( .A1(n3529), .A2(n3882), .A3(n3878), .A4(n6876), .Y(n6881)
         );
  NAND2X0_LVT U8274 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[63]), .Y(n6905) );
  NAND2X0_LVT U8275 ( .A1(n6899), .A2(n_T_918[63]), .Y(n6904) );
  NAND2X0_LVT U8276 ( .A1(n_T_1165[63]), .A2(n6900), .Y(n6903) );
  NAND2X0_LVT U8277 ( .A1(n6901), .A2(n_T_635[63]), .Y(n6902) );
  NAND4X0_LVT U8278 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .Y(
        n_T_702[63]) );
  NAND2X0_LVT U8279 ( .A1(ibuf_io_inst_0_bits_rvc), .A2(n6912), .Y(n6913) );
  NAND2X0_LVT U8280 ( .A1(n4001), .A2(n_T_427[1728]), .Y(n6918) );
  OA21X1_LVT U8281 ( .A1(n3747), .A2(n3138), .A3(n6918), .Y(n6921) );
  NAND2X0_LVT U8282 ( .A1(n3648), .A2(n_T_427[1600]), .Y(n6920) );
  NAND2X0_LVT U8283 ( .A1(n3657), .A2(n_T_427[1664]), .Y(n6919) );
  NAND2X0_LVT U8284 ( .A1(n3670), .A2(n_T_427[1088]), .Y(n6925) );
  OA21X1_LVT U8285 ( .A1(n3416), .A2(n2897), .A3(n6925), .Y(n6929) );
  NAND2X0_LVT U8286 ( .A1(n3621), .A2(n_T_427[1536]), .Y(n6928) );
  NAND2X0_LVT U8287 ( .A1(n3641), .A2(n_T_427[1216]), .Y(n6927) );
  NAND2X0_LVT U8288 ( .A1(n2966), .A2(n_T_427[1408]), .Y(n6930) );
  OA21X1_LVT U8289 ( .A1(n3987), .A2(n3654), .A3(n6930), .Y(n6934) );
  NAND2X0_LVT U8290 ( .A1(n3606), .A2(n_T_427[1344]), .Y(n6933) );
  NAND2X0_LVT U8291 ( .A1(n3999), .A2(n_T_427[1280]), .Y(n6932) );
  AND2X1_LVT U8292 ( .A1(n6937), .A2(n6936), .Y(n6938) );
  NAND2X0_LVT U8293 ( .A1(n3991), .A2(n_T_427[1883]), .Y(n6942) );
  NAND2X0_LVT U8294 ( .A1(n3712), .A2(n_T_427[960]), .Y(n6970) );
  AND2X1_LVT U8295 ( .A1(n4051), .A2(n_T_427[1]), .Y(n6953) );
  AO22X1_LVT U8296 ( .A1(n4023), .A2(n_T_427[896]), .A3(n4020), .A4(
        n_T_427[641]), .Y(n6952) );
  AND2X1_LVT U8297 ( .A1(n6974), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n8980) );
  AO22X1_LVT U8298 ( .A1(n3977), .A2(n_T_427[513]), .A3(n4027), .A4(
        n_T_427[832]), .Y(n6951) );
  AO22X1_LVT U8299 ( .A1(n4033), .A2(n_T_427[577]), .A3(n3985), .A4(
        n_T_427[193]), .Y(n6950) );
  NOR4X1_LVT U8300 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .Y(n6968)
         );
  AO22X1_LVT U8301 ( .A1(n3968), .A2(n_T_427[385]), .A3(n3964), .A4(
        n_T_427[257]), .Y(n6961) );
  AO22X1_LVT U8302 ( .A1(n2858), .A2(n_T_427[129]), .A3(n4039), .A4(
        n_T_427[321]), .Y(n6960) );
  AND2X1_LVT U8303 ( .A1(n6954), .A2(n2825), .Y(n8981) );
  AO22X1_LVT U8304 ( .A1(n3981), .A2(n_T_427[768]), .A3(n4047), .A4(
        n_T_427[705]), .Y(n6959) );
  AND2X1_LVT U8305 ( .A1(n6957), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n8900) );
  AO22X1_LVT U8306 ( .A1(n3962), .A2(n_T_427[449]), .A3(n4044), .A4(
        n_T_427[65]), .Y(n6958) );
  NOR4X1_LVT U8307 ( .A1(n6961), .A2(n6960), .A3(n6959), .A4(n6958), .Y(n6967)
         );
  AND3X1_LVT U8308 ( .A1(n6971), .A2(n6970), .A3(n6969), .Y(n6978) );
  NAND2X0_LVT U8309 ( .A1(n2611), .A2(n_T_427[1152]), .Y(n6977) );
  NAND2X0_LVT U8310 ( .A1(n4014), .A2(n_T_427[1024]), .Y(n6976) );
  NAND2X0_LVT U8311 ( .A1(n4002), .A2(n_T_427[1727]), .Y(n6979) );
  OA21X1_LVT U8312 ( .A1(n3601), .A2(n3311), .A3(n6979), .Y(n6982) );
  NAND2X0_LVT U8313 ( .A1(n3651), .A2(n_T_427[1599]), .Y(n6981) );
  NAND2X0_LVT U8314 ( .A1(n2922), .A2(n_T_427[1663]), .Y(n6980) );
  NAND2X0_LVT U8315 ( .A1(n3671), .A2(n_T_427[1087]), .Y(n6983) );
  OA21X1_LVT U8316 ( .A1(n3417), .A2(n3653), .A3(n6983), .Y(n6986) );
  NAND2X0_LVT U8317 ( .A1(n3616), .A2(n_T_427[1535]), .Y(n6985) );
  NAND2X0_LVT U8318 ( .A1(n3636), .A2(n_T_427[1215]), .Y(n6984) );
  NAND2X0_LVT U8319 ( .A1(n3630), .A2(n_T_427[1407]), .Y(n6987) );
  OA21X1_LVT U8320 ( .A1(n2969), .A2(n3633), .A3(n6987), .Y(n6990) );
  NAND2X0_LVT U8321 ( .A1(n3607), .A2(n_T_427[1343]), .Y(n6989) );
  NAND2X0_LVT U8322 ( .A1(n3997), .A2(n_T_427[1279]), .Y(n6988) );
  NAND3X0_LVT U8323 ( .A1(n6995), .A2(n9288), .A3(n6994), .Y(n6998) );
  NAND2X0_LVT U8324 ( .A1(n2882), .A2(n_T_427[1882]), .Y(n6996) );
  NAND2X0_LVT U8325 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[0]), .Y(n7011)
         );
  NAND2X0_LVT U8326 ( .A1(n3712), .A2(n_T_427[959]), .Y(n7010) );
  AND2X1_LVT U8327 ( .A1(n4049), .A2(n_T_427[0]), .Y(n7002) );
  AO22X1_LVT U8328 ( .A1(n4026), .A2(n_T_427[895]), .A3(n4018), .A4(
        n_T_427[640]), .Y(n7001) );
  AO22X1_LVT U8329 ( .A1(n3976), .A2(n_T_427[512]), .A3(n4030), .A4(
        n_T_427[831]), .Y(n7000) );
  AO22X1_LVT U8330 ( .A1(n4032), .A2(n_T_427[576]), .A3(n3983), .A4(
        n_T_427[192]), .Y(n6999) );
  NOR4X1_LVT U8331 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .Y(n7008)
         );
  AO22X1_LVT U8332 ( .A1(n3968), .A2(n_T_427[384]), .A3(n3964), .A4(
        n_T_427[256]), .Y(n7006) );
  AO22X1_LVT U8333 ( .A1(n3975), .A2(n_T_427[128]), .A3(n4039), .A4(
        n_T_427[320]), .Y(n7005) );
  AO22X1_LVT U8334 ( .A1(n3979), .A2(n_T_427[767]), .A3(n4045), .A4(
        n_T_427[704]), .Y(n7004) );
  AO22X1_LVT U8335 ( .A1(n3960), .A2(n_T_427[448]), .A3(n2837), .A4(
        n_T_427[64]), .Y(n7003) );
  NOR4X1_LVT U8336 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .Y(n7007)
         );
  AND3X1_LVT U8337 ( .A1(n7011), .A2(n7010), .A3(n7009), .Y(n7014) );
  NAND2X0_LVT U8338 ( .A1(n2611), .A2(n_T_427[1151]), .Y(n7013) );
  NAND2X0_LVT U8339 ( .A1(n4014), .A2(n_T_427[1023]), .Y(n7012) );
  OR2X1_LVT U8340 ( .A1(n2497), .A2(n_T_918[0]), .Y(n7015) );
  AND2X1_LVT U8341 ( .A1(n3101), .A2(n_T_628[1]), .Y(n7017) );
  AO22X1_LVT U8342 ( .A1(n7019), .A2(n7015), .A3(n7017), .A4(
        io_imem_sfence_bits_addr[0]), .Y(n7016) );
  NAND2X0_LVT U8343 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[1]), .Y(n7022)
         );
  NAND3X0_LVT U8344 ( .A1(n7019), .A2(n_T_628[1]), .A3(
        io_fpu_dmem_resp_data[1]), .Y(n7018) );
  OA21X1_LVT U8345 ( .A1(n3101), .A2(n3255), .A3(n7018), .Y(n7021) );
  NAND2X0_LVT U8346 ( .A1(n9066), .A2(n_T_918[1]), .Y(n7020) );
  NAND3X0_LVT U8347 ( .A1(n7022), .A2(n7021), .A3(n7020), .Y(
        io_fpu_fromint_data[1]) );
  NAND2X0_LVT U8348 ( .A1(n3997), .A2(n_T_427[1281]), .Y(n7023) );
  OA21X1_LVT U8349 ( .A1(n3377), .A2(n3684), .A3(n7023), .Y(n7026) );
  NAND2X0_LVT U8350 ( .A1(n3990), .A2(n_T_427[1848]), .Y(n7025) );
  NAND2X0_LVT U8351 ( .A1(n_T_427[1792]), .A2(n3715), .Y(n7024) );
  NAND2X0_LVT U8352 ( .A1(n3619), .A2(n_T_427[1537]), .Y(n7027) );
  OA21X1_LVT U8353 ( .A1(n3418), .A2(n3653), .A3(n7027), .Y(n7030) );
  NAND2X0_LVT U8354 ( .A1(n4004), .A2(n_T_427[1729]), .Y(n7029) );
  NAND2X0_LVT U8355 ( .A1(n3652), .A2(n_T_427[1601]), .Y(n7028) );
  NAND2X0_LVT U8356 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[2]), .Y(n7043)
         );
  NAND2X0_LVT U8357 ( .A1(n3717), .A2(n_T_427[1025]), .Y(n7042) );
  AND2X1_LVT U8358 ( .A1(n4049), .A2(n_T_427[2]), .Y(n7034) );
  AO22X1_LVT U8359 ( .A1(n4024), .A2(n_T_427[897]), .A3(n4018), .A4(
        n_T_427[642]), .Y(n7033) );
  AO22X1_LVT U8360 ( .A1(n3976), .A2(n_T_427[514]), .A3(n4030), .A4(
        n_T_427[833]), .Y(n7032) );
  AO22X1_LVT U8361 ( .A1(n4031), .A2(n_T_427[578]), .A3(n3984), .A4(
        n_T_427[194]), .Y(n7031) );
  NOR4X1_LVT U8362 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .Y(n7040)
         );
  AO22X1_LVT U8363 ( .A1(n3968), .A2(n_T_427[386]), .A3(n3964), .A4(
        n_T_427[258]), .Y(n7038) );
  AO22X1_LVT U8364 ( .A1(n2858), .A2(n_T_427[130]), .A3(n4039), .A4(
        n_T_427[322]), .Y(n7037) );
  AO22X1_LVT U8365 ( .A1(n3979), .A2(n_T_427[769]), .A3(n4045), .A4(
        n_T_427[706]), .Y(n7036) );
  AO22X1_LVT U8366 ( .A1(n3960), .A2(n_T_427[450]), .A3(n4043), .A4(
        n_T_427[66]), .Y(n7035) );
  NOR4X1_LVT U8367 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .Y(n7039)
         );
  NAND2X0_LVT U8368 ( .A1(n3639), .A2(n_T_427[1217]), .Y(n7044) );
  NAND2X0_LVT U8369 ( .A1(n3673), .A2(n_T_427[1089]), .Y(n7046) );
  NAND2X0_LVT U8370 ( .A1(n3712), .A2(n_T_427[961]), .Y(n7045) );
  NAND2X0_LVT U8371 ( .A1(n2967), .A2(n_T_427[1409]), .Y(n7047) );
  OA21X1_LVT U8372 ( .A1(n3196), .A2(n2089), .A3(n7047), .Y(n7050) );
  NAND2X0_LVT U8373 ( .A1(n3609), .A2(n_T_427[1345]), .Y(n7049) );
  NAND2X0_LVT U8374 ( .A1(n3992), .A2(n_T_427[1884]), .Y(n7048) );
  NAND2X0_LVT U8375 ( .A1(n3996), .A2(n_T_427[1282]), .Y(n7051) );
  OA21X1_LVT U8376 ( .A1(n3378), .A2(n3684), .A3(n7051), .Y(n7054) );
  NAND2X0_LVT U8377 ( .A1(n_T_427[1849]), .A2(n3764), .Y(n7053) );
  NAND2X0_LVT U8378 ( .A1(n_T_427[1793]), .A2(n3715), .Y(n7052) );
  NAND2X0_LVT U8379 ( .A1(n3620), .A2(n_T_427[1538]), .Y(n7055) );
  OA21X1_LVT U8380 ( .A1(n3420), .A2(n2897), .A3(n7055), .Y(n7058) );
  NAND2X0_LVT U8381 ( .A1(n4004), .A2(n_T_427[1730]), .Y(n7057) );
  NAND2X0_LVT U8382 ( .A1(n3643), .A2(n_T_427[1602]), .Y(n7056) );
  NAND2X0_LVT U8383 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[3]), .Y(n7071)
         );
  NAND2X0_LVT U8384 ( .A1(n4014), .A2(n_T_427[1026]), .Y(n7070) );
  AND2X1_LVT U8385 ( .A1(n4049), .A2(n_T_427[3]), .Y(n7062) );
  AO22X1_LVT U8386 ( .A1(n4025), .A2(n_T_427[898]), .A3(n4018), .A4(
        n_T_427[643]), .Y(n7061) );
  AO22X1_LVT U8387 ( .A1(n3976), .A2(n_T_427[515]), .A3(n4030), .A4(
        n_T_427[834]), .Y(n7060) );
  AO22X1_LVT U8388 ( .A1(n4032), .A2(n_T_427[579]), .A3(n3983), .A4(
        n_T_427[195]), .Y(n7059) );
  NOR4X1_LVT U8389 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .Y(n7068)
         );
  AO22X1_LVT U8390 ( .A1(n3968), .A2(n_T_427[387]), .A3(n3964), .A4(
        n_T_427[259]), .Y(n7066) );
  AO22X1_LVT U8391 ( .A1(n3975), .A2(n_T_427[131]), .A3(n4038), .A4(
        n_T_427[323]), .Y(n7065) );
  AO22X1_LVT U8392 ( .A1(n3980), .A2(n_T_427[770]), .A3(n4045), .A4(
        n_T_427[707]), .Y(n7064) );
  AO22X1_LVT U8393 ( .A1(n3961), .A2(n_T_427[451]), .A3(n4042), .A4(
        n_T_427[67]), .Y(n7063) );
  NOR4X1_LVT U8394 ( .A1(n7066), .A2(n7065), .A3(n7064), .A4(n7063), .Y(n7067)
         );
  NAND2X0_LVT U8395 ( .A1(n_T_427[1218]), .A2(n3639), .Y(n7072) );
  OA21X1_LVT U8396 ( .A1(n3421), .A2(n3664), .A3(n7072), .Y(n7075) );
  NAND2X0_LVT U8397 ( .A1(n3667), .A2(n_T_427[1090]), .Y(n7074) );
  NAND2X0_LVT U8398 ( .A1(n3759), .A2(n_T_427[962]), .Y(n7073) );
  NAND2X0_LVT U8399 ( .A1(n2966), .A2(n_T_427[1410]), .Y(n7076) );
  OA21X1_LVT U8400 ( .A1(n3187), .A2(n2090), .A3(n7076), .Y(n7079) );
  NAND2X0_LVT U8401 ( .A1(n3602), .A2(n_T_427[1346]), .Y(n7078) );
  NAND2X0_LVT U8402 ( .A1(n2093), .A2(n_T_427[1283]), .Y(n7080) );
  OA21X1_LVT U8403 ( .A1(n3379), .A2(n3684), .A3(n7080), .Y(n7083) );
  NAND2X0_LVT U8404 ( .A1(n_T_427[1850]), .A2(n3990), .Y(n7082) );
  NAND2X0_LVT U8405 ( .A1(n_T_427[1794]), .A2(n3715), .Y(n7081) );
  NAND2X0_LVT U8406 ( .A1(n3615), .A2(n_T_427[1539]), .Y(n7084) );
  OA21X1_LVT U8407 ( .A1(n3422), .A2(n3653), .A3(n7084), .Y(n7087) );
  NAND2X0_LVT U8408 ( .A1(n4003), .A2(n_T_427[1731]), .Y(n7086) );
  NAND2X0_LVT U8409 ( .A1(n3643), .A2(n_T_427[1603]), .Y(n7085) );
  NAND2X0_LVT U8410 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[4]), .Y(n7100)
         );
  NAND2X0_LVT U8411 ( .A1(n3716), .A2(n_T_427[1027]), .Y(n7099) );
  AND2X1_LVT U8412 ( .A1(n4049), .A2(n_T_427[4]), .Y(n7091) );
  AO22X1_LVT U8413 ( .A1(n4026), .A2(n_T_427[899]), .A3(n4018), .A4(
        n_T_427[644]), .Y(n7090) );
  AO22X1_LVT U8414 ( .A1(n3976), .A2(n_T_427[516]), .A3(n4030), .A4(
        n_T_427[835]), .Y(n7089) );
  AO22X1_LVT U8415 ( .A1(n4032), .A2(n_T_427[580]), .A3(n3983), .A4(
        n_T_427[196]), .Y(n7088) );
  NOR4X1_LVT U8416 ( .A1(n7091), .A2(n7090), .A3(n7089), .A4(n7088), .Y(n7097)
         );
  AO22X1_LVT U8417 ( .A1(n3968), .A2(n_T_427[388]), .A3(n3964), .A4(
        n_T_427[260]), .Y(n7095) );
  AO22X1_LVT U8418 ( .A1(n2859), .A2(n_T_427[132]), .A3(n9040), .A4(
        n_T_427[324]), .Y(n7094) );
  AO22X1_LVT U8419 ( .A1(n3980), .A2(n_T_427[771]), .A3(n4045), .A4(
        n_T_427[708]), .Y(n7093) );
  AO22X1_LVT U8420 ( .A1(n3961), .A2(n_T_427[452]), .A3(n4042), .A4(
        n_T_427[68]), .Y(n7092) );
  NOR4X1_LVT U8421 ( .A1(n7095), .A2(n7094), .A3(n7093), .A4(n7092), .Y(n7096)
         );
  NAND3X0_LVT U8422 ( .A1(n7100), .A2(n7099), .A3(n7098), .Y(n7107) );
  NAND2X0_LVT U8423 ( .A1(n3674), .A2(n_T_427[1091]), .Y(n7102) );
  NAND2X0_LVT U8424 ( .A1(n3758), .A2(n_T_427[963]), .Y(n7101) );
  NAND2X0_LVT U8425 ( .A1(n_T_427[1347]), .A2(n3611), .Y(n7104) );
  NAND2X0_LVT U8426 ( .A1(n2986), .A2(n_T_427[1885]), .Y(n7103) );
  OR3X1_LVT U8427 ( .A1(n7108), .A2(n7109), .A3(n7110), .Y(N684) );
  NAND2X0_LVT U8428 ( .A1(n3999), .A2(n_T_427[1284]), .Y(n7111) );
  OA21X1_LVT U8429 ( .A1(n3380), .A2(n3684), .A3(n7111), .Y(n7114) );
  NAND2X0_LVT U8430 ( .A1(n_T_427[1851]), .A2(n3764), .Y(n7113) );
  NAND2X0_LVT U8431 ( .A1(n_T_427[1795]), .A2(n3715), .Y(n7112) );
  NAND2X0_LVT U8432 ( .A1(n3616), .A2(n_T_427[1540]), .Y(n7115) );
  OA21X1_LVT U8433 ( .A1(n3423), .A2(n2897), .A3(n7115), .Y(n7118) );
  NAND2X0_LVT U8434 ( .A1(n4002), .A2(n_T_427[1732]), .Y(n7117) );
  NAND2X0_LVT U8435 ( .A1(n3642), .A2(n_T_427[1604]), .Y(n7116) );
  NAND2X0_LVT U8436 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[5]), .Y(n7131)
         );
  NAND2X0_LVT U8437 ( .A1(n3717), .A2(n_T_427[1028]), .Y(n7130) );
  AND2X1_LVT U8438 ( .A1(n4049), .A2(n_T_427[5]), .Y(n7122) );
  AO22X1_LVT U8439 ( .A1(n4026), .A2(n_T_427[900]), .A3(n4018), .A4(
        n_T_427[645]), .Y(n7121) );
  AO22X1_LVT U8440 ( .A1(n3976), .A2(n_T_427[517]), .A3(n4030), .A4(
        n_T_427[836]), .Y(n7120) );
  AO22X1_LVT U8441 ( .A1(n4032), .A2(n_T_427[581]), .A3(n3984), .A4(
        n_T_427[197]), .Y(n7119) );
  NOR4X1_LVT U8442 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .Y(n7128)
         );
  AO22X1_LVT U8443 ( .A1(n3968), .A2(n_T_427[389]), .A3(n3964), .A4(
        n_T_427[261]), .Y(n7126) );
  AO22X1_LVT U8444 ( .A1(n3974), .A2(n_T_427[133]), .A3(n4037), .A4(
        n_T_427[325]), .Y(n7125) );
  AO22X1_LVT U8445 ( .A1(n3980), .A2(n_T_427[772]), .A3(n4045), .A4(
        n_T_427[709]), .Y(n7124) );
  AO22X1_LVT U8446 ( .A1(n3961), .A2(n_T_427[453]), .A3(n4042), .A4(
        n_T_427[69]), .Y(n7123) );
  NOR4X1_LVT U8447 ( .A1(n7126), .A2(n7125), .A3(n7124), .A4(n7123), .Y(n7127)
         );
  AO21X1_LVT U8448 ( .A1(n7128), .A2(n7127), .A3(n2645), .Y(n7129) );
  NAND2X0_LVT U8449 ( .A1(n3641), .A2(n_T_427[1220]), .Y(n7132) );
  NAND2X0_LVT U8450 ( .A1(n3674), .A2(n_T_427[1092]), .Y(n7134) );
  NAND2X0_LVT U8451 ( .A1(n3756), .A2(n_T_427[964]), .Y(n7133) );
  NAND2X0_LVT U8452 ( .A1(n3629), .A2(n_T_427[1412]), .Y(n7135) );
  OA21X1_LVT U8453 ( .A1(n3197), .A2(n2089), .A3(n7135), .Y(n7138) );
  NAND2X0_LVT U8454 ( .A1(n3608), .A2(n_T_427[1348]), .Y(n7137) );
  NAND2X0_LVT U8455 ( .A1(n2986), .A2(n_T_427[1886]), .Y(n7136) );
  NAND2X0_LVT U8456 ( .A1(n4000), .A2(n_T_427[1285]), .Y(n7139) );
  OA21X1_LVT U8457 ( .A1(n3381), .A2(n3684), .A3(n7139), .Y(n7142) );
  NAND2X0_LVT U8458 ( .A1(n_T_427[1852]), .A2(n3990), .Y(n7141) );
  NAND2X0_LVT U8459 ( .A1(n_T_427[1796]), .A2(n3715), .Y(n7140) );
  NAND2X0_LVT U8460 ( .A1(n3617), .A2(n_T_427[1541]), .Y(n7143) );
  OA21X1_LVT U8461 ( .A1(n3425), .A2(n3653), .A3(n7143), .Y(n7146) );
  NAND2X0_LVT U8462 ( .A1(n4002), .A2(n_T_427[1733]), .Y(n7145) );
  NAND2X0_LVT U8463 ( .A1(n3651), .A2(n_T_427[1605]), .Y(n7144) );
  NAND2X0_LVT U8464 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[6]), .Y(n7159)
         );
  NAND2X0_LVT U8465 ( .A1(n4014), .A2(n_T_427[1029]), .Y(n7158) );
  AND2X1_LVT U8466 ( .A1(n4049), .A2(n_T_427[6]), .Y(n7150) );
  AO22X1_LVT U8467 ( .A1(n4023), .A2(n_T_427[901]), .A3(n4018), .A4(
        n_T_427[646]), .Y(n7149) );
  AO22X1_LVT U8468 ( .A1(n3977), .A2(n_T_427[518]), .A3(n4030), .A4(
        n_T_427[837]), .Y(n7148) );
  AO22X1_LVT U8469 ( .A1(n4032), .A2(n_T_427[582]), .A3(n3983), .A4(
        n_T_427[198]), .Y(n7147) );
  NOR4X1_LVT U8470 ( .A1(n7150), .A2(n7149), .A3(n7148), .A4(n7147), .Y(n7156)
         );
  AO22X1_LVT U8471 ( .A1(n3968), .A2(n_T_427[390]), .A3(n3964), .A4(
        n_T_427[262]), .Y(n7154) );
  AO22X1_LVT U8472 ( .A1(n2859), .A2(n_T_427[134]), .A3(n4039), .A4(
        n_T_427[326]), .Y(n7153) );
  AO22X1_LVT U8473 ( .A1(n3980), .A2(n_T_427[773]), .A3(n4045), .A4(
        n_T_427[710]), .Y(n7152) );
  AO22X1_LVT U8474 ( .A1(n3961), .A2(n_T_427[454]), .A3(n4041), .A4(
        n_T_427[70]), .Y(n7151) );
  NOR4X1_LVT U8475 ( .A1(n7154), .A2(n7153), .A3(n7152), .A4(n7151), .Y(n7155)
         );
  AO21X1_LVT U8476 ( .A1(n7156), .A2(n7155), .A3(n2154), .Y(n7157) );
  NAND2X0_LVT U8477 ( .A1(n_T_427[1221]), .A2(n3640), .Y(n7160) );
  OA21X1_LVT U8478 ( .A1(n3426), .A2(n2081), .A3(n7160), .Y(n7163) );
  NAND2X0_LVT U8479 ( .A1(n3675), .A2(n_T_427[1093]), .Y(n7162) );
  NAND2X0_LVT U8480 ( .A1(n3760), .A2(n_T_427[965]), .Y(n7161) );
  NAND2X0_LVT U8481 ( .A1(n3629), .A2(n_T_427[1413]), .Y(n7164) );
  OA21X1_LVT U8482 ( .A1(n3194), .A2(n2090), .A3(n7164), .Y(n7167) );
  NAND2X0_LVT U8483 ( .A1(n3605), .A2(n_T_427[1349]), .Y(n7166) );
  NAND2X0_LVT U8484 ( .A1(n2985), .A2(n_T_427[1887]), .Y(n7165) );
  NAND2X0_LVT U8485 ( .A1(n2093), .A2(n_T_427[1286]), .Y(n7168) );
  OA21X1_LVT U8486 ( .A1(n3382), .A2(n3684), .A3(n7168), .Y(n7171) );
  NAND2X0_LVT U8487 ( .A1(n_T_427[1853]), .A2(n3990), .Y(n7170) );
  NAND2X0_LVT U8488 ( .A1(n_T_427[1797]), .A2(n3715), .Y(n7169) );
  NAND2X0_LVT U8489 ( .A1(n3618), .A2(n_T_427[1542]), .Y(n7172) );
  NAND2X0_LVT U8490 ( .A1(n4005), .A2(n_T_427[1734]), .Y(n7174) );
  NAND2X0_LVT U8491 ( .A1(n3651), .A2(n_T_427[1606]), .Y(n7173) );
  NAND2X0_LVT U8492 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[7]), .Y(n7187)
         );
  NAND2X0_LVT U8493 ( .A1(n3717), .A2(n_T_427[1030]), .Y(n7186) );
  AND2X1_LVT U8494 ( .A1(n4049), .A2(n_T_427[7]), .Y(n7178) );
  AO22X1_LVT U8495 ( .A1(n4026), .A2(n_T_427[902]), .A3(n4018), .A4(
        n_T_427[647]), .Y(n7177) );
  AO22X1_LVT U8496 ( .A1(n3977), .A2(n_T_427[519]), .A3(n4030), .A4(
        n_T_427[838]), .Y(n7176) );
  AO22X1_LVT U8497 ( .A1(n4032), .A2(n_T_427[583]), .A3(n3983), .A4(
        n_T_427[199]), .Y(n7175) );
  NOR4X1_LVT U8498 ( .A1(n7178), .A2(n7177), .A3(n7176), .A4(n7175), .Y(n7184)
         );
  AO22X1_LVT U8499 ( .A1(n3968), .A2(n_T_427[391]), .A3(n3964), .A4(
        n_T_427[263]), .Y(n7182) );
  AO22X1_LVT U8500 ( .A1(n3975), .A2(n_T_427[135]), .A3(n4037), .A4(
        n_T_427[327]), .Y(n7181) );
  AO22X1_LVT U8501 ( .A1(n3980), .A2(n_T_427[774]), .A3(n4045), .A4(
        n_T_427[711]), .Y(n7180) );
  AO22X1_LVT U8502 ( .A1(n3961), .A2(n_T_427[455]), .A3(n4043), .A4(
        n_T_427[71]), .Y(n7179) );
  NOR4X1_LVT U8503 ( .A1(n7182), .A2(n7181), .A3(n7180), .A4(n7179), .Y(n7183)
         );
  AO21X1_LVT U8504 ( .A1(n7184), .A2(n7183), .A3(n3631), .Y(n7185) );
  NAND2X0_LVT U8505 ( .A1(n_T_427[1222]), .A2(n3638), .Y(n7188) );
  NAND2X0_LVT U8506 ( .A1(n3667), .A2(n_T_427[1094]), .Y(n7190) );
  NAND2X0_LVT U8507 ( .A1(n3756), .A2(n_T_427[966]), .Y(n7189) );
  NAND2X0_LVT U8508 ( .A1(n2967), .A2(n_T_427[1414]), .Y(n7191) );
  NAND2X0_LVT U8509 ( .A1(n3607), .A2(n_T_427[1350]), .Y(n7193) );
  NAND2X0_LVT U8510 ( .A1(n2985), .A2(n_T_427[1888]), .Y(n7192) );
  NAND2X0_LVT U8511 ( .A1(n4000), .A2(n_T_427[1287]), .Y(n7194) );
  OA21X1_LVT U8512 ( .A1(n3383), .A2(n3684), .A3(n7194), .Y(n7197) );
  NAND2X0_LVT U8513 ( .A1(n_T_427[1854]), .A2(n3764), .Y(n7196) );
  NAND2X0_LVT U8514 ( .A1(n_T_427[1798]), .A2(n3715), .Y(n7195) );
  NAND2X0_LVT U8515 ( .A1(n3619), .A2(n_T_427[1543]), .Y(n7198) );
  OA21X1_LVT U8516 ( .A1(n3429), .A2(n2897), .A3(n7198), .Y(n7201) );
  NAND2X0_LVT U8517 ( .A1(n4001), .A2(n_T_427[1735]), .Y(n7200) );
  NAND2X0_LVT U8518 ( .A1(n3643), .A2(n_T_427[1607]), .Y(n7199) );
  NAND2X0_LVT U8519 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[8]), .Y(n7214)
         );
  NAND2X0_LVT U8520 ( .A1(n3716), .A2(n_T_427[1031]), .Y(n7213) );
  AND2X1_LVT U8521 ( .A1(n4049), .A2(n_T_427[8]), .Y(n7205) );
  AO22X1_LVT U8522 ( .A1(n4026), .A2(n_T_427[903]), .A3(n4018), .A4(
        n_T_427[648]), .Y(n7204) );
  AO22X1_LVT U8523 ( .A1(n3977), .A2(n_T_427[520]), .A3(n4030), .A4(
        n_T_427[839]), .Y(n7203) );
  AO22X1_LVT U8524 ( .A1(n4032), .A2(n_T_427[584]), .A3(n3983), .A4(
        n_T_427[200]), .Y(n7202) );
  NOR4X1_LVT U8525 ( .A1(n7205), .A2(n7204), .A3(n7203), .A4(n7202), .Y(n7211)
         );
  AO22X1_LVT U8526 ( .A1(n3968), .A2(n_T_427[392]), .A3(n3964), .A4(
        n_T_427[264]), .Y(n7209) );
  AO22X1_LVT U8527 ( .A1(n3974), .A2(n_T_427[136]), .A3(n4039), .A4(
        n_T_427[328]), .Y(n7208) );
  AO22X1_LVT U8528 ( .A1(n3980), .A2(n_T_427[775]), .A3(n4045), .A4(
        n_T_427[712]), .Y(n7207) );
  AO22X1_LVT U8529 ( .A1(n3961), .A2(n_T_427[456]), .A3(n4044), .A4(
        n_T_427[72]), .Y(n7206) );
  NOR4X1_LVT U8530 ( .A1(n7209), .A2(n7208), .A3(n7207), .A4(n7206), .Y(n7210)
         );
  AO21X1_LVT U8531 ( .A1(n7211), .A2(n7210), .A3(n3656), .Y(n7212) );
  NAND2X0_LVT U8532 ( .A1(n3637), .A2(n_T_427[1223]), .Y(n7215) );
  OA21X1_LVT U8533 ( .A1(n3430), .A2(n4010), .A3(n7215), .Y(n7218) );
  NAND2X0_LVT U8534 ( .A1(n3675), .A2(n_T_427[1095]), .Y(n7217) );
  NAND2X0_LVT U8535 ( .A1(n3756), .A2(n_T_427[967]), .Y(n7216) );
  NAND2X0_LVT U8536 ( .A1(n3629), .A2(n_T_427[1415]), .Y(n7219) );
  OA21X1_LVT U8537 ( .A1(n3192), .A2(n2089), .A3(n7219), .Y(n7222) );
  NAND2X0_LVT U8538 ( .A1(n3608), .A2(n_T_427[1351]), .Y(n7221) );
  NAND2X0_LVT U8539 ( .A1(n2986), .A2(n_T_427[1889]), .Y(n7220) );
  NAND2X0_LVT U8540 ( .A1(n2093), .A2(n_T_427[1288]), .Y(n7223) );
  OA21X1_LVT U8541 ( .A1(n3384), .A2(n3684), .A3(n7223), .Y(n7226) );
  NAND2X0_LVT U8542 ( .A1(n_T_427[1855]), .A2(n3990), .Y(n7225) );
  NAND2X0_LVT U8543 ( .A1(n_T_427[1799]), .A2(n3715), .Y(n7224) );
  NAND2X0_LVT U8544 ( .A1(n3620), .A2(n_T_427[1544]), .Y(n7227) );
  OA21X1_LVT U8545 ( .A1(n3431), .A2(n2897), .A3(n7227), .Y(n7230) );
  NAND2X0_LVT U8546 ( .A1(n4001), .A2(n_T_427[1736]), .Y(n7229) );
  NAND2X0_LVT U8547 ( .A1(n3652), .A2(n_T_427[1608]), .Y(n7228) );
  NAND2X0_LVT U8548 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[9]), .Y(n7243)
         );
  NAND2X0_LVT U8549 ( .A1(n4014), .A2(n_T_427[1032]), .Y(n7242) );
  AND2X1_LVT U8550 ( .A1(n4049), .A2(n_T_427[9]), .Y(n7234) );
  AO22X1_LVT U8551 ( .A1(n4026), .A2(n_T_427[904]), .A3(n4019), .A4(
        n_T_427[649]), .Y(n7233) );
  AO22X1_LVT U8552 ( .A1(n3977), .A2(n_T_427[521]), .A3(n4029), .A4(
        n_T_427[840]), .Y(n7232) );
  AO22X1_LVT U8553 ( .A1(n4032), .A2(n_T_427[585]), .A3(n3984), .A4(
        n_T_427[201]), .Y(n7231) );
  NOR4X1_LVT U8554 ( .A1(n7234), .A2(n7233), .A3(n7232), .A4(n7231), .Y(n7240)
         );
  AO22X1_LVT U8555 ( .A1(n3969), .A2(n_T_427[393]), .A3(n3965), .A4(
        n_T_427[265]), .Y(n7238) );
  AO22X1_LVT U8556 ( .A1(n3975), .A2(n_T_427[137]), .A3(n4039), .A4(
        n_T_427[329]), .Y(n7237) );
  AO22X1_LVT U8557 ( .A1(n3980), .A2(n_T_427[776]), .A3(n4045), .A4(
        n_T_427[713]), .Y(n7236) );
  AO22X1_LVT U8558 ( .A1(n3961), .A2(n_T_427[457]), .A3(n2837), .A4(
        n_T_427[73]), .Y(n7235) );
  NOR4X1_LVT U8559 ( .A1(n7238), .A2(n7237), .A3(n7236), .A4(n7235), .Y(n7239)
         );
  AO21X1_LVT U8560 ( .A1(n7240), .A2(n7239), .A3(n2155), .Y(n7241) );
  NAND2X0_LVT U8561 ( .A1(n3636), .A2(n_T_427[1224]), .Y(n7244) );
  NAND2X0_LVT U8562 ( .A1(n3672), .A2(n_T_427[1096]), .Y(n7246) );
  NAND2X0_LVT U8563 ( .A1(n3761), .A2(n_T_427[968]), .Y(n7245) );
  NAND2X0_LVT U8564 ( .A1(n3626), .A2(n_T_427[1416]), .Y(n7247) );
  NAND2X0_LVT U8565 ( .A1(n2882), .A2(n_T_427[1890]), .Y(n7248) );
  NAND2X0_LVT U8566 ( .A1(n3998), .A2(n_T_427[1289]), .Y(n7249) );
  OA21X1_LVT U8567 ( .A1(n3385), .A2(n3684), .A3(n7249), .Y(n7252) );
  NAND2X0_LVT U8568 ( .A1(n_T_427[1856]), .A2(n3764), .Y(n7251) );
  NAND2X0_LVT U8569 ( .A1(n_T_427[1800]), .A2(n3715), .Y(n7250) );
  NAND2X0_LVT U8570 ( .A1(n3621), .A2(n_T_427[1545]), .Y(n7253) );
  OA21X1_LVT U8571 ( .A1(n3433), .A2(n3653), .A3(n7253), .Y(n7256) );
  NAND2X0_LVT U8572 ( .A1(n2091), .A2(n_T_427[1737]), .Y(n7255) );
  NAND2X0_LVT U8573 ( .A1(n3648), .A2(n_T_427[1609]), .Y(n7254) );
  NAND2X0_LVT U8574 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[10]), .Y(n7269)
         );
  NAND2X0_LVT U8575 ( .A1(n3717), .A2(n_T_427[1033]), .Y(n7268) );
  AND2X1_LVT U8576 ( .A1(n4049), .A2(n_T_427[10]), .Y(n7260) );
  AO22X1_LVT U8577 ( .A1(n4026), .A2(n_T_427[905]), .A3(n4018), .A4(
        n_T_427[650]), .Y(n7259) );
  AO22X1_LVT U8578 ( .A1(n3977), .A2(n_T_427[522]), .A3(n4029), .A4(
        n_T_427[841]), .Y(n7258) );
  AO22X1_LVT U8579 ( .A1(n4032), .A2(n_T_427[586]), .A3(n3984), .A4(
        n_T_427[202]), .Y(n7257) );
  NOR4X1_LVT U8580 ( .A1(n7260), .A2(n7259), .A3(n7258), .A4(n7257), .Y(n7266)
         );
  AO22X1_LVT U8581 ( .A1(n3968), .A2(n_T_427[394]), .A3(n3964), .A4(
        n_T_427[266]), .Y(n7264) );
  AO22X1_LVT U8582 ( .A1(n3973), .A2(n_T_427[138]), .A3(n4039), .A4(
        n_T_427[330]), .Y(n7263) );
  AO22X1_LVT U8583 ( .A1(n3980), .A2(n_T_427[777]), .A3(n4045), .A4(
        n_T_427[714]), .Y(n7262) );
  AO22X1_LVT U8584 ( .A1(n3961), .A2(n_T_427[458]), .A3(n2836), .A4(
        n_T_427[74]), .Y(n7261) );
  NOR4X1_LVT U8585 ( .A1(n7264), .A2(n7263), .A3(n7262), .A4(n7261), .Y(n7265)
         );
  AO21X1_LVT U8586 ( .A1(n7266), .A2(n7265), .A3(n2645), .Y(n7267) );
  NAND2X0_LVT U8587 ( .A1(n3637), .A2(n_T_427[1225]), .Y(n7270) );
  OA21X1_LVT U8588 ( .A1(n3434), .A2(n3664), .A3(n7270), .Y(n7273) );
  NAND2X0_LVT U8589 ( .A1(n3671), .A2(n_T_427[1097]), .Y(n7272) );
  NAND2X0_LVT U8590 ( .A1(n3757), .A2(n_T_427[969]), .Y(n7271) );
  NAND2X0_LVT U8591 ( .A1(n2966), .A2(n_T_427[1417]), .Y(n7274) );
  OA21X1_LVT U8592 ( .A1(n3188), .A2(n2090), .A3(n7274), .Y(n7277) );
  NAND2X0_LVT U8593 ( .A1(n3602), .A2(n_T_427[1353]), .Y(n7276) );
  NAND2X0_LVT U8594 ( .A1(n2998), .A2(n_T_427[1891]), .Y(n7275) );
  NAND2X0_LVT U8595 ( .A1(n4000), .A2(n_T_427[1290]), .Y(n7278) );
  OA21X1_LVT U8596 ( .A1(n3435), .A2(n3684), .A3(n7278), .Y(n7281) );
  NAND2X0_LVT U8597 ( .A1(n_T_427[1857]), .A2(n3764), .Y(n7280) );
  NAND2X0_LVT U8598 ( .A1(n_T_427[1801]), .A2(n3715), .Y(n7279) );
  NAND2X0_LVT U8599 ( .A1(n3619), .A2(n_T_427[1546]), .Y(n7282) );
  OA21X1_LVT U8600 ( .A1(n3386), .A2(n3653), .A3(n7282), .Y(n7285) );
  NAND2X0_LVT U8601 ( .A1(n2092), .A2(n_T_427[1738]), .Y(n7284) );
  NAND2X0_LVT U8602 ( .A1(n3642), .A2(n_T_427[1610]), .Y(n7283) );
  NAND2X0_LVT U8603 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[11]), .Y(n7298)
         );
  NAND2X0_LVT U8604 ( .A1(n4014), .A2(n_T_427[1034]), .Y(n7297) );
  AND2X1_LVT U8605 ( .A1(n4049), .A2(n_T_427[11]), .Y(n7289) );
  AO22X1_LVT U8606 ( .A1(n4026), .A2(n_T_427[906]), .A3(n4019), .A4(
        n_T_427[651]), .Y(n7288) );
  AO22X1_LVT U8607 ( .A1(n3977), .A2(n_T_427[523]), .A3(n4029), .A4(
        n_T_427[842]), .Y(n7287) );
  AO22X1_LVT U8608 ( .A1(n4032), .A2(n_T_427[587]), .A3(n3984), .A4(
        n_T_427[203]), .Y(n7286) );
  NOR4X1_LVT U8609 ( .A1(n7289), .A2(n7288), .A3(n7287), .A4(n7286), .Y(n7295)
         );
  AO22X1_LVT U8610 ( .A1(n3969), .A2(n_T_427[395]), .A3(n3964), .A4(
        n_T_427[267]), .Y(n7293) );
  AO22X1_LVT U8611 ( .A1(n3973), .A2(n_T_427[139]), .A3(n4037), .A4(
        n_T_427[331]), .Y(n7292) );
  AO22X1_LVT U8612 ( .A1(n3980), .A2(n_T_427[778]), .A3(n4045), .A4(
        n_T_427[715]), .Y(n7291) );
  AO22X1_LVT U8613 ( .A1(n3961), .A2(n_T_427[459]), .A3(n4042), .A4(
        n_T_427[75]), .Y(n7290) );
  NOR4X1_LVT U8614 ( .A1(n7293), .A2(n7292), .A3(n7291), .A4(n7290), .Y(n7294)
         );
  AO21X1_LVT U8615 ( .A1(n7295), .A2(n7294), .A3(n3631), .Y(n7296) );
  NAND2X0_LVT U8616 ( .A1(n3667), .A2(n_T_427[1098]), .Y(n7300) );
  NAND2X0_LVT U8617 ( .A1(n3758), .A2(n_T_427[970]), .Y(n7299) );
  NAND2X0_LVT U8618 ( .A1(n3630), .A2(n_T_427[1418]), .Y(n7302) );
  NAND2X0_LVT U8619 ( .A1(n3603), .A2(n_T_427[1354]), .Y(n7304) );
  NAND2X0_LVT U8620 ( .A1(n2985), .A2(n_T_427[1892]), .Y(n7303) );
  NAND2X0_LVT U8621 ( .A1(n2093), .A2(n_T_427[1291]), .Y(n7305) );
  OA21X1_LVT U8622 ( .A1(n3387), .A2(n3684), .A3(n7305), .Y(n7308) );
  NAND2X0_LVT U8623 ( .A1(n_T_427[1858]), .A2(n3990), .Y(n7307) );
  NAND2X0_LVT U8624 ( .A1(n_T_427[1802]), .A2(n3995), .Y(n7306) );
  NAND2X0_LVT U8625 ( .A1(n3615), .A2(n_T_427[1547]), .Y(n7309) );
  OA21X1_LVT U8626 ( .A1(n3436), .A2(n2897), .A3(n7309), .Y(n7312) );
  NAND2X0_LVT U8627 ( .A1(n4005), .A2(n_T_427[1739]), .Y(n7311) );
  NAND2X0_LVT U8628 ( .A1(n3648), .A2(n_T_427[1611]), .Y(n7310) );
  NAND2X0_LVT U8629 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[12]), .Y(n7325)
         );
  NAND2X0_LVT U8630 ( .A1(n3716), .A2(n_T_427[1035]), .Y(n7324) );
  AND2X1_LVT U8631 ( .A1(n4049), .A2(n_T_427[12]), .Y(n7316) );
  AO22X1_LVT U8632 ( .A1(n4026), .A2(n_T_427[907]), .A3(n4019), .A4(
        n_T_427[652]), .Y(n7315) );
  AO22X1_LVT U8633 ( .A1(n3977), .A2(n_T_427[524]), .A3(n4029), .A4(
        n_T_427[843]), .Y(n7314) );
  AO22X1_LVT U8634 ( .A1(n4032), .A2(n_T_427[588]), .A3(n3984), .A4(
        n_T_427[204]), .Y(n7313) );
  NOR4X1_LVT U8635 ( .A1(n7316), .A2(n7315), .A3(n7314), .A4(n7313), .Y(n7322)
         );
  AO22X1_LVT U8636 ( .A1(n3968), .A2(n_T_427[396]), .A3(n3965), .A4(
        n_T_427[268]), .Y(n7320) );
  AO22X1_LVT U8637 ( .A1(n3973), .A2(n_T_427[140]), .A3(n4036), .A4(
        n_T_427[332]), .Y(n7319) );
  AO22X1_LVT U8638 ( .A1(n3980), .A2(n_T_427[779]), .A3(n4046), .A4(
        n_T_427[716]), .Y(n7318) );
  AO22X1_LVT U8639 ( .A1(n3961), .A2(n_T_427[460]), .A3(n4044), .A4(
        n_T_427[76]), .Y(n7317) );
  NOR4X1_LVT U8640 ( .A1(n7320), .A2(n7319), .A3(n7318), .A4(n7317), .Y(n7321)
         );
  NAND2X0_LVT U8641 ( .A1(n_T_427[1227]), .A2(n3640), .Y(n7326) );
  OA21X1_LVT U8642 ( .A1(n3437), .A2(n4008), .A3(n7326), .Y(n7329) );
  NAND2X0_LVT U8643 ( .A1(n3674), .A2(n_T_427[1099]), .Y(n7328) );
  NAND2X0_LVT U8644 ( .A1(n3761), .A2(n_T_427[971]), .Y(n7327) );
  NAND2X0_LVT U8645 ( .A1(n2966), .A2(n_T_427[1419]), .Y(n7330) );
  OA21X1_LVT U8646 ( .A1(n3193), .A2(n2089), .A3(n7330), .Y(n7333) );
  NAND2X0_LVT U8647 ( .A1(n3604), .A2(n_T_427[1355]), .Y(n7332) );
  NAND2X0_LVT U8648 ( .A1(n2986), .A2(n_T_427[1893]), .Y(n7331) );
  NAND2X0_LVT U8649 ( .A1(n2094), .A2(n_T_427[1292]), .Y(n7334) );
  OA21X1_LVT U8650 ( .A1(n3388), .A2(n3684), .A3(n7334), .Y(n7337) );
  NAND2X0_LVT U8651 ( .A1(n_T_427[1859]), .A2(n3990), .Y(n7336) );
  NAND2X0_LVT U8652 ( .A1(n_T_427[1803]), .A2(n3995), .Y(n7335) );
  NAND2X0_LVT U8653 ( .A1(n3616), .A2(n_T_427[1548]), .Y(n7338) );
  OA21X1_LVT U8654 ( .A1(n3438), .A2(n3653), .A3(n7338), .Y(n7341) );
  NAND2X0_LVT U8655 ( .A1(n2092), .A2(n_T_427[1740]), .Y(n7340) );
  NAND2X0_LVT U8656 ( .A1(n3652), .A2(n_T_427[1612]), .Y(n7339) );
  NAND2X0_LVT U8657 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[13]), .Y(n7354)
         );
  NAND2X0_LVT U8658 ( .A1(n3716), .A2(n_T_427[1036]), .Y(n7353) );
  AND2X1_LVT U8659 ( .A1(n4050), .A2(n_T_427[13]), .Y(n7345) );
  AO22X1_LVT U8660 ( .A1(n4026), .A2(n_T_427[908]), .A3(n4019), .A4(
        n_T_427[653]), .Y(n7344) );
  AO22X1_LVT U8661 ( .A1(n3977), .A2(n_T_427[525]), .A3(n4029), .A4(
        n_T_427[844]), .Y(n7343) );
  AO22X1_LVT U8662 ( .A1(n4032), .A2(n_T_427[589]), .A3(n3984), .A4(
        n_T_427[205]), .Y(n7342) );
  NOR4X1_LVT U8663 ( .A1(n7345), .A2(n7344), .A3(n7343), .A4(n7342), .Y(n7351)
         );
  AO22X1_LVT U8664 ( .A1(n3969), .A2(n_T_427[397]), .A3(n3965), .A4(
        n_T_427[269]), .Y(n7349) );
  AO22X1_LVT U8665 ( .A1(n3974), .A2(n_T_427[141]), .A3(n4037), .A4(
        n_T_427[333]), .Y(n7348) );
  AO22X1_LVT U8666 ( .A1(n3980), .A2(n_T_427[780]), .A3(n4046), .A4(
        n_T_427[717]), .Y(n7347) );
  AO22X1_LVT U8667 ( .A1(n3961), .A2(n_T_427[461]), .A3(n2836), .A4(
        n_T_427[77]), .Y(n7346) );
  NOR4X1_LVT U8668 ( .A1(n7349), .A2(n7348), .A3(n7347), .A4(n7346), .Y(n7350)
         );
  NAND2X0_LVT U8669 ( .A1(n_T_427[1228]), .A2(n3638), .Y(n7355) );
  NAND2X0_LVT U8670 ( .A1(n_T_427[1100]), .A2(n3674), .Y(n7357) );
  NAND2X0_LVT U8671 ( .A1(n3757), .A2(n_T_427[972]), .Y(n7356) );
  NAND2X0_LVT U8672 ( .A1(n3610), .A2(n_T_427[1356]), .Y(n7359) );
  NAND2X0_LVT U8673 ( .A1(n2998), .A2(n_T_427[1894]), .Y(n7358) );
  NAND2X0_LVT U8674 ( .A1(n3998), .A2(n_T_427[1293]), .Y(n7361) );
  OA21X1_LVT U8675 ( .A1(n3389), .A2(n3684), .A3(n7361), .Y(n7364) );
  NAND2X0_LVT U8676 ( .A1(n_T_427[1860]), .A2(n3990), .Y(n7363) );
  NAND2X0_LVT U8677 ( .A1(n_T_427[1804]), .A2(n3995), .Y(n7362) );
  NAND2X0_LVT U8678 ( .A1(n3617), .A2(n_T_427[1549]), .Y(n7365) );
  OA21X1_LVT U8679 ( .A1(n3440), .A2(n2897), .A3(n7365), .Y(n7368) );
  NAND2X0_LVT U8680 ( .A1(n4001), .A2(n_T_427[1741]), .Y(n7367) );
  NAND2X0_LVT U8681 ( .A1(n3651), .A2(n_T_427[1613]), .Y(n7366) );
  NAND2X0_LVT U8682 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[14]), .Y(n7381)
         );
  NAND2X0_LVT U8683 ( .A1(n3716), .A2(n_T_427[1037]), .Y(n7380) );
  AND2X1_LVT U8684 ( .A1(n4050), .A2(n_T_427[14]), .Y(n7372) );
  AO22X1_LVT U8685 ( .A1(n4026), .A2(n_T_427[909]), .A3(n4019), .A4(
        n_T_427[654]), .Y(n7371) );
  AO22X1_LVT U8686 ( .A1(n3977), .A2(n_T_427[526]), .A3(n4029), .A4(
        n_T_427[845]), .Y(n7370) );
  AO22X1_LVT U8687 ( .A1(n4032), .A2(n_T_427[590]), .A3(n3984), .A4(
        n_T_427[206]), .Y(n7369) );
  NOR4X1_LVT U8688 ( .A1(n7372), .A2(n7371), .A3(n7370), .A4(n7369), .Y(n7378)
         );
  AO22X1_LVT U8689 ( .A1(n3969), .A2(n_T_427[398]), .A3(n3965), .A4(
        n_T_427[270]), .Y(n7376) );
  AO22X1_LVT U8690 ( .A1(n2859), .A2(n_T_427[142]), .A3(n4036), .A4(
        n_T_427[334]), .Y(n7375) );
  AO22X1_LVT U8691 ( .A1(n3980), .A2(n_T_427[781]), .A3(n4046), .A4(
        n_T_427[718]), .Y(n7374) );
  AO22X1_LVT U8692 ( .A1(n3961), .A2(n_T_427[462]), .A3(n2837), .A4(
        n_T_427[78]), .Y(n7373) );
  NOR4X1_LVT U8693 ( .A1(n7376), .A2(n7375), .A3(n7374), .A4(n7373), .Y(n7377)
         );
  NAND2X0_LVT U8694 ( .A1(n_T_427[1229]), .A2(n3636), .Y(n7382) );
  OA21X1_LVT U8695 ( .A1(n3441), .A2(n3664), .A3(n7382), .Y(n7385) );
  NAND2X0_LVT U8696 ( .A1(n3673), .A2(n_T_427[1101]), .Y(n7384) );
  NAND2X0_LVT U8697 ( .A1(n3758), .A2(n_T_427[973]), .Y(n7383) );
  NAND2X0_LVT U8698 ( .A1(n3629), .A2(n_T_427[1421]), .Y(n7386) );
  OA21X1_LVT U8699 ( .A1(n3195), .A2(n2089), .A3(n7386), .Y(n7389) );
  NAND2X0_LVT U8700 ( .A1(n3604), .A2(n_T_427[1357]), .Y(n7388) );
  NAND2X0_LVT U8701 ( .A1(n3992), .A2(n_T_427[1895]), .Y(n7387) );
  NAND2X0_LVT U8702 ( .A1(n3996), .A2(n_T_427[1294]), .Y(n7390) );
  OA21X1_LVT U8703 ( .A1(n3390), .A2(n3684), .A3(n7390), .Y(n7393) );
  NAND2X0_LVT U8704 ( .A1(n_T_427[1861]), .A2(n3764), .Y(n7392) );
  NAND2X0_LVT U8705 ( .A1(n_T_427[1805]), .A2(n3995), .Y(n7391) );
  NAND2X0_LVT U8706 ( .A1(n3618), .A2(n_T_427[1550]), .Y(n7394) );
  OA21X1_LVT U8707 ( .A1(n3442), .A2(n3653), .A3(n7394), .Y(n7397) );
  NAND2X0_LVT U8708 ( .A1(n4005), .A2(n_T_427[1742]), .Y(n7396) );
  NAND2X0_LVT U8709 ( .A1(n3649), .A2(n_T_427[1614]), .Y(n7395) );
  NAND2X0_LVT U8710 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[15]), .Y(n7410)
         );
  NAND2X0_LVT U8711 ( .A1(n3716), .A2(n_T_427[1038]), .Y(n7409) );
  AND2X1_LVT U8712 ( .A1(n4050), .A2(n_T_427[15]), .Y(n7401) );
  AO22X1_LVT U8713 ( .A1(n4026), .A2(n_T_427[910]), .A3(n4019), .A4(
        n_T_427[655]), .Y(n7400) );
  AO22X1_LVT U8714 ( .A1(n3977), .A2(n_T_427[527]), .A3(n4029), .A4(
        n_T_427[846]), .Y(n7399) );
  AO22X1_LVT U8715 ( .A1(n4033), .A2(n_T_427[591]), .A3(n3984), .A4(
        n_T_427[207]), .Y(n7398) );
  NOR4X1_LVT U8716 ( .A1(n7401), .A2(n7400), .A3(n7399), .A4(n7398), .Y(n7407)
         );
  AO22X1_LVT U8717 ( .A1(n3969), .A2(n_T_427[399]), .A3(n3965), .A4(
        n_T_427[271]), .Y(n7405) );
  AO22X1_LVT U8718 ( .A1(n3973), .A2(n_T_427[143]), .A3(n4039), .A4(
        n_T_427[335]), .Y(n7404) );
  AO22X1_LVT U8719 ( .A1(n3980), .A2(n_T_427[782]), .A3(n4046), .A4(
        n_T_427[719]), .Y(n7403) );
  AO22X1_LVT U8720 ( .A1(n3961), .A2(n_T_427[463]), .A3(n4043), .A4(
        n_T_427[79]), .Y(n7402) );
  NOR4X1_LVT U8721 ( .A1(n7405), .A2(n7404), .A3(n7403), .A4(n7402), .Y(n7406)
         );
  AO21X1_LVT U8722 ( .A1(n7407), .A2(n7406), .A3(n3632), .Y(n7408) );
  NAND2X0_LVT U8723 ( .A1(n3641), .A2(n_T_427[1230]), .Y(n7411) );
  NAND2X0_LVT U8724 ( .A1(n3673), .A2(n_T_427[1102]), .Y(n7413) );
  NAND2X0_LVT U8725 ( .A1(n3756), .A2(n_T_427[974]), .Y(n7412) );
  NAND2X0_LVT U8726 ( .A1(n3627), .A2(n_T_427[1422]), .Y(n7414) );
  NAND2X0_LVT U8727 ( .A1(n3607), .A2(n_T_427[1358]), .Y(n7416) );
  NAND2X0_LVT U8728 ( .A1(n2985), .A2(n_T_427[1896]), .Y(n7415) );
  NAND2X0_LVT U8729 ( .A1(n2093), .A2(n_T_427[1295]), .Y(n7417) );
  OA21X1_LVT U8730 ( .A1(n3444), .A2(n3601), .A3(n7417), .Y(n7420) );
  NAND2X0_LVT U8731 ( .A1(n3744), .A2(n_T_427[1679]), .Y(n7419) );
  NAND2X0_LVT U8732 ( .A1(n4005), .A2(n_T_427[1743]), .Y(n7418) );
  NAND2X0_LVT U8733 ( .A1(n3619), .A2(n_T_427[1551]), .Y(n7421) );
  OA21X1_LVT U8734 ( .A1(n3664), .A2(n3312), .A3(n7421), .Y(n7424) );
  NAND2X0_LVT U8735 ( .A1(n3649), .A2(n_T_427[1615]), .Y(n7423) );
  NAND2X0_LVT U8736 ( .A1(n4006), .A2(n_T_427[1487]), .Y(n7422) );
  NAND2X0_LVT U8737 ( .A1(n3757), .A2(n_T_427[975]), .Y(n7425) );
  NAND2X0_LVT U8738 ( .A1(n3636), .A2(n_T_427[1231]), .Y(n7427) );
  NAND2X0_LVT U8739 ( .A1(n3667), .A2(n_T_427[1103]), .Y(n7426) );
  NAND2X0_LVT U8740 ( .A1(n2966), .A2(n_T_427[1423]), .Y(n7429) );
  NAND2X0_LVT U8741 ( .A1(n3608), .A2(n_T_427[1359]), .Y(n7428) );
  AND2X1_LVT U8742 ( .A1(n4050), .A2(n_T_427[16]), .Y(n7433) );
  AO22X1_LVT U8743 ( .A1(n4026), .A2(n_T_427[911]), .A3(n4019), .A4(
        n_T_427[656]), .Y(n7432) );
  AO22X1_LVT U8744 ( .A1(n3977), .A2(n_T_427[528]), .A3(n4029), .A4(
        n_T_427[847]), .Y(n7431) );
  AO22X1_LVT U8745 ( .A1(n4032), .A2(n_T_427[592]), .A3(n3984), .A4(
        n_T_427[208]), .Y(n7430) );
  NOR4X1_LVT U8746 ( .A1(n7433), .A2(n7432), .A3(n7431), .A4(n7430), .Y(n7439)
         );
  AO22X1_LVT U8747 ( .A1(n3969), .A2(n_T_427[400]), .A3(n3965), .A4(
        n_T_427[272]), .Y(n7437) );
  AO22X1_LVT U8748 ( .A1(n3974), .A2(n_T_427[144]), .A3(n4036), .A4(
        n_T_427[336]), .Y(n7436) );
  AO22X1_LVT U8749 ( .A1(n3980), .A2(n_T_427[783]), .A3(n4046), .A4(
        n_T_427[720]), .Y(n7435) );
  AO22X1_LVT U8750 ( .A1(n3961), .A2(n_T_427[464]), .A3(n2836), .A4(
        n_T_427[80]), .Y(n7434) );
  NOR4X1_LVT U8751 ( .A1(n7437), .A2(n7436), .A3(n7435), .A4(n7434), .Y(n7438)
         );
  AO21X1_LVT U8752 ( .A1(n7439), .A2(n7438), .A3(n2154), .Y(n7440) );
  NAND2X0_LVT U8753 ( .A1(n4000), .A2(n_T_427[1296]), .Y(n7443) );
  OA21X1_LVT U8754 ( .A1(n3142), .A2(n3747), .A3(n7443), .Y(n7446) );
  NAND2X0_LVT U8755 ( .A1(n3744), .A2(n_T_427[1680]), .Y(n7445) );
  NAND2X0_LVT U8756 ( .A1(n2092), .A2(n_T_427[1744]), .Y(n7444) );
  NAND2X0_LVT U8757 ( .A1(n3615), .A2(n_T_427[1552]), .Y(n7447) );
  OA21X1_LVT U8758 ( .A1(n4010), .A2(n3313), .A3(n7447), .Y(n7450) );
  NAND2X0_LVT U8759 ( .A1(n3652), .A2(n_T_427[1616]), .Y(n7449) );
  NAND2X0_LVT U8760 ( .A1(n4007), .A2(n_T_427[1488]), .Y(n7448) );
  NAND2X0_LVT U8761 ( .A1(n3758), .A2(n_T_427[976]), .Y(n7451) );
  OA21X1_LVT U8762 ( .A1(n3752), .A2(n3283), .A3(n7451), .Y(n7454) );
  NAND2X0_LVT U8763 ( .A1(n3639), .A2(n_T_427[1232]), .Y(n7453) );
  NAND2X0_LVT U8764 ( .A1(n3669), .A2(n_T_427[1104]), .Y(n7452) );
  NAND2X0_LVT U8765 ( .A1(n3992), .A2(n_T_427[1898]), .Y(n7455) );
  NAND2X0_LVT U8766 ( .A1(n3628), .A2(n_T_427[1424]), .Y(n7457) );
  NAND2X0_LVT U8767 ( .A1(n3605), .A2(n_T_427[1360]), .Y(n7456) );
  NAND2X0_LVT U8768 ( .A1(n3665), .A2(n4367), .Y(n7469) );
  AND2X1_LVT U8769 ( .A1(n4050), .A2(n_T_427[17]), .Y(n7461) );
  AO22X1_LVT U8770 ( .A1(n4025), .A2(n_T_427[912]), .A3(n4019), .A4(
        n_T_427[657]), .Y(n7460) );
  AO22X1_LVT U8771 ( .A1(n3977), .A2(n_T_427[529]), .A3(n4029), .A4(
        n_T_427[848]), .Y(n7459) );
  AO22X1_LVT U8772 ( .A1(n4033), .A2(n_T_427[593]), .A3(n3984), .A4(
        n_T_427[209]), .Y(n7458) );
  NOR4X1_LVT U8773 ( .A1(n7461), .A2(n7460), .A3(n7459), .A4(n7458), .Y(n7467)
         );
  AO22X1_LVT U8774 ( .A1(n3969), .A2(n_T_427[401]), .A3(n3965), .A4(
        n_T_427[273]), .Y(n7465) );
  AO22X1_LVT U8775 ( .A1(n3973), .A2(n_T_427[145]), .A3(n9040), .A4(
        n_T_427[337]), .Y(n7464) );
  AO22X1_LVT U8776 ( .A1(n3981), .A2(n_T_427[784]), .A3(n4046), .A4(
        n_T_427[721]), .Y(n7463) );
  AO22X1_LVT U8777 ( .A1(n3962), .A2(n_T_427[465]), .A3(n4042), .A4(
        n_T_427[81]), .Y(n7462) );
  NOR4X1_LVT U8778 ( .A1(n7465), .A2(n7464), .A3(n7463), .A4(n7462), .Y(n7466)
         );
  NAND2X0_LVT U8779 ( .A1(n3996), .A2(n_T_427[1297]), .Y(n7471) );
  OA21X1_LVT U8780 ( .A1(n3445), .A2(n3601), .A3(n7471), .Y(n7474) );
  NAND2X0_LVT U8781 ( .A1(n3744), .A2(n_T_427[1681]), .Y(n7473) );
  NAND2X0_LVT U8782 ( .A1(n2092), .A2(n_T_427[1745]), .Y(n7472) );
  NAND2X0_LVT U8783 ( .A1(n3620), .A2(n_T_427[1553]), .Y(n7475) );
  OA21X1_LVT U8784 ( .A1(n3663), .A2(n3314), .A3(n7475), .Y(n7478) );
  NAND2X0_LVT U8785 ( .A1(n3649), .A2(n_T_427[1617]), .Y(n7477) );
  NAND2X0_LVT U8786 ( .A1(n4007), .A2(n_T_427[1489]), .Y(n7476) );
  NAND2X0_LVT U8787 ( .A1(n3757), .A2(n_T_427[977]), .Y(n7479) );
  OA21X1_LVT U8788 ( .A1(n3752), .A2(n3315), .A3(n7479), .Y(n7482) );
  NAND2X0_LVT U8789 ( .A1(n3637), .A2(n_T_427[1233]), .Y(n7481) );
  NAND2X0_LVT U8790 ( .A1(n3673), .A2(n_T_427[1105]), .Y(n7480) );
  OA21X1_LVT U8791 ( .A1(n3988), .A2(n3316), .A3(n7483), .Y(n7486) );
  NAND2X0_LVT U8792 ( .A1(n3628), .A2(n_T_427[1425]), .Y(n7485) );
  NAND2X0_LVT U8793 ( .A1(n3602), .A2(n_T_427[1361]), .Y(n7484) );
  NAND2X0_LVT U8794 ( .A1(n4015), .A2(n4370), .Y(n7498) );
  AND2X1_LVT U8795 ( .A1(n4050), .A2(n_T_427[18]), .Y(n7490) );
  AO22X1_LVT U8796 ( .A1(n4026), .A2(n_T_427[913]), .A3(n4019), .A4(
        n_T_427[658]), .Y(n7489) );
  AO22X1_LVT U8797 ( .A1(n3977), .A2(n_T_427[530]), .A3(n4029), .A4(
        n_T_427[849]), .Y(n7488) );
  AO22X1_LVT U8798 ( .A1(n4033), .A2(n_T_427[594]), .A3(n3984), .A4(
        n_T_427[210]), .Y(n7487) );
  NOR4X1_LVT U8799 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .Y(n7496)
         );
  AO22X1_LVT U8800 ( .A1(n3969), .A2(n_T_427[402]), .A3(n3965), .A4(
        n_T_427[274]), .Y(n7494) );
  AO22X1_LVT U8801 ( .A1(n2858), .A2(n_T_427[146]), .A3(n4039), .A4(
        n_T_427[338]), .Y(n7493) );
  AO22X1_LVT U8802 ( .A1(n3981), .A2(n_T_427[785]), .A3(n4046), .A4(
        n_T_427[722]), .Y(n7492) );
  AO22X1_LVT U8803 ( .A1(n3962), .A2(n_T_427[466]), .A3(n2836), .A4(
        n_T_427[82]), .Y(n7491) );
  NOR4X1_LVT U8804 ( .A1(n7494), .A2(n7493), .A3(n7492), .A4(n7491), .Y(n7495)
         );
  AO21X1_LVT U8805 ( .A1(n7496), .A2(n7495), .A3(n2154), .Y(n7497) );
  NAND2X0_LVT U8806 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[18]), .Y(n7503) );
  NAND2X0_LVT U8807 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[18]), .Y(n7502)
         );
  NAND2X0_LVT U8808 ( .A1(n2497), .A2(n_T_628[18]), .Y(n7501) );
  NAND2X0_LVT U8809 ( .A1(n9066), .A2(n_T_918[18]), .Y(n7500) );
  NAND4X0_LVT U8810 ( .A1(n7503), .A2(n7502), .A3(n7501), .A4(n7500), .Y(
        io_fpu_fromint_data[18]) );
  NAND2X0_LVT U8811 ( .A1(n3997), .A2(n_T_427[1298]), .Y(n7504) );
  OA21X1_LVT U8812 ( .A1(n3446), .A2(n3751), .A3(n7504), .Y(n7507) );
  NAND2X0_LVT U8813 ( .A1(n3744), .A2(n_T_427[1682]), .Y(n7506) );
  NAND2X0_LVT U8814 ( .A1(n4002), .A2(n_T_427[1746]), .Y(n7505) );
  NAND2X0_LVT U8815 ( .A1(n3616), .A2(n_T_427[1554]), .Y(n7508) );
  OA21X1_LVT U8816 ( .A1(n4008), .A2(n3317), .A3(n7508), .Y(n7511) );
  NAND2X0_LVT U8817 ( .A1(n3648), .A2(n_T_427[1618]), .Y(n7510) );
  NAND2X0_LVT U8818 ( .A1(n4006), .A2(n_T_427[1490]), .Y(n7509) );
  NAND2X0_LVT U8819 ( .A1(n3712), .A2(n_T_427[978]), .Y(n7512) );
  OA21X1_LVT U8820 ( .A1(n3752), .A2(n3318), .A3(n7512), .Y(n7515) );
  NAND2X0_LVT U8821 ( .A1(n3640), .A2(n_T_427[1234]), .Y(n7514) );
  NAND2X0_LVT U8822 ( .A1(n3668), .A2(n_T_427[1106]), .Y(n7513) );
  NAND2X0_LVT U8823 ( .A1(n2882), .A2(n_T_427[1900]), .Y(n7516) );
  OA21X1_LVT U8824 ( .A1(n3987), .A2(n3319), .A3(n7516), .Y(n7519) );
  NAND2X0_LVT U8825 ( .A1(n3630), .A2(n_T_427[1426]), .Y(n7518) );
  NAND2X0_LVT U8826 ( .A1(n3608), .A2(n_T_427[1362]), .Y(n7517) );
  NAND2X0_LVT U8827 ( .A1(n3665), .A2(n4373), .Y(n7531) );
  AND2X1_LVT U8828 ( .A1(n4050), .A2(n_T_427[19]), .Y(n7523) );
  AO22X1_LVT U8829 ( .A1(n4025), .A2(n_T_427[914]), .A3(n4019), .A4(
        n_T_427[659]), .Y(n7522) );
  AO22X1_LVT U8830 ( .A1(n3978), .A2(n_T_427[531]), .A3(n4029), .A4(
        n_T_427[850]), .Y(n7521) );
  AO22X1_LVT U8831 ( .A1(n4033), .A2(n_T_427[595]), .A3(n3984), .A4(
        n_T_427[211]), .Y(n7520) );
  NOR4X1_LVT U8832 ( .A1(n7523), .A2(n7522), .A3(n7521), .A4(n7520), .Y(n7529)
         );
  AO22X1_LVT U8833 ( .A1(n3969), .A2(n_T_427[403]), .A3(n3965), .A4(
        n_T_427[275]), .Y(n7527) );
  AO22X1_LVT U8834 ( .A1(n3975), .A2(n_T_427[147]), .A3(n4038), .A4(
        n_T_427[339]), .Y(n7526) );
  AO22X1_LVT U8835 ( .A1(n3981), .A2(n_T_427[786]), .A3(n4046), .A4(
        n_T_427[723]), .Y(n7525) );
  AO22X1_LVT U8836 ( .A1(n3962), .A2(n_T_427[467]), .A3(n2837), .A4(
        n_T_427[83]), .Y(n7524) );
  NOR4X1_LVT U8837 ( .A1(n7527), .A2(n7526), .A3(n7525), .A4(n7524), .Y(n7528)
         );
  AO21X1_LVT U8838 ( .A1(n7529), .A2(n7528), .A3(n3632), .Y(n7530) );
  NAND2X0_LVT U8839 ( .A1(n3999), .A2(n_T_427[1299]), .Y(n7533) );
  OA21X1_LVT U8840 ( .A1(n3447), .A2(n3601), .A3(n7533), .Y(n7536) );
  NAND2X0_LVT U8841 ( .A1(n3744), .A2(n_T_427[1683]), .Y(n7535) );
  NAND2X0_LVT U8842 ( .A1(n4005), .A2(n_T_427[1747]), .Y(n7534) );
  NAND2X0_LVT U8843 ( .A1(n3617), .A2(n_T_427[1555]), .Y(n7537) );
  OA21X1_LVT U8844 ( .A1(n3663), .A2(n3320), .A3(n7537), .Y(n7540) );
  NAND2X0_LVT U8845 ( .A1(n3651), .A2(n_T_427[1619]), .Y(n7539) );
  NAND2X0_LVT U8846 ( .A1(n4007), .A2(n_T_427[1491]), .Y(n7538) );
  NAND2X0_LVT U8847 ( .A1(n3755), .A2(n_T_427[979]), .Y(n7541) );
  OA21X1_LVT U8848 ( .A1(n3752), .A2(n3321), .A3(n7541), .Y(n7544) );
  NAND2X0_LVT U8849 ( .A1(n3641), .A2(n_T_427[1235]), .Y(n7543) );
  NAND2X0_LVT U8850 ( .A1(n3670), .A2(n_T_427[1107]), .Y(n7542) );
  NAND2X0_LVT U8851 ( .A1(n3628), .A2(n_T_427[1427]), .Y(n7546) );
  NAND2X0_LVT U8852 ( .A1(n3604), .A2(n_T_427[1363]), .Y(n7545) );
  NAND2X0_LVT U8853 ( .A1(n2982), .A2(n4376), .Y(n7558) );
  AND2X1_LVT U8854 ( .A1(n4050), .A2(n_T_427[20]), .Y(n7550) );
  AO22X1_LVT U8855 ( .A1(n4025), .A2(n_T_427[915]), .A3(n4019), .A4(
        n_T_427[660]), .Y(n7549) );
  AO22X1_LVT U8856 ( .A1(n3978), .A2(n_T_427[532]), .A3(n4029), .A4(
        n_T_427[851]), .Y(n7548) );
  AO22X1_LVT U8857 ( .A1(n4033), .A2(n_T_427[596]), .A3(n3985), .A4(
        n_T_427[212]), .Y(n7547) );
  NOR4X1_LVT U8858 ( .A1(n7550), .A2(n7549), .A3(n7548), .A4(n7547), .Y(n7556)
         );
  AO22X1_LVT U8859 ( .A1(n3969), .A2(n_T_427[404]), .A3(n3965), .A4(
        n_T_427[276]), .Y(n7554) );
  AO22X1_LVT U8860 ( .A1(n2858), .A2(n_T_427[148]), .A3(n4038), .A4(
        n_T_427[340]), .Y(n7553) );
  AO22X1_LVT U8861 ( .A1(n3981), .A2(n_T_427[787]), .A3(n4046), .A4(
        n_T_427[724]), .Y(n7552) );
  AO22X1_LVT U8862 ( .A1(n3962), .A2(n_T_427[468]), .A3(n2836), .A4(
        n_T_427[84]), .Y(n7551) );
  NOR4X1_LVT U8863 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .Y(n7555)
         );
  AO21X1_LVT U8864 ( .A1(n7556), .A2(n7555), .A3(n3632), .Y(n7557) );
  NAND2X0_LVT U8865 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[20]), .Y(n7563) );
  NAND2X0_LVT U8866 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[20]), .Y(n7562)
         );
  NAND2X0_LVT U8867 ( .A1(n2497), .A2(n_T_628[20]), .Y(n7561) );
  NAND2X0_LVT U8868 ( .A1(n9066), .A2(n_T_918[20]), .Y(n7560) );
  NAND4X0_LVT U8869 ( .A1(n7563), .A2(n7562), .A3(n7561), .A4(n7560), .Y(
        io_fpu_fromint_data[20]) );
  NAND2X0_LVT U8870 ( .A1(n3996), .A2(n_T_427[1300]), .Y(n7564) );
  OA21X1_LVT U8871 ( .A1(n3391), .A2(n3601), .A3(n7564), .Y(n7567) );
  NAND2X0_LVT U8872 ( .A1(n3744), .A2(n_T_427[1684]), .Y(n7566) );
  NAND2X0_LVT U8873 ( .A1(n2091), .A2(n_T_427[1748]), .Y(n7565) );
  NAND2X0_LVT U8874 ( .A1(n3618), .A2(n_T_427[1556]), .Y(n7568) );
  OA21X1_LVT U8875 ( .A1(n3664), .A2(n3284), .A3(n7568), .Y(n7571) );
  NAND2X0_LVT U8876 ( .A1(n3648), .A2(n_T_427[1620]), .Y(n7570) );
  NAND2X0_LVT U8877 ( .A1(n4006), .A2(n_T_427[1492]), .Y(n7569) );
  NAND2X0_LVT U8878 ( .A1(n3758), .A2(n_T_427[980]), .Y(n7572) );
  OA21X1_LVT U8879 ( .A1(n3752), .A2(n3285), .A3(n7572), .Y(n7575) );
  NAND2X0_LVT U8880 ( .A1(n3639), .A2(n_T_427[1236]), .Y(n7574) );
  NAND2X0_LVT U8881 ( .A1(n3671), .A2(n_T_427[1108]), .Y(n7573) );
  NAND2X0_LVT U8882 ( .A1(n3992), .A2(n_T_427[1902]), .Y(n7576) );
  NAND2X0_LVT U8883 ( .A1(n3630), .A2(n_T_427[1428]), .Y(n7578) );
  NAND2X0_LVT U8884 ( .A1(n3602), .A2(n_T_427[1364]), .Y(n7577) );
  NAND2X0_LVT U8885 ( .A1(n3060), .A2(n4378), .Y(n7590) );
  AND2X1_LVT U8886 ( .A1(n4050), .A2(n_T_427[21]), .Y(n7582) );
  AO22X1_LVT U8887 ( .A1(n4025), .A2(n_T_427[916]), .A3(n4019), .A4(
        n_T_427[661]), .Y(n7581) );
  AO22X1_LVT U8888 ( .A1(n3978), .A2(n_T_427[533]), .A3(n4029), .A4(
        n_T_427[852]), .Y(n7580) );
  AO22X1_LVT U8889 ( .A1(n4033), .A2(n_T_427[597]), .A3(n3985), .A4(
        n_T_427[213]), .Y(n7579) );
  NOR4X1_LVT U8890 ( .A1(n7582), .A2(n7581), .A3(n7580), .A4(n7579), .Y(n7588)
         );
  AO22X1_LVT U8891 ( .A1(n3969), .A2(n_T_427[405]), .A3(n3965), .A4(
        n_T_427[277]), .Y(n7586) );
  AO22X1_LVT U8892 ( .A1(n2859), .A2(n_T_427[149]), .A3(n4038), .A4(
        n_T_427[341]), .Y(n7585) );
  AO22X1_LVT U8893 ( .A1(n3981), .A2(n_T_427[788]), .A3(n4046), .A4(
        n_T_427[725]), .Y(n7584) );
  AO22X1_LVT U8894 ( .A1(n3962), .A2(n_T_427[469]), .A3(n4041), .A4(
        n_T_427[85]), .Y(n7583) );
  NOR4X1_LVT U8895 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .Y(n7587)
         );
  NAND2X0_LVT U8896 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[21]), .Y(n7595) );
  NAND2X0_LVT U8897 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[21]), .Y(n7594)
         );
  NAND2X0_LVT U8898 ( .A1(n2497), .A2(n_T_628[21]), .Y(n7593) );
  NAND2X0_LVT U8899 ( .A1(n9066), .A2(n_T_918[21]), .Y(n7592) );
  NAND4X0_LVT U8900 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .Y(
        io_fpu_fromint_data[21]) );
  NAND2X0_LVT U8901 ( .A1(n2094), .A2(n_T_427[1301]), .Y(n7596) );
  OA21X1_LVT U8902 ( .A1(n3392), .A2(n3601), .A3(n7596), .Y(n7599) );
  NAND2X0_LVT U8903 ( .A1(n3744), .A2(n_T_427[1685]), .Y(n7598) );
  NAND2X0_LVT U8904 ( .A1(n4004), .A2(n_T_427[1749]), .Y(n7597) );
  NAND2X0_LVT U8905 ( .A1(n3619), .A2(n_T_427[1557]), .Y(n7600) );
  OA21X1_LVT U8906 ( .A1(n4010), .A2(n3286), .A3(n7600), .Y(n7603) );
  NAND2X0_LVT U8907 ( .A1(n3649), .A2(n_T_427[1621]), .Y(n7602) );
  NAND2X0_LVT U8908 ( .A1(n4006), .A2(n_T_427[1493]), .Y(n7601) );
  NAND2X0_LVT U8909 ( .A1(n3755), .A2(n_T_427[981]), .Y(n7604) );
  OA21X1_LVT U8910 ( .A1(n3752), .A2(n3287), .A3(n7604), .Y(n7607) );
  NAND2X0_LVT U8911 ( .A1(n_T_427[1237]), .A2(n3638), .Y(n7606) );
  NAND2X0_LVT U8912 ( .A1(n3670), .A2(n_T_427[1109]), .Y(n7605) );
  NAND2X0_LVT U8913 ( .A1(n2967), .A2(n_T_427[1429]), .Y(n7609) );
  NAND2X0_LVT U8914 ( .A1(n3609), .A2(n_T_427[1365]), .Y(n7608) );
  NAND2X0_LVT U8915 ( .A1(n3060), .A2(n4380), .Y(n7621) );
  AND2X1_LVT U8916 ( .A1(n4050), .A2(n_T_427[22]), .Y(n7613) );
  AO22X1_LVT U8917 ( .A1(n4025), .A2(n_T_427[917]), .A3(n4019), .A4(
        n_T_427[662]), .Y(n7612) );
  AO22X1_LVT U8918 ( .A1(n3978), .A2(n_T_427[534]), .A3(n4028), .A4(
        n_T_427[853]), .Y(n7611) );
  AO22X1_LVT U8919 ( .A1(n4033), .A2(n_T_427[598]), .A3(n3985), .A4(
        n_T_427[214]), .Y(n7610) );
  NOR4X1_LVT U8920 ( .A1(n7613), .A2(n7612), .A3(n7611), .A4(n7610), .Y(n7619)
         );
  AO22X1_LVT U8921 ( .A1(n3969), .A2(n_T_427[406]), .A3(n3965), .A4(
        n_T_427[278]), .Y(n7617) );
  AO22X1_LVT U8922 ( .A1(n2859), .A2(n_T_427[150]), .A3(n4038), .A4(
        n_T_427[342]), .Y(n7616) );
  AO22X1_LVT U8923 ( .A1(n3981), .A2(n_T_427[789]), .A3(n4046), .A4(
        n_T_427[726]), .Y(n7615) );
  AO22X1_LVT U8924 ( .A1(n3962), .A2(n_T_427[470]), .A3(n2837), .A4(
        n_T_427[86]), .Y(n7614) );
  NOR4X1_LVT U8925 ( .A1(n7617), .A2(n7616), .A3(n7615), .A4(n7614), .Y(n7618)
         );
  AO21X1_LVT U8926 ( .A1(n7619), .A2(n7618), .A3(n2155), .Y(n7620) );
  NAND2X0_LVT U8927 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[22]), .Y(n7626) );
  NAND2X0_LVT U8928 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[22]), .Y(n7625)
         );
  NAND2X0_LVT U8929 ( .A1(n2497), .A2(n_T_628[22]), .Y(n7624) );
  NAND2X0_LVT U8930 ( .A1(n9066), .A2(n_T_918[22]), .Y(n7623) );
  NAND4X0_LVT U8931 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .Y(
        io_fpu_fromint_data[22]) );
  NAND2X0_LVT U8932 ( .A1(n2094), .A2(n_T_427[1302]), .Y(n7627) );
  OA21X1_LVT U8933 ( .A1(n3448), .A2(n3751), .A3(n7627), .Y(n7630) );
  NAND2X0_LVT U8934 ( .A1(n3657), .A2(n_T_427[1686]), .Y(n7629) );
  NAND2X0_LVT U8935 ( .A1(n2092), .A2(n_T_427[1750]), .Y(n7628) );
  NAND2X0_LVT U8936 ( .A1(n3621), .A2(n_T_427[1558]), .Y(n7631) );
  OA21X1_LVT U8937 ( .A1(n2081), .A2(n3323), .A3(n7631), .Y(n7634) );
  NAND2X0_LVT U8938 ( .A1(n3642), .A2(n_T_427[1622]), .Y(n7633) );
  NAND2X0_LVT U8939 ( .A1(n4006), .A2(n_T_427[1494]), .Y(n7632) );
  NAND2X0_LVT U8940 ( .A1(n3760), .A2(n_T_427[982]), .Y(n7635) );
  OA21X1_LVT U8941 ( .A1(n3752), .A2(n3324), .A3(n7635), .Y(n7638) );
  NAND2X0_LVT U8942 ( .A1(n_T_427[1238]), .A2(n3638), .Y(n7637) );
  NAND2X0_LVT U8943 ( .A1(n3672), .A2(n_T_427[1110]), .Y(n7636) );
  NAND2X0_LVT U8944 ( .A1(n3991), .A2(n_T_427[1904]), .Y(n7639) );
  OA21X1_LVT U8945 ( .A1(n3989), .A2(n3325), .A3(n7639), .Y(n7642) );
  NAND2X0_LVT U8946 ( .A1(n3626), .A2(n_T_427[1430]), .Y(n7641) );
  NAND2X0_LVT U8947 ( .A1(n3602), .A2(n_T_427[1366]), .Y(n7640) );
  NAND2X0_LVT U8948 ( .A1(n4015), .A2(n4383), .Y(n7654) );
  AND2X1_LVT U8949 ( .A1(n4050), .A2(n_T_427[23]), .Y(n7646) );
  AO22X1_LVT U8950 ( .A1(n4025), .A2(n_T_427[918]), .A3(n4020), .A4(
        n_T_427[663]), .Y(n7645) );
  AO22X1_LVT U8951 ( .A1(n3978), .A2(n_T_427[535]), .A3(n4028), .A4(
        n_T_427[854]), .Y(n7644) );
  AO22X1_LVT U8952 ( .A1(n4033), .A2(n_T_427[599]), .A3(n3985), .A4(
        n_T_427[215]), .Y(n7643) );
  NOR4X1_LVT U8953 ( .A1(n7646), .A2(n7645), .A3(n7644), .A4(n7643), .Y(n7652)
         );
  AO22X1_LVT U8954 ( .A1(n3969), .A2(n_T_427[407]), .A3(n3965), .A4(
        n_T_427[279]), .Y(n7650) );
  AO22X1_LVT U8955 ( .A1(n3973), .A2(n_T_427[151]), .A3(n4038), .A4(
        n_T_427[343]), .Y(n7649) );
  AO22X1_LVT U8956 ( .A1(n3981), .A2(n_T_427[790]), .A3(n4046), .A4(
        n_T_427[727]), .Y(n7648) );
  AO22X1_LVT U8957 ( .A1(n3962), .A2(n_T_427[471]), .A3(n2837), .A4(
        n_T_427[87]), .Y(n7647) );
  NOR4X1_LVT U8958 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .Y(n7651)
         );
  AO21X1_LVT U8959 ( .A1(n7652), .A2(n7651), .A3(n2155), .Y(n7653) );
  NAND2X0_LVT U8960 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[23]), .Y(n7659) );
  NAND2X0_LVT U8961 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[23]), .Y(n7658)
         );
  NAND2X0_LVT U8962 ( .A1(n2497), .A2(n_T_628[23]), .Y(n7657) );
  NAND2X0_LVT U8963 ( .A1(n9066), .A2(n_T_918[23]), .Y(n7656) );
  NAND4X0_LVT U8964 ( .A1(n7659), .A2(n7658), .A3(n7657), .A4(n7656), .Y(
        io_fpu_fromint_data[23]) );
  NAND2X0_LVT U8965 ( .A1(n4000), .A2(n_T_427[1303]), .Y(n7660) );
  OA21X1_LVT U8966 ( .A1(n3449), .A2(n3747), .A3(n7660), .Y(n7663) );
  NAND2X0_LVT U8967 ( .A1(n2922), .A2(n_T_427[1687]), .Y(n7662) );
  NAND2X0_LVT U8968 ( .A1(n2091), .A2(n_T_427[1751]), .Y(n7661) );
  NAND3X0_LVT U8969 ( .A1(n7663), .A2(n7662), .A3(n7661), .Y(n7685) );
  NAND2X0_LVT U8970 ( .A1(n3620), .A2(n_T_427[1559]), .Y(n7664) );
  OA21X1_LVT U8971 ( .A1(n4010), .A2(n3326), .A3(n7664), .Y(n7667) );
  NAND2X0_LVT U8972 ( .A1(n3651), .A2(n_T_427[1623]), .Y(n7666) );
  NAND2X0_LVT U8973 ( .A1(n4006), .A2(n_T_427[1495]), .Y(n7665) );
  NAND3X0_LVT U8974 ( .A1(n7667), .A2(n7666), .A3(n7665), .Y(n7684) );
  NAND2X0_LVT U8975 ( .A1(n3759), .A2(n_T_427[983]), .Y(n7668) );
  NAND2X0_LVT U8976 ( .A1(n3640), .A2(n_T_427[1239]), .Y(n7670) );
  NAND2X0_LVT U8977 ( .A1(n3672), .A2(n_T_427[1111]), .Y(n7669) );
  NAND2X0_LVT U8978 ( .A1(n2882), .A2(n_T_427[1905]), .Y(n7671) );
  NAND2X0_LVT U8979 ( .A1(n3604), .A2(n_T_427[1367]), .Y(n7672) );
  NAND2X0_LVT U8980 ( .A1(n3665), .A2(n4386), .Y(n7682) );
  AND2X1_LVT U8981 ( .A1(n4050), .A2(n_T_427[24]), .Y(n7676) );
  AO22X1_LVT U8982 ( .A1(n4025), .A2(n_T_427[919]), .A3(n4020), .A4(
        n_T_427[664]), .Y(n7675) );
  AO22X1_LVT U8983 ( .A1(n3978), .A2(n_T_427[536]), .A3(n4028), .A4(
        n_T_427[855]), .Y(n7674) );
  AO22X1_LVT U8984 ( .A1(n4033), .A2(n_T_427[600]), .A3(n3985), .A4(
        n_T_427[216]), .Y(n7673) );
  AO22X1_LVT U8985 ( .A1(n3969), .A2(n_T_427[408]), .A3(n3966), .A4(
        n_T_427[280]), .Y(n7680) );
  AO22X1_LVT U8986 ( .A1(n3973), .A2(n_T_427[152]), .A3(n4038), .A4(
        n_T_427[344]), .Y(n7679) );
  AO22X1_LVT U8987 ( .A1(n3981), .A2(n_T_427[791]), .A3(n4047), .A4(
        n_T_427[728]), .Y(n7678) );
  AO22X1_LVT U8988 ( .A1(n3962), .A2(n_T_427[472]), .A3(n4042), .A4(
        n_T_427[88]), .Y(n7677) );
  NAND2X0_LVT U8989 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[24]), .Y(n7689) );
  NAND2X0_LVT U8990 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[24]), .Y(n7688)
         );
  NAND2X0_LVT U8991 ( .A1(n2497), .A2(n_T_628[24]), .Y(n7687) );
  NAND2X0_LVT U8992 ( .A1(n9066), .A2(n_T_918[24]), .Y(n7686) );
  NAND4X0_LVT U8993 ( .A1(n7689), .A2(n7688), .A3(n7687), .A4(n7686), .Y(
        io_fpu_fromint_data[24]) );
  NAND2X0_LVT U8994 ( .A1(n3999), .A2(n_T_427[1304]), .Y(n7690) );
  OA21X1_LVT U8995 ( .A1(n3393), .A2(n3747), .A3(n7690), .Y(n7693) );
  NAND2X0_LVT U8996 ( .A1(n3744), .A2(n_T_427[1688]), .Y(n7692) );
  NAND2X0_LVT U8997 ( .A1(n2091), .A2(n_T_427[1752]), .Y(n7691) );
  NAND2X0_LVT U8998 ( .A1(n3621), .A2(n_T_427[1560]), .Y(n7694) );
  OA21X1_LVT U8999 ( .A1(n4009), .A2(n3288), .A3(n7694), .Y(n7697) );
  NAND2X0_LVT U9000 ( .A1(n3643), .A2(n_T_427[1624]), .Y(n7696) );
  NAND2X0_LVT U9001 ( .A1(n4007), .A2(n_T_427[1496]), .Y(n7695) );
  NAND2X0_LVT U9002 ( .A1(n3758), .A2(n_T_427[984]), .Y(n7698) );
  OA21X1_LVT U9003 ( .A1(n3752), .A2(n3289), .A3(n7698), .Y(n7701) );
  NAND2X0_LVT U9004 ( .A1(n3636), .A2(n_T_427[1240]), .Y(n7700) );
  NAND2X0_LVT U9005 ( .A1(n3674), .A2(n_T_427[1112]), .Y(n7699) );
  NAND2X0_LVT U9006 ( .A1(n2998), .A2(n_T_427[1906]), .Y(n7702) );
  OA21X1_LVT U9007 ( .A1(n3989), .A2(n3372), .A3(n7702), .Y(n7705) );
  NAND2X0_LVT U9008 ( .A1(n3626), .A2(n_T_427[1432]), .Y(n7704) );
  NAND2X0_LVT U9009 ( .A1(n3603), .A2(n_T_427[1368]), .Y(n7703) );
  NAND2X0_LVT U9010 ( .A1(n3060), .A2(n4388), .Y(n7717) );
  AND2X1_LVT U9011 ( .A1(n4051), .A2(n_T_427[25]), .Y(n7709) );
  AO22X1_LVT U9012 ( .A1(n4025), .A2(n_T_427[920]), .A3(n4020), .A4(
        n_T_427[665]), .Y(n7708) );
  AO22X1_LVT U9013 ( .A1(n3976), .A2(n_T_427[537]), .A3(n4028), .A4(
        n_T_427[856]), .Y(n7707) );
  AO22X1_LVT U9014 ( .A1(n4033), .A2(n_T_427[601]), .A3(n3985), .A4(
        n_T_427[217]), .Y(n7706) );
  NOR4X1_LVT U9015 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .Y(n7715)
         );
  AO22X1_LVT U9016 ( .A1(n3970), .A2(n_T_427[409]), .A3(n3966), .A4(
        n_T_427[281]), .Y(n7713) );
  AO22X1_LVT U9017 ( .A1(n2858), .A2(n_T_427[153]), .A3(n4038), .A4(
        n_T_427[345]), .Y(n7712) );
  AO22X1_LVT U9018 ( .A1(n3981), .A2(n_T_427[792]), .A3(n4047), .A4(
        n_T_427[729]), .Y(n7711) );
  AO22X1_LVT U9019 ( .A1(n3962), .A2(n_T_427[473]), .A3(n4044), .A4(
        n_T_427[89]), .Y(n7710) );
  NOR4X1_LVT U9020 ( .A1(n7713), .A2(n7712), .A3(n7711), .A4(n7710), .Y(n7714)
         );
  AO21X1_LVT U9021 ( .A1(n7715), .A2(n7714), .A3(n2645), .Y(n7716) );
  NAND2X0_LVT U9022 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[25]), .Y(n7722) );
  NAND2X0_LVT U9023 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[25]), .Y(n7721)
         );
  NAND2X0_LVT U9024 ( .A1(n2497), .A2(n_T_628[25]), .Y(n7720) );
  NAND2X0_LVT U9025 ( .A1(n9066), .A2(n_T_918[25]), .Y(n7719) );
  NAND4X0_LVT U9026 ( .A1(n7722), .A2(n7721), .A3(n7720), .A4(n7719), .Y(
        io_fpu_fromint_data[25]) );
  NAND2X0_LVT U9027 ( .A1(n3997), .A2(n_T_427[1305]), .Y(n7723) );
  OA21X1_LVT U9028 ( .A1(n3394), .A2(n3747), .A3(n7723), .Y(n7726) );
  NAND2X0_LVT U9029 ( .A1(n3744), .A2(n_T_427[1689]), .Y(n7725) );
  NAND2X0_LVT U9030 ( .A1(n4001), .A2(n_T_427[1753]), .Y(n7724) );
  NAND2X0_LVT U9031 ( .A1(n3621), .A2(n_T_427[1561]), .Y(n7727) );
  OA21X1_LVT U9032 ( .A1(n2081), .A2(n3290), .A3(n7727), .Y(n7730) );
  NAND2X0_LVT U9033 ( .A1(n3652), .A2(n_T_427[1625]), .Y(n7729) );
  NAND2X0_LVT U9034 ( .A1(n4006), .A2(n_T_427[1497]), .Y(n7728) );
  NAND2X0_LVT U9035 ( .A1(n3756), .A2(n_T_427[985]), .Y(n7731) );
  OA21X1_LVT U9036 ( .A1(n3752), .A2(n3291), .A3(n7731), .Y(n7734) );
  NAND2X0_LVT U9037 ( .A1(n3637), .A2(n_T_427[1241]), .Y(n7733) );
  NAND2X0_LVT U9038 ( .A1(n3675), .A2(n_T_427[1113]), .Y(n7732) );
  NAND2X0_LVT U9039 ( .A1(n2998), .A2(n_T_427[1907]), .Y(n7735) );
  OA21X1_LVT U9040 ( .A1(n3987), .A2(n3373), .A3(n7735), .Y(n7738) );
  NAND2X0_LVT U9041 ( .A1(n3628), .A2(n_T_427[1433]), .Y(n7737) );
  NAND2X0_LVT U9042 ( .A1(n3603), .A2(n_T_427[1369]), .Y(n7736) );
  NAND2X0_LVT U9043 ( .A1(n2982), .A2(n4390), .Y(n7750) );
  AND2X1_LVT U9044 ( .A1(n4051), .A2(n_T_427[26]), .Y(n7742) );
  AO22X1_LVT U9045 ( .A1(n4025), .A2(n_T_427[921]), .A3(n4020), .A4(
        n_T_427[666]), .Y(n7741) );
  AO22X1_LVT U9046 ( .A1(n3978), .A2(n_T_427[538]), .A3(n4028), .A4(
        n_T_427[857]), .Y(n7740) );
  AO22X1_LVT U9047 ( .A1(n4033), .A2(n_T_427[602]), .A3(n3985), .A4(
        n_T_427[218]), .Y(n7739) );
  NOR4X1_LVT U9048 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .Y(n7748)
         );
  AO22X1_LVT U9049 ( .A1(n3970), .A2(n_T_427[410]), .A3(n3966), .A4(
        n_T_427[282]), .Y(n7746) );
  AO22X1_LVT U9050 ( .A1(n3975), .A2(n_T_427[154]), .A3(n4038), .A4(
        n_T_427[346]), .Y(n7745) );
  AO22X1_LVT U9051 ( .A1(n3981), .A2(n_T_427[793]), .A3(n4047), .A4(
        n_T_427[730]), .Y(n7744) );
  AO22X1_LVT U9052 ( .A1(n3962), .A2(n_T_427[474]), .A3(n4041), .A4(
        n_T_427[90]), .Y(n7743) );
  NOR4X1_LVT U9053 ( .A1(n7746), .A2(n7745), .A3(n7744), .A4(n7743), .Y(n7747)
         );
  NAND2X0_LVT U9054 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[26]), .Y(n7755) );
  NAND2X0_LVT U9055 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[26]), .Y(n7754)
         );
  NAND2X0_LVT U9056 ( .A1(n2497), .A2(n_T_628[26]), .Y(n7753) );
  NAND2X0_LVT U9057 ( .A1(n9066), .A2(n_T_918[26]), .Y(n7752) );
  NAND4X0_LVT U9058 ( .A1(n7755), .A2(n7754), .A3(n7753), .A4(n7752), .Y(
        io_fpu_fromint_data[26]) );
  NAND2X0_LVT U9059 ( .A1(n3999), .A2(n_T_427[1306]), .Y(n7756) );
  OA21X1_LVT U9060 ( .A1(n3450), .A2(n3751), .A3(n7756), .Y(n7759) );
  NAND2X0_LVT U9061 ( .A1(n3744), .A2(n_T_427[1690]), .Y(n7758) );
  NAND2X0_LVT U9062 ( .A1(n4002), .A2(n_T_427[1754]), .Y(n7757) );
  NAND2X0_LVT U9063 ( .A1(n3618), .A2(n_T_427[1562]), .Y(n7760) );
  OA21X1_LVT U9064 ( .A1(n2081), .A2(n3328), .A3(n7760), .Y(n7762) );
  NAND2X0_LVT U9065 ( .A1(n4007), .A2(n_T_427[1498]), .Y(n7761) );
  NAND2X0_LVT U9066 ( .A1(n3757), .A2(n_T_427[986]), .Y(n7763) );
  OA21X1_LVT U9067 ( .A1(n3752), .A2(n3329), .A3(n7763), .Y(n7766) );
  NAND2X0_LVT U9068 ( .A1(n3636), .A2(n_T_427[1242]), .Y(n7765) );
  NAND2X0_LVT U9069 ( .A1(n3672), .A2(n_T_427[1114]), .Y(n7764) );
  NAND2X0_LVT U9070 ( .A1(n2985), .A2(n_T_427[1908]), .Y(n7767) );
  OA21X1_LVT U9071 ( .A1(n2120), .A2(n3330), .A3(n7767), .Y(n7770) );
  NAND2X0_LVT U9072 ( .A1(n2966), .A2(n_T_427[1434]), .Y(n7769) );
  NAND2X0_LVT U9073 ( .A1(n3607), .A2(n_T_427[1370]), .Y(n7768) );
  NAND2X0_LVT U9074 ( .A1(n4015), .A2(n4393), .Y(n7782) );
  AND2X1_LVT U9075 ( .A1(n4051), .A2(n_T_427[27]), .Y(n7774) );
  AO22X1_LVT U9076 ( .A1(n4025), .A2(n_T_427[922]), .A3(n4020), .A4(
        n_T_427[667]), .Y(n7773) );
  AO22X1_LVT U9077 ( .A1(n3978), .A2(n_T_427[539]), .A3(n4028), .A4(
        n_T_427[858]), .Y(n7772) );
  AO22X1_LVT U9078 ( .A1(n4033), .A2(n_T_427[603]), .A3(n3985), .A4(
        n_T_427[219]), .Y(n7771) );
  NOR4X1_LVT U9079 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .Y(n7780)
         );
  AO22X1_LVT U9080 ( .A1(n3970), .A2(n_T_427[411]), .A3(n3966), .A4(
        n_T_427[283]), .Y(n7778) );
  AO22X1_LVT U9081 ( .A1(n3973), .A2(n_T_427[155]), .A3(n4038), .A4(
        n_T_427[347]), .Y(n7777) );
  AO22X1_LVT U9082 ( .A1(n3981), .A2(n_T_427[794]), .A3(n4047), .A4(
        n_T_427[731]), .Y(n7776) );
  AO22X1_LVT U9083 ( .A1(n3962), .A2(n_T_427[475]), .A3(n2836), .A4(
        n_T_427[91]), .Y(n7775) );
  NOR4X1_LVT U9084 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .Y(n7779)
         );
  NAND2X0_LVT U9085 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[27]), .Y(n7787) );
  NAND2X0_LVT U9086 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[27]), .Y(n7786)
         );
  NAND2X0_LVT U9087 ( .A1(n2497), .A2(n_T_628[27]), .Y(n7785) );
  NAND2X0_LVT U9088 ( .A1(n9066), .A2(n_T_918[27]), .Y(n7784) );
  NAND4X0_LVT U9089 ( .A1(n7787), .A2(n7786), .A3(n7785), .A4(n7784), .Y(
        io_fpu_fromint_data[27]) );
  NAND2X0_LVT U9090 ( .A1(n2093), .A2(n_T_427[1307]), .Y(n7788) );
  OA21X1_LVT U9091 ( .A1(n3395), .A2(n3601), .A3(n7788), .Y(n7791) );
  NAND2X0_LVT U9092 ( .A1(n3744), .A2(n_T_427[1691]), .Y(n7790) );
  NAND2X0_LVT U9093 ( .A1(n4004), .A2(n_T_427[1755]), .Y(n7789) );
  NAND2X0_LVT U9094 ( .A1(n3615), .A2(n_T_427[1563]), .Y(n7792) );
  OA21X1_LVT U9095 ( .A1(n4008), .A2(n3292), .A3(n7792), .Y(n7794) );
  NAND2X0_LVT U9096 ( .A1(n4007), .A2(n_T_427[1499]), .Y(n7793) );
  NAND2X0_LVT U9097 ( .A1(n3760), .A2(n_T_427[987]), .Y(n7795) );
  OA21X1_LVT U9098 ( .A1(n4012), .A2(n3293), .A3(n7795), .Y(n7798) );
  NAND2X0_LVT U9099 ( .A1(n3639), .A2(n_T_427[1243]), .Y(n7797) );
  NAND2X0_LVT U9100 ( .A1(n3672), .A2(n_T_427[1115]), .Y(n7796) );
  NAND2X0_LVT U9101 ( .A1(n3992), .A2(n_T_427[1909]), .Y(n7799) );
  OA21X1_LVT U9102 ( .A1(n3767), .A2(n3374), .A3(n7799), .Y(n7802) );
  NAND2X0_LVT U9103 ( .A1(n3630), .A2(n_T_427[1435]), .Y(n7801) );
  NAND2X0_LVT U9104 ( .A1(n3604), .A2(n_T_427[1371]), .Y(n7800) );
  AND2X1_LVT U9105 ( .A1(n4051), .A2(n_T_427[28]), .Y(n7806) );
  AO22X1_LVT U9106 ( .A1(n4025), .A2(n_T_427[923]), .A3(n4020), .A4(
        n_T_427[668]), .Y(n7805) );
  AO22X1_LVT U9107 ( .A1(n3978), .A2(n_T_427[540]), .A3(n4028), .A4(
        n_T_427[859]), .Y(n7804) );
  AO22X1_LVT U9108 ( .A1(n4033), .A2(n_T_427[604]), .A3(n3985), .A4(
        n_T_427[220]), .Y(n7803) );
  NOR4X1_LVT U9109 ( .A1(n7806), .A2(n7805), .A3(n7804), .A4(n7803), .Y(n7812)
         );
  AO22X1_LVT U9110 ( .A1(n3970), .A2(n_T_427[412]), .A3(n3966), .A4(
        n_T_427[284]), .Y(n7810) );
  AO22X1_LVT U9111 ( .A1(n3974), .A2(n_T_427[156]), .A3(n4038), .A4(
        n_T_427[348]), .Y(n7809) );
  AO22X1_LVT U9112 ( .A1(n3981), .A2(n_T_427[795]), .A3(n4047), .A4(
        n_T_427[732]), .Y(n7808) );
  AO22X1_LVT U9113 ( .A1(n3962), .A2(n_T_427[476]), .A3(n4043), .A4(
        n_T_427[92]), .Y(n7807) );
  NOR4X1_LVT U9114 ( .A1(n7810), .A2(n7809), .A3(n7808), .A4(n7807), .Y(n7811)
         );
  NAND2X0_LVT U9115 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[28]), .Y(n7819) );
  NAND2X0_LVT U9116 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[28]), .Y(n7818)
         );
  NAND2X0_LVT U9117 ( .A1(n2493), .A2(n_T_628[28]), .Y(n7817) );
  NAND2X0_LVT U9118 ( .A1(n9066), .A2(n_T_918[28]), .Y(n7816) );
  NAND4X0_LVT U9119 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .Y(
        io_fpu_fromint_data[28]) );
  NAND2X0_LVT U9120 ( .A1(n4000), .A2(n_T_427[1308]), .Y(n7820) );
  OA21X1_LVT U9121 ( .A1(n3396), .A2(n3601), .A3(n7820), .Y(n7823) );
  NAND2X0_LVT U9122 ( .A1(n3744), .A2(n_T_427[1692]), .Y(n7822) );
  NAND2X0_LVT U9123 ( .A1(n4003), .A2(n_T_427[1756]), .Y(n7821) );
  NAND2X0_LVT U9124 ( .A1(n3616), .A2(n_T_427[1564]), .Y(n7824) );
  OA21X1_LVT U9125 ( .A1(n4008), .A2(n3294), .A3(n7824), .Y(n7827) );
  NAND2X0_LVT U9126 ( .A1(n3642), .A2(n_T_427[1628]), .Y(n7826) );
  NAND2X0_LVT U9127 ( .A1(n4007), .A2(n_T_427[1500]), .Y(n7825) );
  NAND2X0_LVT U9128 ( .A1(n3755), .A2(n_T_427[988]), .Y(n7828) );
  OA21X1_LVT U9129 ( .A1(n4013), .A2(n3295), .A3(n7828), .Y(n7831) );
  NAND2X0_LVT U9130 ( .A1(n3640), .A2(n_T_427[1244]), .Y(n7830) );
  NAND2X0_LVT U9131 ( .A1(n3675), .A2(n_T_427[1116]), .Y(n7829) );
  NAND2X0_LVT U9132 ( .A1(n2986), .A2(n_T_427[1910]), .Y(n7832) );
  OA21X1_LVT U9133 ( .A1(n2120), .A2(n3375), .A3(n7832), .Y(n7835) );
  NAND2X0_LVT U9134 ( .A1(n2967), .A2(n_T_427[1436]), .Y(n7834) );
  NAND2X0_LVT U9135 ( .A1(n3603), .A2(n_T_427[1372]), .Y(n7833) );
  AND2X1_LVT U9136 ( .A1(n4051), .A2(n_T_427[29]), .Y(n7839) );
  AO22X1_LVT U9137 ( .A1(n4025), .A2(n_T_427[924]), .A3(n4020), .A4(
        n_T_427[669]), .Y(n7838) );
  AO22X1_LVT U9138 ( .A1(n3978), .A2(n_T_427[541]), .A3(n4028), .A4(
        n_T_427[860]), .Y(n7837) );
  AO22X1_LVT U9139 ( .A1(n4034), .A2(n_T_427[605]), .A3(n3985), .A4(
        n_T_427[221]), .Y(n7836) );
  NOR4X1_LVT U9140 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .Y(n7845)
         );
  AO22X1_LVT U9141 ( .A1(n3970), .A2(n_T_427[413]), .A3(n3966), .A4(
        n_T_427[285]), .Y(n7843) );
  AO22X1_LVT U9142 ( .A1(n3974), .A2(n_T_427[157]), .A3(n4038), .A4(
        n_T_427[349]), .Y(n7842) );
  AO22X1_LVT U9143 ( .A1(n3981), .A2(n_T_427[796]), .A3(n4047), .A4(
        n_T_427[733]), .Y(n7841) );
  AO22X1_LVT U9144 ( .A1(n3962), .A2(n_T_427[477]), .A3(n4041), .A4(
        n_T_427[93]), .Y(n7840) );
  NOR4X1_LVT U9145 ( .A1(n7843), .A2(n7842), .A3(n7841), .A4(n7840), .Y(n7844)
         );
  AO21X1_LVT U9146 ( .A1(n7845), .A2(n7844), .A3(n3656), .Y(n7846) );
  NAND2X0_LVT U9147 ( .A1(n3998), .A2(n_T_427[1309]), .Y(n7849) );
  OA21X1_LVT U9148 ( .A1(n3451), .A2(n3601), .A3(n7849), .Y(n7852) );
  NAND2X0_LVT U9149 ( .A1(n3744), .A2(n_T_427[1693]), .Y(n7851) );
  NAND2X0_LVT U9150 ( .A1(n2091), .A2(n_T_427[1757]), .Y(n7850) );
  NAND2X0_LVT U9151 ( .A1(n3617), .A2(n_T_427[1565]), .Y(n7853) );
  OA21X1_LVT U9152 ( .A1(n4010), .A2(n3331), .A3(n7853), .Y(n7856) );
  NAND2X0_LVT U9153 ( .A1(n3651), .A2(n_T_427[1629]), .Y(n7855) );
  NAND2X0_LVT U9154 ( .A1(n3769), .A2(n_T_427[1501]), .Y(n7854) );
  NAND2X0_LVT U9155 ( .A1(n_T_427[1245]), .A2(n3638), .Y(n7858) );
  NAND2X0_LVT U9156 ( .A1(n3671), .A2(n_T_427[1117]), .Y(n7857) );
  NAND2X0_LVT U9157 ( .A1(n3992), .A2(n_T_427[1911]), .Y(n7860) );
  NAND2X0_LVT U9158 ( .A1(n3627), .A2(n_T_427[1437]), .Y(n7862) );
  NAND2X0_LVT U9159 ( .A1(n3605), .A2(n_T_427[1373]), .Y(n7861) );
  AND2X1_LVT U9160 ( .A1(n4051), .A2(n_T_427[30]), .Y(n7866) );
  AO22X1_LVT U9161 ( .A1(n4024), .A2(n_T_427[925]), .A3(n4020), .A4(
        n_T_427[670]), .Y(n7865) );
  AO22X1_LVT U9162 ( .A1(n3978), .A2(n_T_427[542]), .A3(n4028), .A4(
        n_T_427[861]), .Y(n7864) );
  AO22X1_LVT U9163 ( .A1(n4034), .A2(n_T_427[606]), .A3(n3985), .A4(
        n_T_427[222]), .Y(n7863) );
  NOR4X1_LVT U9164 ( .A1(n7866), .A2(n7865), .A3(n7864), .A4(n7863), .Y(n7872)
         );
  AO22X1_LVT U9165 ( .A1(n3970), .A2(n_T_427[414]), .A3(n3966), .A4(
        n_T_427[286]), .Y(n7870) );
  AO22X1_LVT U9166 ( .A1(n3974), .A2(n_T_427[158]), .A3(n4037), .A4(
        n_T_427[350]), .Y(n7869) );
  AO22X1_LVT U9167 ( .A1(n3982), .A2(n_T_427[797]), .A3(n4047), .A4(
        n_T_427[734]), .Y(n7868) );
  AO22X1_LVT U9168 ( .A1(n3963), .A2(n_T_427[478]), .A3(n4044), .A4(
        n_T_427[94]), .Y(n7867) );
  NOR4X1_LVT U9169 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .Y(n7871)
         );
  NAND2X0_LVT U9170 ( .A1(n2094), .A2(n_T_427[1310]), .Y(n7876) );
  OA21X1_LVT U9171 ( .A1(n3397), .A2(n3751), .A3(n7876), .Y(n7879) );
  NAND2X0_LVT U9172 ( .A1(n3689), .A2(n_T_427[1694]), .Y(n7878) );
  NAND2X0_LVT U9173 ( .A1(n4001), .A2(n_T_427[1758]), .Y(n7877) );
  NAND2X0_LVT U9174 ( .A1(n3618), .A2(n_T_427[1566]), .Y(n7880) );
  OA21X1_LVT U9175 ( .A1(n3664), .A2(n3296), .A3(n7880), .Y(n7882) );
  NAND2X0_LVT U9176 ( .A1(n4007), .A2(n_T_427[1502]), .Y(n7881) );
  NAND2X0_LVT U9177 ( .A1(n3759), .A2(n_T_427[990]), .Y(n7883) );
  OA21X1_LVT U9178 ( .A1(n4011), .A2(n3297), .A3(n7883), .Y(n7886) );
  NAND2X0_LVT U9179 ( .A1(n3641), .A2(n_T_427[1246]), .Y(n7885) );
  NAND2X0_LVT U9180 ( .A1(n3672), .A2(n_T_427[1118]), .Y(n7884) );
  NAND2X0_LVT U9181 ( .A1(n2985), .A2(n_T_427[1912]), .Y(n7887) );
  OA21X1_LVT U9182 ( .A1(n3767), .A2(n3376), .A3(n7887), .Y(n7890) );
  NAND2X0_LVT U9183 ( .A1(n3630), .A2(n_T_427[1438]), .Y(n7889) );
  NAND2X0_LVT U9184 ( .A1(n_T_427[1374]), .A2(n3611), .Y(n7888) );
  NAND2X0_LVT U9185 ( .A1(n4015), .A2(n4403), .Y(n7902) );
  AND2X1_LVT U9186 ( .A1(n4051), .A2(n_T_427[31]), .Y(n7894) );
  AO22X1_LVT U9187 ( .A1(n4024), .A2(n_T_427[926]), .A3(n4020), .A4(
        n_T_427[671]), .Y(n7893) );
  AO22X1_LVT U9188 ( .A1(n3978), .A2(n_T_427[543]), .A3(n4028), .A4(
        n_T_427[862]), .Y(n7892) );
  AO22X1_LVT U9189 ( .A1(n4034), .A2(n_T_427[607]), .A3(n3985), .A4(
        n_T_427[223]), .Y(n7891) );
  NOR4X1_LVT U9190 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .Y(n7900)
         );
  AO22X1_LVT U9191 ( .A1(n3970), .A2(n_T_427[415]), .A3(n3966), .A4(
        n_T_427[287]), .Y(n7898) );
  AO22X1_LVT U9192 ( .A1(n2858), .A2(n_T_427[159]), .A3(n4037), .A4(
        n_T_427[351]), .Y(n7897) );
  AO22X1_LVT U9193 ( .A1(n3982), .A2(n_T_427[798]), .A3(n4047), .A4(
        n_T_427[735]), .Y(n7896) );
  AO22X1_LVT U9194 ( .A1(n3963), .A2(n_T_427[479]), .A3(n4043), .A4(
        n_T_427[95]), .Y(n7895) );
  NOR4X1_LVT U9195 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .Y(n7899)
         );
  AO21X1_LVT U9196 ( .A1(n7900), .A2(n7899), .A3(n3632), .Y(n7901) );
  AO22X1_LVT U9197 ( .A1(n2497), .A2(n_T_628[31]), .A3(n9064), .A4(
        io_fpu_dmem_resp_data[31]), .Y(n7905) );
  AO22X1_LVT U9198 ( .A1(n9066), .A2(n_T_918[31]), .A3(n9065), .A4(
        io_imem_sfence_bits_addr[31]), .Y(n7904) );
  NAND2X0_LVT U9199 ( .A1(n3757), .A2(n_T_427[991]), .Y(n7906) );
  OA21X1_LVT U9200 ( .A1(n4012), .A2(n3333), .A3(n7906), .Y(n7909) );
  NAND2X0_LVT U9201 ( .A1(n3637), .A2(n_T_427[1247]), .Y(n7908) );
  NAND2X0_LVT U9202 ( .A1(n3672), .A2(n_T_427[1119]), .Y(n7907) );
  AND2X1_LVT U9203 ( .A1(n3976), .A2(n8105), .Y(n9035) );
  NAND2X0_LVT U9204 ( .A1(n3786), .A2(n_T_427[544]), .Y(n7921) );
  NAND2X0_LVT U9205 ( .A1(n3060), .A2(n4406), .Y(n7920) );
  AO22X1_LVT U9206 ( .A1(n4024), .A2(n_T_427[927]), .A3(n4041), .A4(
        n_T_427[96]), .Y(n7917) );
  AO22X1_LVT U9207 ( .A1(n3970), .A2(n_T_427[416]), .A3(n4037), .A4(
        n_T_427[352]), .Y(n7916) );
  AOI22X1_LVT U9208 ( .A1(n4035), .A2(n_T_427[608]), .A3(n4027), .A4(
        n_T_427[863]), .Y(n7914) );
  AOI22X1_LVT U9209 ( .A1(n2858), .A2(n_T_427[160]), .A3(n4051), .A4(
        n_T_427[32]), .Y(n7913) );
  AOI22X1_LVT U9210 ( .A1(n4022), .A2(n_T_427[672]), .A3(n3983), .A4(
        n_T_427[224]), .Y(n7912) );
  NAND3X0_LVT U9211 ( .A1(n7914), .A2(n7913), .A3(n7912), .Y(n7915) );
  OR3X1_LVT U9212 ( .A1(n7917), .A2(n7916), .A3(n7915), .Y(n7918) );
  NAND2X0_LVT U9213 ( .A1(n4053), .A2(n7918), .Y(n7919) );
  AND3X1_LVT U9214 ( .A1(n7921), .A2(n7920), .A3(n7919), .Y(n7924) );
  AND2X1_LVT U9215 ( .A1(n3964), .A2(n8105), .Y(n9053) );
  NAND2X0_LVT U9216 ( .A1(n3789), .A2(n_T_427[288]), .Y(n7922) );
  NAND2X0_LVT U9217 ( .A1(n3689), .A2(n_T_427[1695]), .Y(n7925) );
  OA21X1_LVT U9218 ( .A1(n3143), .A2(n3751), .A3(n7925), .Y(n7928) );
  NAND2X0_LVT U9219 ( .A1(n4000), .A2(n_T_427[1311]), .Y(n7927) );
  NAND2X0_LVT U9220 ( .A1(n2091), .A2(n_T_427[1759]), .Y(n7926) );
  NAND2X0_LVT U9221 ( .A1(n3769), .A2(n_T_427[1503]), .Y(n7929) );
  OA21X1_LVT U9222 ( .A1(n2081), .A2(n3334), .A3(n7929), .Y(n7932) );
  NAND2X0_LVT U9223 ( .A1(n3616), .A2(n_T_427[1567]), .Y(n7931) );
  NAND2X0_LVT U9224 ( .A1(n3652), .A2(n_T_427[1631]), .Y(n7930) );
  NAND2X0_LVT U9225 ( .A1(n9056), .A2(n_T_427[799]), .Y(n7933) );
  OA21X1_LVT U9226 ( .A1(n3398), .A2(n3691), .A3(n7933), .Y(n7938) );
  NAND2X0_LVT U9227 ( .A1(n3629), .A2(n_T_427[1439]), .Y(n7934) );
  NAND2X0_LVT U9228 ( .A1(n3603), .A2(n_T_427[1375]), .Y(n7935) );
  NAND2X0_LVT U9229 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[32]), .Y(n7942) );
  NAND2X0_LVT U9230 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[32]), .Y(n7941)
         );
  NAND2X0_LVT U9231 ( .A1(n2497), .A2(n_T_628[32]), .Y(n7940) );
  NAND2X0_LVT U9232 ( .A1(n9066), .A2(n_T_918[32]), .Y(n7939) );
  NAND4X0_LVT U9233 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .Y(
        io_fpu_fromint_data[32]) );
  NAND2X0_LVT U9234 ( .A1(n3787), .A2(n_T_427[545]), .Y(n7952) );
  NAND2X0_LVT U9235 ( .A1(n3665), .A2(n4408), .Y(n7951) );
  AO22X1_LVT U9236 ( .A1(n4021), .A2(n_T_427[673]), .A3(n3966), .A4(
        n_T_427[289]), .Y(n7948) );
  AO22X1_LVT U9237 ( .A1(n4036), .A2(n_T_427[353]), .A3(n4047), .A4(
        n_T_427[737]), .Y(n7947) );
  AO22X1_LVT U9238 ( .A1(n4024), .A2(n_T_427[928]), .A3(n4031), .A4(
        n_T_427[609]), .Y(n7945) );
  AO22X1_LVT U9239 ( .A1(n2858), .A2(n_T_427[161]), .A3(n4051), .A4(
        n_T_427[33]), .Y(n7944) );
  AO22X1_LVT U9240 ( .A1(n3963), .A2(n_T_427[481]), .A3(n2836), .A4(
        n_T_427[97]), .Y(n7943) );
  OR3X1_LVT U9241 ( .A1(n7945), .A2(n7944), .A3(n7943), .Y(n7946) );
  OR3X1_LVT U9242 ( .A1(n7948), .A2(n7947), .A3(n7946), .Y(n7949) );
  NAND2X0_LVT U9243 ( .A1(n4053), .A2(n7949), .Y(n7950) );
  AND2X1_LVT U9244 ( .A1(n3983), .A2(n8105), .Y(n9058) );
  NAND2X0_LVT U9245 ( .A1(n3624), .A2(n_T_427[225]), .Y(n7954) );
  NAND2X0_LVT U9246 ( .A1(n3661), .A2(n_T_427[864]), .Y(n7953) );
  NAND2X0_LVT U9247 ( .A1(n3635), .A2(n_T_427[1248]), .Y(n7956) );
  NAND2X0_LVT U9248 ( .A1(n3668), .A2(n_T_427[1120]), .Y(n7955) );
  NAND2X0_LVT U9249 ( .A1(n3760), .A2(n_T_427[992]), .Y(n7958) );
  NAND2X0_LVT U9250 ( .A1(n4014), .A2(n_T_427[1056]), .Y(n7957) );
  NAND2X0_LVT U9251 ( .A1(n3605), .A2(n_T_427[1376]), .Y(n7959) );
  NAND2X0_LVT U9252 ( .A1(n2966), .A2(n_T_427[1440]), .Y(n7961) );
  NAND2X0_LVT U9253 ( .A1(n3991), .A2(n_T_427[1913]), .Y(n7960) );
  AND3X1_LVT U9254 ( .A1(n7962), .A2(n7961), .A3(n7960), .Y(n7965) );
  NAND2X0_LVT U9255 ( .A1(n3600), .A2(n_T_427[800]), .Y(n7964) );
  OA21X1_LVT U9256 ( .A1(n3399), .A2(n3601), .A3(n7966), .Y(n7969) );
  NAND2X0_LVT U9257 ( .A1(n2093), .A2(n_T_427[1312]), .Y(n7968) );
  NAND2X0_LVT U9258 ( .A1(n2092), .A2(n_T_427[1760]), .Y(n7967) );
  NAND3X0_LVT U9259 ( .A1(n7969), .A2(n7968), .A3(n7967), .Y(n7974) );
  NAND2X0_LVT U9260 ( .A1(n3769), .A2(n_T_427[1504]), .Y(n7970) );
  NAND2X0_LVT U9261 ( .A1(n3621), .A2(n_T_427[1568]), .Y(n7972) );
  NAND2X0_LVT U9262 ( .A1(n3650), .A2(n_T_427[1632]), .Y(n7971) );
  NAND2X0_LVT U9263 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[33]), .Y(n7978) );
  NAND2X0_LVT U9264 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[33]), .Y(n7977)
         );
  NAND2X0_LVT U9265 ( .A1(n2493), .A2(n_T_628[33]), .Y(n7976) );
  NAND2X0_LVT U9266 ( .A1(n9066), .A2(n_T_918[33]), .Y(n7975) );
  NAND4X0_LVT U9267 ( .A1(n7978), .A2(n7977), .A3(n7976), .A4(n7975), .Y(
        io_fpu_fromint_data[33]) );
  AND2X1_LVT U9268 ( .A1(n4031), .A2(n2135), .Y(n8837) );
  NAND2X0_LVT U9269 ( .A1(n8837), .A2(n_T_427[610]), .Y(n7986) );
  NAND2X0_LVT U9270 ( .A1(n3665), .A2(n4411), .Y(n7985) );
  AO22X1_LVT U9271 ( .A1(n3970), .A2(n_T_427[418]), .A3(n4020), .A4(
        n_T_427[674]), .Y(n7982) );
  AO22X1_LVT U9272 ( .A1(n4024), .A2(n_T_427[929]), .A3(n3986), .A4(
        n_T_427[226]), .Y(n7981) );
  AO22X1_LVT U9273 ( .A1(n2837), .A2(n_T_427[98]), .A3(n4037), .A4(
        n_T_427[354]), .Y(n7980) );
  AO22X1_LVT U9274 ( .A1(n3982), .A2(n_T_427[801]), .A3(n4051), .A4(
        n_T_427[34]), .Y(n7979) );
  NOR4X1_LVT U9275 ( .A1(n7982), .A2(n7981), .A3(n7980), .A4(n7979), .Y(n7983)
         );
  OR2X1_LVT U9276 ( .A1(n7983), .A2(n2154), .Y(n7984) );
  AND3X1_LVT U9277 ( .A1(n7986), .A2(n7985), .A3(n7984), .Y(n7989) );
  NAND2X0_LVT U9278 ( .A1(n3788), .A2(n_T_427[546]), .Y(n7988) );
  NAND2X0_LVT U9279 ( .A1(n_T_427[482]), .A2(n3614), .Y(n7987) );
  NAND2X0_LVT U9280 ( .A1(n8991), .A2(n_T_427[865]), .Y(n7990) );
  OA21X1_LVT U9281 ( .A1(n3691), .A2(n3141), .A3(n7990), .Y(n7993) );
  NAND2X0_LVT U9282 ( .A1(n3790), .A2(n_T_427[290]), .Y(n7992) );
  NAND2X0_LVT U9283 ( .A1(n3713), .A2(n_T_427[162]), .Y(n7991) );
  NAND2X0_LVT U9284 ( .A1(n3605), .A2(n_T_427[1377]), .Y(n7994) );
  OA21X1_LVT U9285 ( .A1(n3452), .A2(n3767), .A3(n7994), .Y(n7997) );
  NAND2X0_LVT U9286 ( .A1(n3628), .A2(n_T_427[1441]), .Y(n7996) );
  NAND2X0_LVT U9287 ( .A1(n2998), .A2(n_T_427[1914]), .Y(n7995) );
  NAND2X0_LVT U9288 ( .A1(n2922), .A2(n_T_427[1697]), .Y(n7998) );
  OA21X1_LVT U9289 ( .A1(n3453), .A2(n3601), .A3(n7998), .Y(n8001) );
  NAND2X0_LVT U9290 ( .A1(n2094), .A2(n_T_427[1313]), .Y(n8000) );
  NAND2X0_LVT U9291 ( .A1(n4003), .A2(n_T_427[1761]), .Y(n7999) );
  NAND2X0_LVT U9292 ( .A1(n3769), .A2(n_T_427[1505]), .Y(n8002) );
  OA21X1_LVT U9293 ( .A1(n4010), .A2(n3335), .A3(n8002), .Y(n8005) );
  NAND2X0_LVT U9294 ( .A1(n3619), .A2(n_T_427[1569]), .Y(n8004) );
  NAND2X0_LVT U9295 ( .A1(n_T_427[1633]), .A2(n3643), .Y(n8003) );
  NAND2X0_LVT U9296 ( .A1(n_T_427[1249]), .A2(n3641), .Y(n8007) );
  NAND2X0_LVT U9297 ( .A1(n3674), .A2(n_T_427[1121]), .Y(n8006) );
  NAND2X0_LVT U9298 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[34]), .Y(n8012) );
  NAND2X0_LVT U9299 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[34]), .Y(n8011)
         );
  NAND2X0_LVT U9300 ( .A1(n2493), .A2(n_T_628[34]), .Y(n8010) );
  NAND2X0_LVT U9301 ( .A1(n9066), .A2(n_T_918[34]), .Y(n8009) );
  NAND4X0_LVT U9302 ( .A1(n8012), .A2(n8011), .A3(n8010), .A4(n8009), .Y(
        io_fpu_fromint_data[34]) );
  NAND2X0_LVT U9303 ( .A1(n3661), .A2(n_T_427[866]), .Y(n8013) );
  OA21X1_LVT U9304 ( .A1(n3400), .A2(n3691), .A3(n8013), .Y(n8022) );
  AO22X1_LVT U9305 ( .A1(n4024), .A2(n_T_427[930]), .A3(n3960), .A4(
        n_T_427[483]), .Y(n8017) );
  AO22X1_LVT U9306 ( .A1(n3967), .A2(n_T_427[291]), .A3(n4037), .A4(
        n_T_427[355]), .Y(n8016) );
  AO22X1_LVT U9307 ( .A1(n3975), .A2(n_T_427[163]), .A3(n4052), .A4(
        n_T_427[35]), .Y(n8015) );
  AO22X1_LVT U9308 ( .A1(n4034), .A2(n_T_427[611]), .A3(n3986), .A4(
        n_T_427[227]), .Y(n8014) );
  NOR4X1_LVT U9309 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .Y(n8019)
         );
  NAND2X0_LVT U9310 ( .A1(n2982), .A2(n4413), .Y(n8018) );
  OA21X1_LVT U9311 ( .A1(n8019), .A2(n3612), .A3(n8018), .Y(n8021) );
  NAND2X0_LVT U9312 ( .A1(n3788), .A2(n_T_427[547]), .Y(n8020) );
  NAND2X0_LVT U9313 ( .A1(n2135), .A2(n4022), .Y(n8996) );
  NAND2X0_LVT U9314 ( .A1(n_T_427[99]), .A2(n3707), .Y(n8023) );
  OA21X1_LVT U9315 ( .A1(n3369), .A2(n8996), .A3(n8023), .Y(n8026) );
  NAND2X0_LVT U9316 ( .A1(n3600), .A2(n_T_427[802]), .Y(n8024) );
  NAND2X0_LVT U9317 ( .A1(n3609), .A2(n_T_427[1378]), .Y(n8027) );
  NAND2X0_LVT U9318 ( .A1(n2966), .A2(n_T_427[1442]), .Y(n8029) );
  NAND2X0_LVT U9319 ( .A1(n2882), .A2(n_T_427[1915]), .Y(n8028) );
  NAND2X0_LVT U9320 ( .A1(n2922), .A2(n_T_427[1698]), .Y(n8031) );
  OA21X1_LVT U9321 ( .A1(n3401), .A2(n3601), .A3(n8031), .Y(n8034) );
  NAND2X0_LVT U9322 ( .A1(n2094), .A2(n_T_427[1314]), .Y(n8033) );
  NAND2X0_LVT U9323 ( .A1(n2092), .A2(n_T_427[1762]), .Y(n8032) );
  NAND2X0_LVT U9324 ( .A1(n3769), .A2(n_T_427[1506]), .Y(n8035) );
  OA21X1_LVT U9325 ( .A1(n2081), .A2(n3299), .A3(n8035), .Y(n8038) );
  NAND2X0_LVT U9326 ( .A1(n3618), .A2(n_T_427[1570]), .Y(n8037) );
  NAND2X0_LVT U9327 ( .A1(n3648), .A2(n_T_427[1634]), .Y(n8036) );
  NAND2X0_LVT U9328 ( .A1(n_T_427[1250]), .A2(n3635), .Y(n8040) );
  NAND2X0_LVT U9329 ( .A1(n3674), .A2(n_T_427[1122]), .Y(n8039) );
  NAND2X0_LVT U9330 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[35]), .Y(n8045) );
  NAND2X0_LVT U9331 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[35]), .Y(n8044)
         );
  NAND2X0_LVT U9332 ( .A1(n2493), .A2(n_T_628[35]), .Y(n8043) );
  NAND2X0_LVT U9333 ( .A1(n9066), .A2(n_T_918[35]), .Y(n8042) );
  NAND4X0_LVT U9334 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .Y(
        io_fpu_fromint_data[35]) );
  NAND2X0_LVT U9335 ( .A1(n2967), .A2(n_T_427[1443]), .Y(n8047) );
  AND3X1_LVT U9336 ( .A1(n8048), .A2(n8047), .A3(n8046), .Y(n8051) );
  NAND2X0_LVT U9337 ( .A1(n3789), .A2(n_T_427[292]), .Y(n8050) );
  NAND2X0_LVT U9338 ( .A1(n3771), .A2(n_T_427[739]), .Y(n8049) );
  NAND2X0_LVT U9339 ( .A1(n3998), .A2(n_T_427[1315]), .Y(n8053) );
  NAND2X0_LVT U9340 ( .A1(n4003), .A2(n_T_427[1763]), .Y(n8052) );
  NAND3X0_LVT U9341 ( .A1(n8053), .A2(n8052), .A3(n8054), .Y(n8060) );
  NAND2X0_LVT U9342 ( .A1(n2922), .A2(n_T_427[1699]), .Y(n8055) );
  OA21X1_LVT U9343 ( .A1(n3753), .A2(n3454), .A3(n8055), .Y(n8058) );
  NAND2X0_LVT U9344 ( .A1(n3620), .A2(n_T_427[1571]), .Y(n8057) );
  NAND2X0_LVT U9345 ( .A1(n_T_427[1635]), .A2(n3650), .Y(n8056) );
  NAND3X0_LVT U9346 ( .A1(n8058), .A2(n8057), .A3(n8056), .Y(n8059) );
  NAND2X0_LVT U9347 ( .A1(n3673), .A2(n_T_427[1123]), .Y(n8062) );
  NAND2X0_LVT U9348 ( .A1(n3759), .A2(n_T_427[995]), .Y(n8061) );
  NAND2X0_LVT U9349 ( .A1(n8062), .A2(n8061), .Y(n8079) );
  NAND2X0_LVT U9350 ( .A1(n3661), .A2(n_T_427[867]), .Y(n8073) );
  AO22X1_LVT U9351 ( .A1(n4039), .A2(n_T_427[356]), .A3(n4041), .A4(
        n_T_427[100]), .Y(n8069) );
  AO22X1_LVT U9352 ( .A1(n3973), .A2(n_T_427[164]), .A3(n3979), .A4(
        n_T_427[803]), .Y(n8068) );
  AOI22X1_LVT U9353 ( .A1(n4025), .A2(n_T_427[931]), .A3(n4031), .A4(
        n_T_427[612]), .Y(n8066) );
  AOI22X1_LVT U9354 ( .A1(n4022), .A2(n_T_427[676]), .A3(n3976), .A4(
        n_T_427[548]), .Y(n8065) );
  AOI22X1_LVT U9355 ( .A1(n3971), .A2(n_T_427[420]), .A3(n3960), .A4(
        n_T_427[484]), .Y(n8064) );
  NAND2X0_LVT U9356 ( .A1(n4052), .A2(n_T_427[36]), .Y(n8063) );
  NAND4X0_LVT U9357 ( .A1(n8066), .A2(n8065), .A3(n8064), .A4(n8063), .Y(n8067) );
  OR3X1_LVT U9358 ( .A1(n8069), .A2(n8068), .A3(n8067), .Y(n8070) );
  NAND2X0_LVT U9359 ( .A1(n4053), .A2(n8070), .Y(n8071) );
  NAND3X0_LVT U9360 ( .A1(n8073), .A2(n8072), .A3(n8071), .Y(n8078) );
  NAND2X0_LVT U9361 ( .A1(n3635), .A2(n_T_427[1251]), .Y(n8074) );
  NAND2X0_LVT U9362 ( .A1(n4014), .A2(n_T_427[1059]), .Y(n8075) );
  NAND2X0_LVT U9363 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[36]), .Y(n8084) );
  NAND2X0_LVT U9364 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[36]), .Y(n8083)
         );
  NAND2X0_LVT U9365 ( .A1(n2497), .A2(n_T_628[36]), .Y(n8082) );
  NAND2X0_LVT U9366 ( .A1(n9066), .A2(n_T_918[36]), .Y(n8081) );
  NAND4X0_LVT U9367 ( .A1(n8084), .A2(n8083), .A3(n8082), .A4(n8081), .Y(
        io_fpu_fromint_data[36]) );
  NAND2X0_LVT U9368 ( .A1(n3789), .A2(n_T_427[293]), .Y(n8094) );
  NAND2X0_LVT U9369 ( .A1(n3060), .A2(n4419), .Y(n8093) );
  AO22X1_LVT U9370 ( .A1(n8980), .A2(n_T_427[549]), .A3(n4043), .A4(
        n_T_427[101]), .Y(n8090) );
  AO22X1_LVT U9371 ( .A1(n4021), .A2(n_T_427[677]), .A3(n4037), .A4(
        n_T_427[357]), .Y(n8089) );
  AO22X1_LVT U9372 ( .A1(n4024), .A2(n_T_427[932]), .A3(n3960), .A4(
        n_T_427[485]), .Y(n8087) );
  AO22X1_LVT U9373 ( .A1(n3982), .A2(n_T_427[804]), .A3(n4047), .A4(
        n_T_427[740]), .Y(n8086) );
  AO22X1_LVT U9374 ( .A1(n4034), .A2(n_T_427[613]), .A3(n4028), .A4(
        n_T_427[868]), .Y(n8085) );
  OR3X1_LVT U9375 ( .A1(n8087), .A2(n8086), .A3(n8085), .Y(n8088) );
  OR3X1_LVT U9376 ( .A1(n8090), .A2(n8089), .A3(n8088), .Y(n8091) );
  NAND2X0_LVT U9377 ( .A1(n4053), .A2(n8091), .Y(n8092) );
  NAND2X0_LVT U9378 ( .A1(n3745), .A2(n_T_427[229]), .Y(n8096) );
  NAND2X0_LVT U9379 ( .A1(n3713), .A2(n_T_427[165]), .Y(n8095) );
  NAND2X0_LVT U9380 ( .A1(n3635), .A2(n_T_427[1252]), .Y(n8098) );
  NAND2X0_LVT U9381 ( .A1(n3670), .A2(n_T_427[1124]), .Y(n8097) );
  NAND2X0_LVT U9382 ( .A1(n3761), .A2(n_T_427[996]), .Y(n8100) );
  NAND2X0_LVT U9383 ( .A1(n3716), .A2(n_T_427[1060]), .Y(n8099) );
  NAND2X0_LVT U9384 ( .A1(n3607), .A2(n_T_427[1380]), .Y(n8101) );
  NAND2X0_LVT U9385 ( .A1(n3630), .A2(n_T_427[1444]), .Y(n8103) );
  NAND2X0_LVT U9386 ( .A1(n2985), .A2(n_T_427[1917]), .Y(n8102) );
  AND3X1_LVT U9387 ( .A1(n8104), .A2(n8103), .A3(n8102), .Y(n8108) );
  NAND2X0_LVT U9388 ( .A1(n3647), .A2(n_T_427[37]), .Y(n8107) );
  NAND2X0_LVT U9389 ( .A1(n3689), .A2(n_T_427[1700]), .Y(n8109) );
  OA21X1_LVT U9390 ( .A1(n3456), .A2(n3601), .A3(n8109), .Y(n8112) );
  NAND2X0_LVT U9391 ( .A1(n4000), .A2(n_T_427[1316]), .Y(n8111) );
  NAND2X0_LVT U9392 ( .A1(n4001), .A2(n_T_427[1764]), .Y(n8110) );
  NAND2X0_LVT U9393 ( .A1(n3769), .A2(n_T_427[1508]), .Y(n8113) );
  NAND2X0_LVT U9394 ( .A1(n3618), .A2(n_T_427[1572]), .Y(n8115) );
  NAND2X0_LVT U9395 ( .A1(n3642), .A2(n_T_427[1636]), .Y(n8114) );
  NAND2X0_LVT U9396 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[37]), .Y(n8120) );
  NAND2X0_LVT U9397 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[37]), .Y(n8119)
         );
  NAND2X0_LVT U9398 ( .A1(n2493), .A2(n_T_628[37]), .Y(n8118) );
  NAND2X0_LVT U9399 ( .A1(n9066), .A2(n_T_918[37]), .Y(n8117) );
  NAND4X0_LVT U9400 ( .A1(n8120), .A2(n8119), .A3(n8118), .A4(n8117), .Y(
        io_fpu_fromint_data[37]) );
  NAND2X0_LVT U9401 ( .A1(n8994), .A2(n_T_427[102]), .Y(n8123) );
  NAND2X0_LVT U9402 ( .A1(n3630), .A2(n_T_427[1445]), .Y(n8122) );
  NAND2X0_LVT U9403 ( .A1(n2985), .A2(n_T_427[1918]), .Y(n8121) );
  AND3X1_LVT U9404 ( .A1(n8123), .A2(n8122), .A3(n8121), .Y(n8126) );
  NAND2X0_LVT U9405 ( .A1(n3771), .A2(n_T_427[741]), .Y(n8124) );
  NAND2X0_LVT U9406 ( .A1(n3606), .A2(n_T_427[1381]), .Y(n8127) );
  OA21X1_LVT U9407 ( .A1(n3481), .A2(n9006), .A3(n8127), .Y(n8130) );
  NAND2X0_LVT U9408 ( .A1(n3999), .A2(n_T_427[1317]), .Y(n8129) );
  NAND2X0_LVT U9409 ( .A1(n4001), .A2(n_T_427[1765]), .Y(n8128) );
  OA21X1_LVT U9410 ( .A1(n3402), .A2(n3753), .A3(n8131), .Y(n8134) );
  NAND2X0_LVT U9411 ( .A1(n3621), .A2(n_T_427[1573]), .Y(n8133) );
  NAND2X0_LVT U9412 ( .A1(n3642), .A2(n_T_427[1637]), .Y(n8132) );
  NAND2X0_LVT U9413 ( .A1(n3670), .A2(n_T_427[1125]), .Y(n8136) );
  NAND2X0_LVT U9414 ( .A1(n3756), .A2(n_T_427[997]), .Y(n8135) );
  NAND2X0_LVT U9415 ( .A1(n3714), .A2(n_T_427[166]), .Y(n8147) );
  NAND2X0_LVT U9416 ( .A1(n2982), .A2(n4421), .Y(n8146) );
  AO22X1_LVT U9417 ( .A1(n3970), .A2(n_T_427[422]), .A3(n4037), .A4(
        n_T_427[358]), .Y(n8143) );
  AO22X1_LVT U9418 ( .A1(n3967), .A2(n_T_427[294]), .A3(n3979), .A4(
        n_T_427[805]), .Y(n8142) );
  AOI22X1_LVT U9419 ( .A1(n4035), .A2(n_T_427[614]), .A3(n4027), .A4(
        n_T_427[869]), .Y(n8140) );
  AOI22X1_LVT U9420 ( .A1(n3978), .A2(n_T_427[550]), .A3(n3983), .A4(
        n_T_427[230]), .Y(n8139) );
  AOI22X1_LVT U9421 ( .A1(n4024), .A2(n_T_427[933]), .A3(n4018), .A4(
        n_T_427[678]), .Y(n8138) );
  NAND2X0_LVT U9422 ( .A1(n4052), .A2(n_T_427[38]), .Y(n8137) );
  NAND4X0_LVT U9423 ( .A1(n8140), .A2(n8139), .A3(n8138), .A4(n8137), .Y(n8141) );
  OR3X1_LVT U9424 ( .A1(n8143), .A2(n8142), .A3(n8141), .Y(n8144) );
  NAND2X0_LVT U9425 ( .A1(n4053), .A2(n8144), .Y(n8145) );
  NAND2X0_LVT U9426 ( .A1(n3635), .A2(n_T_427[1253]), .Y(n8148) );
  NAND2X0_LVT U9427 ( .A1(n2611), .A2(n_T_427[1189]), .Y(n8150) );
  NAND2X0_LVT U9428 ( .A1(n3716), .A2(n_T_427[1061]), .Y(n8149) );
  NAND2X0_LVT U9429 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[38]), .Y(n8154) );
  NAND2X0_LVT U9430 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[38]), .Y(n8153)
         );
  NAND2X0_LVT U9431 ( .A1(n2497), .A2(n_T_628[38]), .Y(n8152) );
  NAND2X0_LVT U9432 ( .A1(n9066), .A2(n_T_918[38]), .Y(n8151) );
  NAND4X0_LVT U9433 ( .A1(n8154), .A2(n8153), .A3(n8152), .A4(n8151), .Y(
        io_fpu_fromint_data[38]) );
  NAND2X0_LVT U9434 ( .A1(n3626), .A2(n_T_427[1446]), .Y(n8156) );
  NAND2X0_LVT U9435 ( .A1(n2986), .A2(n_T_427[1919]), .Y(n8155) );
  AND3X1_LVT U9436 ( .A1(n8157), .A2(n8156), .A3(n8155), .Y(n8160) );
  NAND2X0_LVT U9437 ( .A1(n3789), .A2(n_T_427[295]), .Y(n8159) );
  NAND2X0_LVT U9438 ( .A1(n3647), .A2(n_T_427[39]), .Y(n8158) );
  NAND2X0_LVT U9439 ( .A1(n3606), .A2(n_T_427[1382]), .Y(n8161) );
  OA21X1_LVT U9440 ( .A1(n3457), .A2(n9006), .A3(n8161), .Y(n8164) );
  NAND2X0_LVT U9441 ( .A1(n4000), .A2(n_T_427[1318]), .Y(n8163) );
  NAND2X0_LVT U9442 ( .A1(n2091), .A2(n_T_427[1766]), .Y(n8162) );
  NAND2X0_LVT U9443 ( .A1(n3689), .A2(n_T_427[1702]), .Y(n8165) );
  OA21X1_LVT U9444 ( .A1(n3458), .A2(n3753), .A3(n8165), .Y(n8168) );
  NAND2X0_LVT U9445 ( .A1(n3615), .A2(n_T_427[1574]), .Y(n8167) );
  NAND2X0_LVT U9446 ( .A1(n3649), .A2(n_T_427[1638]), .Y(n8166) );
  NAND2X0_LVT U9447 ( .A1(n3672), .A2(n_T_427[1126]), .Y(n8170) );
  NAND2X0_LVT U9448 ( .A1(n3757), .A2(n_T_427[998]), .Y(n8169) );
  NAND2X0_LVT U9449 ( .A1(n_T_427[167]), .A2(n3713), .Y(n8181) );
  NAND2X0_LVT U9450 ( .A1(n4015), .A2(n4424), .Y(n8180) );
  AO22X1_LVT U9451 ( .A1(n4021), .A2(n_T_427[679]), .A3(n4042), .A4(
        n_T_427[103]), .Y(n8177) );
  AO22X1_LVT U9452 ( .A1(n3982), .A2(n_T_427[806]), .A3(n4037), .A4(
        n_T_427[359]), .Y(n8176) );
  AOI22X1_LVT U9453 ( .A1(n4035), .A2(n_T_427[615]), .A3(n4027), .A4(
        n_T_427[870]), .Y(n8174) );
  AOI22X1_LVT U9454 ( .A1(n3978), .A2(n_T_427[551]), .A3(n3983), .A4(
        n_T_427[231]), .Y(n8173) );
  AOI22X1_LVT U9455 ( .A1(n4026), .A2(n_T_427[934]), .A3(n3960), .A4(
        n_T_427[487]), .Y(n8172) );
  NAND2X0_LVT U9456 ( .A1(n4048), .A2(n_T_427[742]), .Y(n8171) );
  NAND4X0_LVT U9457 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .Y(n8175) );
  OR3X1_LVT U9458 ( .A1(n8177), .A2(n8176), .A3(n8175), .Y(n8178) );
  NAND2X0_LVT U9459 ( .A1(n4053), .A2(n8178), .Y(n8179) );
  NAND2X0_LVT U9460 ( .A1(n3640), .A2(n_T_427[1254]), .Y(n8182) );
  NAND2X0_LVT U9461 ( .A1(n2611), .A2(n_T_427[1190]), .Y(n8184) );
  NAND2X0_LVT U9462 ( .A1(n3717), .A2(n_T_427[1062]), .Y(n8183) );
  NAND2X0_LVT U9463 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[39]), .Y(n8188) );
  NAND2X0_LVT U9464 ( .A1(n9065), .A2(n_T_1165[39]), .Y(n8187) );
  NAND2X0_LVT U9465 ( .A1(n2493), .A2(n_T_628[39]), .Y(n8186) );
  NAND2X0_LVT U9466 ( .A1(n9066), .A2(n_T_918[39]), .Y(n8185) );
  NAND4X0_LVT U9467 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .Y(
        io_fpu_fromint_data[39]) );
  NAND2X0_LVT U9468 ( .A1(n_T_427[1383]), .A2(n3611), .Y(n8189) );
  OA21X1_LVT U9469 ( .A1(n3147), .A2(n3988), .A3(n8189), .Y(n8192) );
  NAND2X0_LVT U9470 ( .A1(n2967), .A2(n_T_427[1447]), .Y(n8191) );
  NAND2X0_LVT U9471 ( .A1(n3992), .A2(n_T_427[1920]), .Y(n8190) );
  NAND3X0_LVT U9472 ( .A1(n8192), .A2(n8191), .A3(n8190), .Y(n8197) );
  NAND2X0_LVT U9473 ( .A1(n3657), .A2(n_T_427[1703]), .Y(n8193) );
  NAND2X0_LVT U9474 ( .A1(n3998), .A2(n_T_427[1319]), .Y(n8195) );
  NAND2X0_LVT U9475 ( .A1(n4003), .A2(n_T_427[1767]), .Y(n8194) );
  NAND2X0_LVT U9476 ( .A1(n3769), .A2(n_T_427[1511]), .Y(n8198) );
  OA21X1_LVT U9477 ( .A1(n4008), .A2(n3337), .A3(n8198), .Y(n8201) );
  NAND2X0_LVT U9478 ( .A1(n3621), .A2(n_T_427[1575]), .Y(n8200) );
  NAND2X0_LVT U9479 ( .A1(n3642), .A2(n_T_427[1639]), .Y(n8199) );
  NAND3X0_LVT U9480 ( .A1(n8201), .A2(n8200), .A3(n8199), .Y(n8206) );
  NAND2X0_LVT U9481 ( .A1(n3760), .A2(n_T_427[999]), .Y(n8202) );
  NAND2X0_LVT U9482 ( .A1(n_T_427[1255]), .A2(n3638), .Y(n8204) );
  NAND2X0_LVT U9483 ( .A1(n3668), .A2(n_T_427[1127]), .Y(n8203) );
  NAND2X0_LVT U9484 ( .A1(n3786), .A2(n_T_427[552]), .Y(n8214) );
  NAND2X0_LVT U9485 ( .A1(n3060), .A2(n4427), .Y(n8213) );
  AO22X1_LVT U9486 ( .A1(n4024), .A2(n_T_427[935]), .A3(n3960), .A4(
        n_T_427[488]), .Y(n8210) );
  AO22X1_LVT U9487 ( .A1(n4021), .A2(n_T_427[680]), .A3(n2836), .A4(
        n_T_427[104]), .Y(n8209) );
  AO22X1_LVT U9488 ( .A1(n3982), .A2(n_T_427[807]), .A3(n4037), .A4(
        n_T_427[360]), .Y(n8208) );
  AO22X1_LVT U9489 ( .A1(n4034), .A2(n_T_427[616]), .A3(n3986), .A4(
        n_T_427[232]), .Y(n8207) );
  NOR4X1_LVT U9490 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .Y(n8211)
         );
  OR2X1_LVT U9491 ( .A1(n8211), .A2(n3656), .Y(n8212) );
  NAND3X0_LVT U9492 ( .A1(n8214), .A2(n8213), .A3(n8212), .Y(n8222) );
  NAND2X0_LVT U9493 ( .A1(n3661), .A2(n_T_427[871]), .Y(n8216) );
  NAND2X0_LVT U9494 ( .A1(n3790), .A2(n_T_427[296]), .Y(n8215) );
  NAND2X0_LVT U9495 ( .A1(n8216), .A2(n8215), .Y(n8221) );
  NAND2X0_LVT U9496 ( .A1(n_T_427[168]), .A2(n3791), .Y(n8217) );
  OA21X1_LVT U9497 ( .A1(n3461), .A2(n3708), .A3(n8217), .Y(n8220) );
  NAND2X0_LVT U9498 ( .A1(n8944), .A2(n_T_427[40]), .Y(n8218) );
  NAND2X0_LVT U9499 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[40]), .Y(n8226) );
  NAND2X0_LVT U9500 ( .A1(n9065), .A2(n_T_1165[40]), .Y(n8225) );
  NAND2X0_LVT U9501 ( .A1(n2493), .A2(n_T_628[40]), .Y(n8224) );
  NAND2X0_LVT U9502 ( .A1(n9066), .A2(n_T_918[40]), .Y(n8223) );
  NAND4X0_LVT U9503 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8223), .Y(
        io_fpu_fromint_data[40]) );
  NAND2X0_LVT U9504 ( .A1(n_T_427[489]), .A2(n9052), .Y(n8228) );
  NAND2X0_LVT U9505 ( .A1(n3790), .A2(n_T_427[297]), .Y(n8227) );
  AND2X1_LVT U9506 ( .A1(n8228), .A2(n8227), .Y(n8237) );
  AO22X1_LVT U9507 ( .A1(n3970), .A2(n_T_427[425]), .A3(n4023), .A4(
        n_T_427[936]), .Y(n8232) );
  AO22X1_LVT U9508 ( .A1(n3982), .A2(n_T_427[808]), .A3(n4048), .A4(
        n_T_427[744]), .Y(n8231) );
  AO22X1_LVT U9509 ( .A1(n4034), .A2(n_T_427[617]), .A3(n3986), .A4(
        n_T_427[233]), .Y(n8230) );
  AO22X1_LVT U9510 ( .A1(n2836), .A2(n_T_427[105]), .A3(n4037), .A4(
        n_T_427[361]), .Y(n8229) );
  NOR4X1_LVT U9511 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8229), .Y(n8234)
         );
  NAND2X0_LVT U9512 ( .A1(n3060), .A2(n4430), .Y(n8233) );
  OA21X1_LVT U9513 ( .A1(n8234), .A2(n3612), .A3(n8233), .Y(n8236) );
  NAND2X0_LVT U9514 ( .A1(n3786), .A2(n_T_427[553]), .Y(n8235) );
  NAND2X0_LVT U9515 ( .A1(n8944), .A2(n_T_427[41]), .Y(n8238) );
  OA21X1_LVT U9516 ( .A1(n3404), .A2(n8996), .A3(n8238), .Y(n8241) );
  NAND2X0_LVT U9517 ( .A1(n3714), .A2(n_T_427[169]), .Y(n8240) );
  NAND2X0_LVT U9518 ( .A1(n8991), .A2(n_T_427[872]), .Y(n8239) );
  NAND2X0_LVT U9519 ( .A1(n3605), .A2(n_T_427[1384]), .Y(n8242) );
  NAND2X0_LVT U9520 ( .A1(n3627), .A2(n_T_427[1448]), .Y(n8244) );
  NAND2X0_LVT U9521 ( .A1(n2986), .A2(n_T_427[1921]), .Y(n8243) );
  NAND2X0_LVT U9522 ( .A1(n2093), .A2(n_T_427[1320]), .Y(n8248) );
  NAND2X0_LVT U9523 ( .A1(n4004), .A2(n_T_427[1768]), .Y(n8247) );
  NAND2X0_LVT U9524 ( .A1(n3770), .A2(n_T_427[1512]), .Y(n8250) );
  NAND2X0_LVT U9525 ( .A1(n_T_427[1576]), .A2(n3617), .Y(n8252) );
  NAND2X0_LVT U9526 ( .A1(n3650), .A2(n_T_427[1640]), .Y(n8251) );
  NAND2X0_LVT U9527 ( .A1(n_T_427[1256]), .A2(n3640), .Y(n8255) );
  NAND2X0_LVT U9528 ( .A1(n3668), .A2(n_T_427[1128]), .Y(n8254) );
  NAND2X0_LVT U9529 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[41]), .Y(n8260) );
  NAND2X0_LVT U9530 ( .A1(n9065), .A2(n_T_1165[41]), .Y(n8259) );
  NAND2X0_LVT U9531 ( .A1(n2497), .A2(n_T_628[41]), .Y(n8258) );
  NAND2X0_LVT U9532 ( .A1(n9066), .A2(n_T_918[41]), .Y(n8257) );
  NAND4X0_LVT U9533 ( .A1(n8260), .A2(n8259), .A3(n8258), .A4(n8257), .Y(
        io_fpu_fromint_data[41]) );
  NAND2X0_LVT U9534 ( .A1(n3771), .A2(n_T_427[745]), .Y(n8263) );
  NAND2X0_LVT U9535 ( .A1(n2966), .A2(n_T_427[1449]), .Y(n8262) );
  NAND2X0_LVT U9536 ( .A1(n2998), .A2(n_T_427[1922]), .Y(n8261) );
  AND3X1_LVT U9537 ( .A1(n8263), .A2(n8262), .A3(n8261), .Y(n8266) );
  NAND2X0_LVT U9538 ( .A1(n3787), .A2(n_T_427[554]), .Y(n8265) );
  NAND2X0_LVT U9539 ( .A1(n_T_427[1385]), .A2(n3611), .Y(n8267) );
  OA21X1_LVT U9540 ( .A1(n3149), .A2(n3989), .A3(n8267), .Y(n8270) );
  NAND2X0_LVT U9541 ( .A1(n3998), .A2(n_T_427[1321]), .Y(n8269) );
  NAND2X0_LVT U9542 ( .A1(n4003), .A2(n_T_427[1769]), .Y(n8268) );
  NAND3X0_LVT U9543 ( .A1(n8268), .A2(n8269), .A3(n8270), .Y(n8276) );
  NAND2X0_LVT U9544 ( .A1(n_T_427[1705]), .A2(n3689), .Y(n8271) );
  OA21X1_LVT U9545 ( .A1(n3462), .A2(n3753), .A3(n8271), .Y(n8274) );
  NAND2X0_LVT U9546 ( .A1(n3621), .A2(n_T_427[1577]), .Y(n8273) );
  NAND3X0_LVT U9547 ( .A1(n8274), .A2(n8273), .A3(n8272), .Y(n8275) );
  NAND2X0_LVT U9548 ( .A1(n3671), .A2(n_T_427[1129]), .Y(n8278) );
  NAND2X0_LVT U9549 ( .A1(n3712), .A2(n_T_427[1001]), .Y(n8277) );
  NAND2X0_LVT U9550 ( .A1(n4015), .A2(n4433), .Y(n8288) );
  AO22X1_LVT U9551 ( .A1(n4039), .A2(n_T_427[362]), .A3(n4044), .A4(
        n_T_427[106]), .Y(n8285) );
  AO22X1_LVT U9552 ( .A1(n2859), .A2(n_T_427[170]), .A3(n3979), .A4(
        n_T_427[809]), .Y(n8284) );
  AOI22X1_LVT U9553 ( .A1(n4035), .A2(n_T_427[618]), .A3(n4027), .A4(
        n_T_427[873]), .Y(n8282) );
  AOI22X1_LVT U9554 ( .A1(n4022), .A2(n_T_427[682]), .A3(n3983), .A4(
        n_T_427[234]), .Y(n8281) );
  AOI22X1_LVT U9555 ( .A1(n3971), .A2(n_T_427[426]), .A3(n4023), .A4(
        n_T_427[937]), .Y(n8280) );
  NAND2X0_LVT U9556 ( .A1(n4052), .A2(n_T_427[42]), .Y(n8279) );
  NAND4X0_LVT U9557 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8279), .Y(n8283) );
  OR3X1_LVT U9558 ( .A1(n8285), .A2(n8284), .A3(n8283), .Y(n8286) );
  NAND2X0_LVT U9559 ( .A1(n4053), .A2(n8286), .Y(n8287) );
  NAND2X0_LVT U9560 ( .A1(n_T_427[1257]), .A2(n3640), .Y(n8290) );
  OA21X1_LVT U9561 ( .A1(n3463), .A2(n2897), .A3(n8290), .Y(n8293) );
  NAND2X0_LVT U9562 ( .A1(n2611), .A2(n_T_427[1193]), .Y(n8292) );
  NAND2X0_LVT U9563 ( .A1(n4014), .A2(n_T_427[1065]), .Y(n8291) );
  NAND2X0_LVT U9564 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[42]), .Y(n8297) );
  NAND2X0_LVT U9565 ( .A1(n9065), .A2(n_T_1165[42]), .Y(n8296) );
  NAND2X0_LVT U9566 ( .A1(n2497), .A2(n_T_628[42]), .Y(n8295) );
  NAND2X0_LVT U9567 ( .A1(n9066), .A2(n_T_918[42]), .Y(n8294) );
  NAND4X0_LVT U9568 ( .A1(n8297), .A2(n8296), .A3(n8295), .A4(n8294), .Y(
        io_fpu_fromint_data[42]) );
  NAND2X0_LVT U9569 ( .A1(n3609), .A2(n_T_427[1386]), .Y(n8298) );
  OA21X1_LVT U9570 ( .A1(n3150), .A2(n3989), .A3(n8298), .Y(n8301) );
  NAND2X0_LVT U9571 ( .A1(n2967), .A2(n_T_427[1450]), .Y(n8300) );
  NAND2X0_LVT U9572 ( .A1(n3991), .A2(n_T_427[1923]), .Y(n8299) );
  NAND2X0_LVT U9573 ( .A1(n3689), .A2(n_T_427[1706]), .Y(n8302) );
  OA21X1_LVT U9574 ( .A1(n3464), .A2(n3994), .A3(n8302), .Y(n8305) );
  NAND2X0_LVT U9575 ( .A1(n3998), .A2(n_T_427[1322]), .Y(n8304) );
  NAND2X0_LVT U9576 ( .A1(n2091), .A2(n_T_427[1770]), .Y(n8303) );
  NAND2X0_LVT U9577 ( .A1(n3769), .A2(n_T_427[1514]), .Y(n8306) );
  OA21X1_LVT U9578 ( .A1(n4008), .A2(n3340), .A3(n8306), .Y(n8309) );
  NAND2X0_LVT U9579 ( .A1(n3616), .A2(n_T_427[1578]), .Y(n8308) );
  NAND2X0_LVT U9580 ( .A1(n_T_427[1642]), .A2(n3648), .Y(n8307) );
  NAND3X0_LVT U9581 ( .A1(n8307), .A2(n8308), .A3(n8309), .Y(n8314) );
  NAND2X0_LVT U9582 ( .A1(n3757), .A2(n_T_427[1002]), .Y(n8310) );
  NAND2X0_LVT U9583 ( .A1(n3637), .A2(n_T_427[1258]), .Y(n8312) );
  NAND2X0_LVT U9584 ( .A1(n3670), .A2(n_T_427[1130]), .Y(n8311) );
  NAND2X0_LVT U9585 ( .A1(n_T_427[938]), .A2(n8873), .Y(n8322) );
  AO22X1_LVT U9586 ( .A1(n3970), .A2(n_T_427[427]), .A3(n4021), .A4(
        n_T_427[683]), .Y(n8318) );
  AO22X1_LVT U9587 ( .A1(n3967), .A2(n_T_427[299]), .A3(n4052), .A4(
        n_T_427[43]), .Y(n8317) );
  AO22X1_LVT U9588 ( .A1(n4034), .A2(n_T_427[619]), .A3(n4027), .A4(
        n_T_427[874]), .Y(n8316) );
  AO22X1_LVT U9589 ( .A1(n2837), .A2(n_T_427[107]), .A3(n4037), .A4(
        n_T_427[363]), .Y(n8315) );
  NOR4X1_LVT U9590 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .Y(n8319)
         );
  NAND3X0_LVT U9591 ( .A1(n8321), .A2(n8322), .A3(n8320), .Y(n8329) );
  NAND2X0_LVT U9592 ( .A1(n_T_427[491]), .A2(n9052), .Y(n8325) );
  NAND2X0_LVT U9593 ( .A1(n_T_427[235]), .A2(n3624), .Y(n8324) );
  NAND3X0_LVT U9594 ( .A1(n8326), .A2(n8325), .A3(n8324), .Y(n8327) );
  NAND2X0_LVT U9595 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[43]), .Y(n8333) );
  NAND2X0_LVT U9596 ( .A1(n9065), .A2(n_T_1165[43]), .Y(n8332) );
  NAND2X0_LVT U9597 ( .A1(n2497), .A2(n_T_628[43]), .Y(n8331) );
  NAND2X0_LVT U9598 ( .A1(n9066), .A2(n_T_918[43]), .Y(n8330) );
  NAND4X0_LVT U9599 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .Y(
        io_fpu_fromint_data[43]) );
  NAND2X0_LVT U9600 ( .A1(n3787), .A2(n_T_427[556]), .Y(n8343) );
  NAND2X0_LVT U9601 ( .A1(n2982), .A2(n4439), .Y(n8342) );
  AO22X1_LVT U9602 ( .A1(n3963), .A2(n_T_427[492]), .A3(n4037), .A4(
        n_T_427[364]), .Y(n8339) );
  AO22X1_LVT U9603 ( .A1(n3970), .A2(n_T_427[428]), .A3(n3966), .A4(
        n_T_427[300]), .Y(n8338) );
  AO22X1_LVT U9604 ( .A1(n4024), .A2(n_T_427[939]), .A3(n4020), .A4(
        n_T_427[684]), .Y(n8336) );
  AO22X1_LVT U9605 ( .A1(n3974), .A2(n_T_427[172]), .A3(n4048), .A4(
        n_T_427[747]), .Y(n8335) );
  AO22X1_LVT U9606 ( .A1(n4034), .A2(n_T_427[620]), .A3(n4027), .A4(
        n_T_427[875]), .Y(n8334) );
  OR3X1_LVT U9607 ( .A1(n8336), .A2(n8335), .A3(n8334), .Y(n8337) );
  OR3X1_LVT U9608 ( .A1(n8339), .A2(n8338), .A3(n8337), .Y(n8340) );
  NAND2X0_LVT U9609 ( .A1(n4053), .A2(n8340), .Y(n8341) );
  NAND2X0_LVT U9610 ( .A1(n8944), .A2(n_T_427[44]), .Y(n8345) );
  NAND2X0_LVT U9611 ( .A1(n3745), .A2(n_T_427[236]), .Y(n8344) );
  NAND2X0_LVT U9612 ( .A1(n3635), .A2(n_T_427[1259]), .Y(n8347) );
  NAND2X0_LVT U9613 ( .A1(n3669), .A2(n_T_427[1131]), .Y(n8346) );
  AND2X1_LVT U9614 ( .A1(n8347), .A2(n8346), .Y(n8350) );
  NAND2X0_LVT U9615 ( .A1(n3761), .A2(n_T_427[1003]), .Y(n8349) );
  NAND2X0_LVT U9616 ( .A1(n3716), .A2(n_T_427[1067]), .Y(n8348) );
  NAND2X0_LVT U9617 ( .A1(n3602), .A2(n_T_427[1387]), .Y(n8351) );
  OA21X1_LVT U9618 ( .A1(n3465), .A2(n3988), .A3(n8351), .Y(n8354) );
  NAND2X0_LVT U9619 ( .A1(n3626), .A2(n_T_427[1451]), .Y(n8353) );
  AND3X1_LVT U9620 ( .A1(n8354), .A2(n8353), .A3(n8352), .Y(n8357) );
  NAND2X0_LVT U9621 ( .A1(n3600), .A2(n_T_427[811]), .Y(n8356) );
  NAND2X0_LVT U9622 ( .A1(n3707), .A2(n_T_427[108]), .Y(n8355) );
  NAND2X0_LVT U9623 ( .A1(n3657), .A2(n_T_427[1707]), .Y(n8358) );
  NAND2X0_LVT U9624 ( .A1(n2093), .A2(n_T_427[1323]), .Y(n8360) );
  NAND2X0_LVT U9625 ( .A1(n2092), .A2(n_T_427[1771]), .Y(n8359) );
  NAND2X0_LVT U9626 ( .A1(n3770), .A2(n_T_427[1515]), .Y(n8362) );
  NAND2X0_LVT U9627 ( .A1(n3619), .A2(n_T_427[1579]), .Y(n8364) );
  NAND2X0_LVT U9628 ( .A1(n3648), .A2(n_T_427[1643]), .Y(n8363) );
  NAND2X0_LVT U9629 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[44]), .Y(n8369) );
  NAND2X0_LVT U9630 ( .A1(n9065), .A2(n_T_1165[44]), .Y(n8368) );
  NAND2X0_LVT U9631 ( .A1(n2493), .A2(n_T_628[44]), .Y(n8367) );
  NAND2X0_LVT U9632 ( .A1(n9066), .A2(n_T_918[44]), .Y(n8366) );
  NAND4X0_LVT U9633 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), .Y(
        io_fpu_fromint_data[44]) );
  NAND2X0_LVT U9634 ( .A1(n_T_427[1388]), .A2(n3611), .Y(n8370) );
  OA21X1_LVT U9635 ( .A1(n3151), .A2(n3987), .A3(n8370), .Y(n8373) );
  NAND2X0_LVT U9636 ( .A1(n3628), .A2(n_T_427[1452]), .Y(n8372) );
  NAND2X0_LVT U9637 ( .A1(n2998), .A2(n_T_427[1925]), .Y(n8371) );
  NAND2X0_LVT U9638 ( .A1(n2922), .A2(n_T_427[1708]), .Y(n8374) );
  NAND2X0_LVT U9639 ( .A1(n3997), .A2(n_T_427[1324]), .Y(n8376) );
  NAND2X0_LVT U9640 ( .A1(n4004), .A2(n_T_427[1772]), .Y(n8375) );
  NAND2X0_LVT U9641 ( .A1(n3770), .A2(n_T_427[1516]), .Y(n8378) );
  OA21X1_LVT U9642 ( .A1(n3664), .A2(n3343), .A3(n8378), .Y(n8381) );
  NAND2X0_LVT U9643 ( .A1(n3615), .A2(n_T_427[1580]), .Y(n8380) );
  NAND2X0_LVT U9644 ( .A1(n3651), .A2(n_T_427[1644]), .Y(n8379) );
  NAND2X0_LVT U9645 ( .A1(n3761), .A2(n_T_427[1004]), .Y(n8382) );
  NAND2X0_LVT U9646 ( .A1(n3639), .A2(n_T_427[1260]), .Y(n8384) );
  NAND2X0_LVT U9647 ( .A1(n3671), .A2(n_T_427[1132]), .Y(n8383) );
  NAND2X0_LVT U9648 ( .A1(n8873), .A2(n_T_427[940]), .Y(n8390) );
  AO22X1_LVT U9649 ( .A1(n4021), .A2(n_T_427[685]), .A3(n3960), .A4(
        n_T_427[493]), .Y(n8387) );
  AO22X1_LVT U9650 ( .A1(n3978), .A2(n_T_427[557]), .A3(n4031), .A4(
        n_T_427[621]), .Y(n8386) );
  AO22X1_LVT U9651 ( .A1(n3967), .A2(n_T_427[301]), .A3(n4036), .A4(
        n_T_427[365]), .Y(n8385) );
  NAND3X0_LVT U9652 ( .A1(n8390), .A2(n8388), .A3(n8389), .Y(n8400) );
  NAND2X0_LVT U9653 ( .A1(n3661), .A2(n_T_427[876]), .Y(n8392) );
  NAND2X0_LVT U9654 ( .A1(n3624), .A2(n_T_427[237]), .Y(n8391) );
  NAND2X0_LVT U9655 ( .A1(n8392), .A2(n8391), .Y(n8399) );
  NAND2X0_LVT U9656 ( .A1(n8944), .A2(n_T_427[45]), .Y(n8394) );
  NAND2X0_LVT U9657 ( .A1(n8994), .A2(n_T_427[109]), .Y(n8393) );
  AND2X1_LVT U9658 ( .A1(n8394), .A2(n8393), .Y(n8397) );
  NAND2X0_LVT U9659 ( .A1(n3714), .A2(n_T_427[173]), .Y(n8396) );
  NAND3X0_LVT U9660 ( .A1(n8397), .A2(n8396), .A3(n8395), .Y(n8398) );
  NAND2X0_LVT U9661 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[45]), .Y(n8404) );
  NAND2X0_LVT U9662 ( .A1(n9065), .A2(n_T_1165[45]), .Y(n8403) );
  NAND2X0_LVT U9663 ( .A1(n2493), .A2(n_T_628[45]), .Y(n8402) );
  NAND2X0_LVT U9664 ( .A1(n9066), .A2(n_T_918[45]), .Y(n8401) );
  NAND4X0_LVT U9665 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .Y(
        io_fpu_fromint_data[45]) );
  NAND2X0_LVT U9666 ( .A1(n3610), .A2(n_T_427[1389]), .Y(n8405) );
  OA21X1_LVT U9667 ( .A1(n3466), .A2(n2969), .A3(n8405), .Y(n8408) );
  NAND2X0_LVT U9668 ( .A1(n2966), .A2(n_T_427[1453]), .Y(n8407) );
  NAND2X0_LVT U9669 ( .A1(n3991), .A2(n_T_427[1926]), .Y(n8406) );
  NAND2X0_LVT U9670 ( .A1(n3689), .A2(n_T_427[1709]), .Y(n8409) );
  OA21X1_LVT U9671 ( .A1(n3467), .A2(n3753), .A3(n8409), .Y(n8412) );
  NAND2X0_LVT U9672 ( .A1(n3996), .A2(n_T_427[1325]), .Y(n8411) );
  NAND2X0_LVT U9673 ( .A1(n4005), .A2(n_T_427[1773]), .Y(n8410) );
  NAND2X0_LVT U9674 ( .A1(n3770), .A2(n_T_427[1517]), .Y(n8413) );
  OA21X1_LVT U9675 ( .A1(n4008), .A2(n3345), .A3(n8413), .Y(n8416) );
  NAND2X0_LVT U9676 ( .A1(n3617), .A2(n_T_427[1581]), .Y(n8415) );
  NAND2X0_LVT U9677 ( .A1(n3650), .A2(n_T_427[1645]), .Y(n8414) );
  NAND2X0_LVT U9678 ( .A1(n3760), .A2(n_T_427[1005]), .Y(n8417) );
  NAND2X0_LVT U9679 ( .A1(n3640), .A2(n_T_427[1261]), .Y(n8419) );
  NAND2X0_LVT U9680 ( .A1(n3667), .A2(n_T_427[1133]), .Y(n8418) );
  NAND2X0_LVT U9681 ( .A1(n8939), .A2(n_T_427[366]), .Y(n8427) );
  AO22X1_LVT U9682 ( .A1(n4024), .A2(n_T_427[941]), .A3(n4021), .A4(
        n_T_427[686]), .Y(n8423) );
  AO22X1_LVT U9683 ( .A1(n3974), .A2(n_T_427[174]), .A3(n3966), .A4(
        n_T_427[302]), .Y(n8422) );
  AO22X1_LVT U9684 ( .A1(n3971), .A2(n_T_427[430]), .A3(n4041), .A4(
        n_T_427[110]), .Y(n8421) );
  AO22X1_LVT U9685 ( .A1(n4034), .A2(n_T_427[622]), .A3(n3986), .A4(
        n_T_427[238]), .Y(n8420) );
  NOR4X1_LVT U9686 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .Y(n8424)
         );
  NAND2X0_LVT U9687 ( .A1(n3786), .A2(n_T_427[558]), .Y(n8429) );
  NAND2X0_LVT U9688 ( .A1(n8991), .A2(n_T_427[877]), .Y(n8428) );
  NAND2X0_LVT U9689 ( .A1(n9056), .A2(n_T_427[813]), .Y(n8430) );
  OA21X1_LVT U9690 ( .A1(n3406), .A2(n3691), .A3(n8430), .Y(n8433) );
  NAND2X0_LVT U9691 ( .A1(n_T_427[494]), .A2(n9052), .Y(n8432) );
  NAND2X0_LVT U9692 ( .A1(n8944), .A2(n_T_427[46]), .Y(n8431) );
  NAND2X0_LVT U9693 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[46]), .Y(n8437) );
  NAND2X0_LVT U9694 ( .A1(n9065), .A2(n_T_1165[46]), .Y(n8436) );
  NAND2X0_LVT U9695 ( .A1(n2493), .A2(n_T_628[46]), .Y(n8435) );
  NAND2X0_LVT U9696 ( .A1(n9066), .A2(n_T_918[46]), .Y(n8434) );
  NAND4X0_LVT U9697 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .Y(
        io_fpu_fromint_data[46]) );
  NAND2X0_LVT U9698 ( .A1(n3610), .A2(n_T_427[1390]), .Y(n8438) );
  OA21X1_LVT U9699 ( .A1(n3152), .A2(n3989), .A3(n8438), .Y(n8441) );
  NAND2X0_LVT U9700 ( .A1(n3626), .A2(n_T_427[1454]), .Y(n8440) );
  NAND2X0_LVT U9701 ( .A1(n3992), .A2(n_T_427[1927]), .Y(n8439) );
  NAND2X0_LVT U9702 ( .A1(n3689), .A2(n_T_427[1710]), .Y(n8442) );
  NAND2X0_LVT U9703 ( .A1(n2094), .A2(n_T_427[1326]), .Y(n8444) );
  NAND2X0_LVT U9704 ( .A1(n2091), .A2(n_T_427[1774]), .Y(n8443) );
  NAND2X0_LVT U9705 ( .A1(n3770), .A2(n_T_427[1518]), .Y(n8446) );
  NAND2X0_LVT U9706 ( .A1(n3618), .A2(n_T_427[1582]), .Y(n8448) );
  NAND2X0_LVT U9707 ( .A1(n3642), .A2(n_T_427[1646]), .Y(n8447) );
  NAND2X0_LVT U9708 ( .A1(n3758), .A2(n_T_427[1006]), .Y(n8450) );
  NAND2X0_LVT U9709 ( .A1(n3639), .A2(n_T_427[1262]), .Y(n8452) );
  NAND2X0_LVT U9710 ( .A1(n3675), .A2(n_T_427[1134]), .Y(n8451) );
  NAND2X0_LVT U9711 ( .A1(n2982), .A2(n4448), .Y(n8459) );
  AO22X1_LVT U9712 ( .A1(n4024), .A2(n_T_427[942]), .A3(n4031), .A4(
        n_T_427[623]), .Y(n8456) );
  AO22X1_LVT U9713 ( .A1(n3978), .A2(n_T_427[559]), .A3(n3960), .A4(
        n_T_427[495]), .Y(n8455) );
  AO22X1_LVT U9714 ( .A1(n3971), .A2(n_T_427[431]), .A3(n4036), .A4(
        n_T_427[367]), .Y(n8454) );
  AO22X1_LVT U9715 ( .A1(n4052), .A2(n_T_427[47]), .A3(n4047), .A4(
        n_T_427[750]), .Y(n8453) );
  NOR4X1_LVT U9716 ( .A1(n8456), .A2(n8455), .A3(n8454), .A4(n8453), .Y(n8457)
         );
  NAND2X0_LVT U9717 ( .A1(n3714), .A2(n_T_427[175]), .Y(n8461) );
  NAND2X0_LVT U9718 ( .A1(n8991), .A2(n_T_427[878]), .Y(n8460) );
  NAND2X0_LVT U9719 ( .A1(n_T_427[111]), .A2(n8994), .Y(n8462) );
  OA21X1_LVT U9720 ( .A1(n3482), .A2(n8996), .A3(n8462), .Y(n8465) );
  NAND2X0_LVT U9721 ( .A1(n9056), .A2(n_T_427[814]), .Y(n8464) );
  NAND2X0_LVT U9722 ( .A1(n3624), .A2(n_T_427[239]), .Y(n8463) );
  NAND2X0_LVT U9723 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[47]), .Y(n8469) );
  NAND2X0_LVT U9724 ( .A1(n9065), .A2(n_T_1165[47]), .Y(n8468) );
  NAND2X0_LVT U9725 ( .A1(n2493), .A2(n_T_628[47]), .Y(n8467) );
  NAND2X0_LVT U9726 ( .A1(n9066), .A2(n_T_918[47]), .Y(n8466) );
  NAND4X0_LVT U9727 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), .Y(
        io_fpu_fromint_data[47]) );
  NAND2X0_LVT U9728 ( .A1(n3787), .A2(n_T_427[560]), .Y(n8476) );
  NAND2X0_LVT U9729 ( .A1(n3060), .A2(n4451), .Y(n8475) );
  AO22X1_LVT U9730 ( .A1(n4024), .A2(n_T_427[943]), .A3(n3966), .A4(
        n_T_427[304]), .Y(n8472) );
  AO22X1_LVT U9731 ( .A1(n4038), .A2(n_T_427[368]), .A3(n4048), .A4(
        n_T_427[751]), .Y(n8471) );
  OR3X1_LVT U9732 ( .A1(n8472), .A2(n8471), .A3(n8470), .Y(n8473) );
  NAND2X0_LVT U9733 ( .A1(n4053), .A2(n8473), .Y(n8474) );
  NAND2X0_LVT U9734 ( .A1(n_T_427[496]), .A2(n9052), .Y(n8478) );
  NAND2X0_LVT U9735 ( .A1(n9056), .A2(n_T_427[815]), .Y(n8477) );
  NAND2X0_LVT U9736 ( .A1(n3759), .A2(n_T_427[1007]), .Y(n8480) );
  NAND2X0_LVT U9737 ( .A1(n4014), .A2(n_T_427[1071]), .Y(n8479) );
  NAND2X0_LVT U9738 ( .A1(n3604), .A2(n_T_427[1391]), .Y(n8481) );
  OA21X1_LVT U9739 ( .A1(n3153), .A2(n3987), .A3(n8481), .Y(n8484) );
  NAND2X0_LVT U9740 ( .A1(n2966), .A2(n_T_427[1455]), .Y(n8483) );
  NAND2X0_LVT U9741 ( .A1(n3991), .A2(n_T_427[1928]), .Y(n8482) );
  AND3X1_LVT U9742 ( .A1(n8484), .A2(n8483), .A3(n8482), .Y(n8487) );
  NAND2X0_LVT U9743 ( .A1(n3707), .A2(n_T_427[112]), .Y(n8485) );
  NAND2X0_LVT U9744 ( .A1(n3689), .A2(n_T_427[1711]), .Y(n8488) );
  NAND2X0_LVT U9745 ( .A1(n3997), .A2(n_T_427[1327]), .Y(n8490) );
  NAND2X0_LVT U9746 ( .A1(n2091), .A2(n_T_427[1775]), .Y(n8489) );
  NAND3X0_LVT U9747 ( .A1(n8490), .A2(n8491), .A3(n8489), .Y(n8497) );
  OA21X1_LVT U9748 ( .A1(n4009), .A2(n3348), .A3(n8492), .Y(n8495) );
  NAND2X0_LVT U9749 ( .A1(n3620), .A2(n_T_427[1583]), .Y(n8494) );
  NAND3X0_LVT U9750 ( .A1(n8493), .A2(n8494), .A3(n8495), .Y(n8496) );
  NAND2X0_LVT U9751 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[48]), .Y(n8501) );
  NAND2X0_LVT U9752 ( .A1(n9065), .A2(n_T_1165[48]), .Y(n8500) );
  NAND2X0_LVT U9753 ( .A1(n2497), .A2(n_T_628[48]), .Y(n8499) );
  NAND2X0_LVT U9754 ( .A1(n9066), .A2(n_T_918[48]), .Y(n8498) );
  NAND4X0_LVT U9755 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .Y(
        io_fpu_fromint_data[48]) );
  NAND2X0_LVT U9756 ( .A1(n_T_427[1392]), .A2(n3611), .Y(n8502) );
  OA21X1_LVT U9757 ( .A1(n3154), .A2(n3988), .A3(n8502), .Y(n8505) );
  NAND2X0_LVT U9758 ( .A1(n3626), .A2(n_T_427[1456]), .Y(n8504) );
  NAND2X0_LVT U9759 ( .A1(n2986), .A2(n_T_427[1929]), .Y(n8503) );
  NAND2X0_LVT U9760 ( .A1(n3657), .A2(n_T_427[1712]), .Y(n8506) );
  OA21X1_LVT U9761 ( .A1(n3468), .A2(n3994), .A3(n8506), .Y(n8509) );
  NAND2X0_LVT U9762 ( .A1(n3997), .A2(n_T_427[1328]), .Y(n8508) );
  NAND2X0_LVT U9763 ( .A1(n4004), .A2(n_T_427[1776]), .Y(n8507) );
  NAND2X0_LVT U9764 ( .A1(n3769), .A2(n_T_427[1520]), .Y(n8510) );
  NAND2X0_LVT U9765 ( .A1(n3619), .A2(n_T_427[1584]), .Y(n8512) );
  NAND2X0_LVT U9766 ( .A1(n3648), .A2(n_T_427[1648]), .Y(n8511) );
  NAND2X0_LVT U9767 ( .A1(n3756), .A2(n_T_427[1008]), .Y(n8514) );
  NAND2X0_LVT U9768 ( .A1(n_T_427[1264]), .A2(n3636), .Y(n8516) );
  NAND2X0_LVT U9769 ( .A1(n3673), .A2(n_T_427[1136]), .Y(n8515) );
  NAND2X0_LVT U9770 ( .A1(n8837), .A2(n_T_427[625]), .Y(n8524) );
  NAND2X0_LVT U9771 ( .A1(n2982), .A2(n4454), .Y(n8523) );
  AO22X1_LVT U9772 ( .A1(n4021), .A2(n_T_427[689]), .A3(n3976), .A4(
        n_T_427[561]), .Y(n8520) );
  AO22X1_LVT U9773 ( .A1(n3971), .A2(n_T_427[433]), .A3(n4036), .A4(
        n_T_427[369]), .Y(n8519) );
  AO22X1_LVT U9774 ( .A1(n4023), .A2(n_T_427[944]), .A3(n3986), .A4(
        n_T_427[241]), .Y(n8518) );
  AO22X1_LVT U9775 ( .A1(n3967), .A2(n_T_427[305]), .A3(n4048), .A4(
        n_T_427[752]), .Y(n8517) );
  NOR4X1_LVT U9776 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .Y(n8521)
         );
  NAND2X0_LVT U9777 ( .A1(n_T_427[497]), .A2(n9052), .Y(n8526) );
  NAND2X0_LVT U9778 ( .A1(n_T_427[177]), .A2(n3713), .Y(n8525) );
  NAND2X0_LVT U9779 ( .A1(n8991), .A2(n_T_427[880]), .Y(n8528) );
  NAND2X0_LVT U9780 ( .A1(n9056), .A2(n_T_427[816]), .Y(n8527) );
  AND2X1_LVT U9781 ( .A1(n8528), .A2(n8527), .Y(n8531) );
  NAND2X0_LVT U9782 ( .A1(n8944), .A2(n_T_427[49]), .Y(n8530) );
  NAND2X0_LVT U9783 ( .A1(n8994), .A2(n_T_427[113]), .Y(n8529) );
  NAND2X0_LVT U9784 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[49]), .Y(n8535) );
  NAND2X0_LVT U9785 ( .A1(n9065), .A2(n_T_1165[49]), .Y(n8534) );
  NAND2X0_LVT U9786 ( .A1(n2493), .A2(n_T_628[49]), .Y(n8533) );
  NAND2X0_LVT U9787 ( .A1(n9066), .A2(n_T_918[49]), .Y(n8532) );
  NAND4X0_LVT U9788 ( .A1(n8535), .A2(n8534), .A3(n8533), .A4(n8532), .Y(
        io_fpu_fromint_data[49]) );
  NAND2X0_LVT U9789 ( .A1(n3759), .A2(n_T_427[1009]), .Y(n8536) );
  OA21X1_LVT U9790 ( .A1(n4012), .A2(n3351), .A3(n8536), .Y(n8539) );
  NAND2X0_LVT U9791 ( .A1(n3637), .A2(n_T_427[1265]), .Y(n8538) );
  NAND2X0_LVT U9792 ( .A1(n3670), .A2(n_T_427[1137]), .Y(n8537) );
  NAND2X0_LVT U9793 ( .A1(n3788), .A2(n_T_427[562]), .Y(n8549) );
  NAND2X0_LVT U9794 ( .A1(n2982), .A2(n4457), .Y(n8548) );
  AO22X1_LVT U9795 ( .A1(n3971), .A2(n_T_427[434]), .A3(n3966), .A4(
        n_T_427[306]), .Y(n8545) );
  AO22X1_LVT U9796 ( .A1(n3975), .A2(n_T_427[178]), .A3(n4036), .A4(
        n_T_427[370]), .Y(n8544) );
  AO22X1_LVT U9797 ( .A1(n4023), .A2(n_T_427[945]), .A3(n4031), .A4(
        n_T_427[626]), .Y(n8542) );
  AO22X1_LVT U9798 ( .A1(n4021), .A2(n_T_427[690]), .A3(n4043), .A4(
        n_T_427[114]), .Y(n8541) );
  AO22X1_LVT U9799 ( .A1(n3982), .A2(n_T_427[817]), .A3(n4052), .A4(
        n_T_427[50]), .Y(n8540) );
  OR3X1_LVT U9800 ( .A1(n8542), .A2(n8541), .A3(n8540), .Y(n8543) );
  OR3X1_LVT U9801 ( .A1(n8545), .A2(n8544), .A3(n8543), .Y(n8546) );
  NAND2X0_LVT U9802 ( .A1(n4053), .A2(n8546), .Y(n8547) );
  AND3X1_LVT U9803 ( .A1(n8549), .A2(n8548), .A3(n8547), .Y(n8552) );
  NAND2X0_LVT U9804 ( .A1(n8991), .A2(n_T_427[881]), .Y(n8551) );
  NAND2X0_LVT U9805 ( .A1(n2922), .A2(n_T_427[1713]), .Y(n8553) );
  NAND2X0_LVT U9806 ( .A1(n3996), .A2(n_T_427[1329]), .Y(n8555) );
  NAND2X0_LVT U9807 ( .A1(n4002), .A2(n_T_427[1777]), .Y(n8554) );
  NAND2X0_LVT U9808 ( .A1(n3770), .A2(n_T_427[1521]), .Y(n8557) );
  OA21X1_LVT U9809 ( .A1(n2081), .A2(n3352), .A3(n8557), .Y(n8560) );
  NAND2X0_LVT U9810 ( .A1(n3615), .A2(n_T_427[1585]), .Y(n8559) );
  NAND2X0_LVT U9811 ( .A1(n3650), .A2(n_T_427[1649]), .Y(n8558) );
  NAND2X0_LVT U9812 ( .A1(n_T_427[242]), .A2(n9058), .Y(n8561) );
  NAND2X0_LVT U9813 ( .A1(n3606), .A2(n_T_427[1393]), .Y(n8563) );
  OA21X1_LVT U9814 ( .A1(n3155), .A2(n2969), .A3(n8563), .Y(n8564) );
  NAND2X0_LVT U9815 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[50]), .Y(n8568) );
  NAND2X0_LVT U9816 ( .A1(n9065), .A2(n_T_1165[50]), .Y(n8567) );
  NAND2X0_LVT U9817 ( .A1(n2493), .A2(n_T_628[50]), .Y(n8566) );
  NAND2X0_LVT U9818 ( .A1(n9066), .A2(n_T_918[50]), .Y(n8565) );
  NAND4X0_LVT U9819 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .Y(
        io_fpu_fromint_data[50]) );
  NAND2X0_LVT U9820 ( .A1(n3608), .A2(n_T_427[1394]), .Y(n8569) );
  OA21X1_LVT U9821 ( .A1(n3156), .A2(n3988), .A3(n8569), .Y(n8572) );
  NAND2X0_LVT U9822 ( .A1(n3627), .A2(n_T_427[1458]), .Y(n8571) );
  NAND2X0_LVT U9823 ( .A1(n2985), .A2(n_T_427[1930]), .Y(n8570) );
  AND3X1_LVT U9824 ( .A1(n8572), .A2(n8571), .A3(n8570), .Y(n8575) );
  NAND2X0_LVT U9825 ( .A1(n3661), .A2(n_T_427[882]), .Y(n8574) );
  NAND2X0_LVT U9826 ( .A1(n3647), .A2(n_T_427[51]), .Y(n8573) );
  NAND2X0_LVT U9827 ( .A1(n3788), .A2(n_T_427[563]), .Y(n8586) );
  NAND2X0_LVT U9828 ( .A1(n3060), .A2(n4460), .Y(n8585) );
  AO22X1_LVT U9829 ( .A1(n4022), .A2(n_T_427[691]), .A3(n4036), .A4(
        n_T_427[371]), .Y(n8582) );
  AO22X1_LVT U9830 ( .A1(n4043), .A2(n_T_427[115]), .A3(n4048), .A4(
        n_T_427[754]), .Y(n8581) );
  AOI22X1_LVT U9831 ( .A1(n2859), .A2(n_T_427[179]), .A3(n3979), .A4(
        n_T_427[818]), .Y(n8579) );
  AOI22X1_LVT U9832 ( .A1(n3971), .A2(n_T_427[435]), .A3(n4023), .A4(
        n_T_427[946]), .Y(n8578) );
  NAND2X0_LVT U9833 ( .A1(n4031), .A2(n_T_427[627]), .Y(n8577) );
  NAND2X0_LVT U9834 ( .A1(n3986), .A2(n_T_427[243]), .Y(n8576) );
  NAND4X0_LVT U9835 ( .A1(n8579), .A2(n8578), .A3(n8577), .A4(n8576), .Y(n8580) );
  OR3X1_LVT U9836 ( .A1(n8582), .A2(n8581), .A3(n8580), .Y(n8583) );
  NAND2X0_LVT U9837 ( .A1(n4053), .A2(n8583), .Y(n8584) );
  NAND2X0_LVT U9838 ( .A1(n_T_427[499]), .A2(n9052), .Y(n8588) );
  NAND2X0_LVT U9839 ( .A1(n3789), .A2(n_T_427[307]), .Y(n8587) );
  NAND2X0_LVT U9840 ( .A1(n3641), .A2(n_T_427[1266]), .Y(n8590) );
  NAND2X0_LVT U9841 ( .A1(n3668), .A2(n_T_427[1138]), .Y(n8589) );
  NAND2X0_LVT U9842 ( .A1(n3689), .A2(n_T_427[1714]), .Y(n8591) );
  NAND2X0_LVT U9843 ( .A1(n3996), .A2(n_T_427[1330]), .Y(n8593) );
  NAND2X0_LVT U9844 ( .A1(n4005), .A2(n_T_427[1778]), .Y(n8592) );
  NAND3X0_LVT U9845 ( .A1(n8593), .A2(n8594), .A3(n8592), .Y(n8600) );
  NAND2X0_LVT U9846 ( .A1(n3769), .A2(n_T_427[1522]), .Y(n8595) );
  NAND2X0_LVT U9847 ( .A1(n3620), .A2(n_T_427[1586]), .Y(n8597) );
  NAND3X0_LVT U9848 ( .A1(n8598), .A2(n8597), .A3(n8596), .Y(n8599) );
  NAND2X0_LVT U9849 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[51]), .Y(n8604) );
  NAND2X0_LVT U9850 ( .A1(n9065), .A2(n_T_1165[51]), .Y(n8603) );
  NAND2X0_LVT U9851 ( .A1(n_T_628[51]), .A2(n2497), .Y(n8602) );
  NAND2X0_LVT U9852 ( .A1(n9066), .A2(n_T_918[51]), .Y(n8601) );
  NAND4X0_LVT U9853 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .Y(
        io_fpu_fromint_data[51]) );
  NAND2X0_LVT U9854 ( .A1(n3603), .A2(n_T_427[1395]), .Y(n8605) );
  OA21X1_LVT U9855 ( .A1(n3157), .A2(n3987), .A3(n8605), .Y(n8608) );
  NAND2X0_LVT U9856 ( .A1(n3627), .A2(n_T_427[1459]), .Y(n8607) );
  NAND2X0_LVT U9857 ( .A1(n3991), .A2(n_T_427[1931]), .Y(n8606) );
  NAND2X0_LVT U9858 ( .A1(n2922), .A2(n_T_427[1715]), .Y(n8609) );
  OA21X1_LVT U9859 ( .A1(n3469), .A2(n3994), .A3(n8609), .Y(n8612) );
  NAND2X0_LVT U9860 ( .A1(n3996), .A2(n_T_427[1331]), .Y(n8611) );
  NAND2X0_LVT U9861 ( .A1(n4002), .A2(n_T_427[1779]), .Y(n8610) );
  NAND2X0_LVT U9862 ( .A1(n3770), .A2(n_T_427[1523]), .Y(n8613) );
  OA21X1_LVT U9863 ( .A1(n4010), .A2(n3355), .A3(n8613), .Y(n8616) );
  NAND2X0_LVT U9864 ( .A1(n3617), .A2(n_T_427[1587]), .Y(n8615) );
  NAND2X0_LVT U9865 ( .A1(n3652), .A2(n_T_427[1651]), .Y(n8614) );
  NAND2X0_LVT U9866 ( .A1(n3761), .A2(n_T_427[1011]), .Y(n8617) );
  NAND2X0_LVT U9867 ( .A1(n3641), .A2(n_T_427[1267]), .Y(n8619) );
  NAND2X0_LVT U9868 ( .A1(n3673), .A2(n_T_427[1139]), .Y(n8618) );
  NAND2X0_LVT U9869 ( .A1(n3786), .A2(n_T_427[564]), .Y(n8627) );
  NAND2X0_LVT U9870 ( .A1(n3060), .A2(n4463), .Y(n8626) );
  AO22X1_LVT U9871 ( .A1(n4022), .A2(n_T_427[692]), .A3(n4036), .A4(
        n_T_427[372]), .Y(n8623) );
  AO22X1_LVT U9872 ( .A1(n4023), .A2(n_T_427[947]), .A3(n3986), .A4(
        n_T_427[244]), .Y(n8622) );
  AO22X1_LVT U9873 ( .A1(n4034), .A2(n_T_427[628]), .A3(n4027), .A4(
        n_T_427[883]), .Y(n8621) );
  AO22X1_LVT U9874 ( .A1(n3982), .A2(n_T_427[819]), .A3(n4052), .A4(
        n_T_427[52]), .Y(n8620) );
  NOR4X1_LVT U9875 ( .A1(n8623), .A2(n8622), .A3(n8621), .A4(n8620), .Y(n8624)
         );
  NAND2X0_LVT U9876 ( .A1(n_T_427[500]), .A2(n9052), .Y(n8629) );
  NAND2X0_LVT U9877 ( .A1(n3789), .A2(n_T_427[308]), .Y(n8628) );
  NAND2X0_LVT U9878 ( .A1(n_T_427[180]), .A2(n3791), .Y(n8630) );
  OA21X1_LVT U9879 ( .A1(n3408), .A2(n3691), .A3(n8630), .Y(n8632) );
  NAND2X0_LVT U9880 ( .A1(n_T_427[116]), .A2(n8994), .Y(n8631) );
  NAND2X0_LVT U9881 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[52]), .Y(n8636) );
  NAND2X0_LVT U9882 ( .A1(n9065), .A2(n_T_1165[52]), .Y(n8635) );
  NAND2X0_LVT U9883 ( .A1(n2497), .A2(n_T_628[52]), .Y(n8634) );
  NAND2X0_LVT U9884 ( .A1(n9066), .A2(n_T_918[52]), .Y(n8633) );
  NAND4X0_LVT U9885 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .Y(
        io_fpu_fromint_data[52]) );
  NAND2X0_LVT U9886 ( .A1(n3607), .A2(n_T_427[1396]), .Y(n8637) );
  OA21X1_LVT U9887 ( .A1(n3158), .A2(n3989), .A3(n8637), .Y(n8640) );
  NAND2X0_LVT U9888 ( .A1(n3627), .A2(n_T_427[1460]), .Y(n8639) );
  NAND2X0_LVT U9889 ( .A1(n3991), .A2(n_T_427[1932]), .Y(n8638) );
  AND3X1_LVT U9890 ( .A1(n8638), .A2(n8639), .A3(n8640), .Y(n8643) );
  NAND2X0_LVT U9891 ( .A1(n3647), .A2(n_T_427[53]), .Y(n8642) );
  NAND2X0_LVT U9892 ( .A1(n3786), .A2(n_T_427[565]), .Y(n8654) );
  NAND2X0_LVT U9893 ( .A1(n3665), .A2(n4466), .Y(n8653) );
  AO22X1_LVT U9894 ( .A1(n3963), .A2(n_T_427[501]), .A3(n4036), .A4(
        n_T_427[373]), .Y(n8650) );
  AO22X1_LVT U9895 ( .A1(n4042), .A2(n_T_427[117]), .A3(n4048), .A4(
        n_T_427[756]), .Y(n8649) );
  AOI22X1_LVT U9896 ( .A1(n3974), .A2(n_T_427[181]), .A3(n3979), .A4(
        n_T_427[820]), .Y(n8647) );
  AOI22X1_LVT U9897 ( .A1(n4023), .A2(n_T_427[948]), .A3(n4018), .A4(
        n_T_427[693]), .Y(n8646) );
  NAND2X0_LVT U9898 ( .A1(n4031), .A2(n_T_427[629]), .Y(n8645) );
  NAND2X0_LVT U9899 ( .A1(n3986), .A2(n_T_427[245]), .Y(n8644) );
  NAND4X0_LVT U9900 ( .A1(n8647), .A2(n8646), .A3(n8645), .A4(n8644), .Y(n8648) );
  OR3X1_LVT U9901 ( .A1(n8650), .A2(n8649), .A3(n8648), .Y(n8651) );
  NAND2X0_LVT U9902 ( .A1(n4053), .A2(n8651), .Y(n8652) );
  NAND2X0_LVT U9903 ( .A1(n8991), .A2(n_T_427[884]), .Y(n8656) );
  NAND2X0_LVT U9904 ( .A1(n3789), .A2(n_T_427[309]), .Y(n8655) );
  NAND2X0_LVT U9905 ( .A1(n3755), .A2(n_T_427[1012]), .Y(n8657) );
  OA21X1_LVT U9906 ( .A1(n4013), .A2(n3357), .A3(n8657), .Y(n8660) );
  NAND2X0_LVT U9907 ( .A1(n3637), .A2(n_T_427[1268]), .Y(n8659) );
  NAND2X0_LVT U9908 ( .A1(n3667), .A2(n_T_427[1140]), .Y(n8658) );
  NAND2X0_LVT U9909 ( .A1(n3689), .A2(n_T_427[1716]), .Y(n8661) );
  OA21X1_LVT U9910 ( .A1(n3470), .A2(n3601), .A3(n8661), .Y(n8664) );
  NAND2X0_LVT U9911 ( .A1(n2094), .A2(n_T_427[1332]), .Y(n8663) );
  NAND2X0_LVT U9912 ( .A1(n4002), .A2(n_T_427[1780]), .Y(n8662) );
  NAND3X0_LVT U9913 ( .A1(n8663), .A2(n8664), .A3(n8662), .Y(n8670) );
  NAND2X0_LVT U9914 ( .A1(n3770), .A2(n_T_427[1524]), .Y(n8665) );
  OA21X1_LVT U9915 ( .A1(n3663), .A2(n3358), .A3(n8665), .Y(n8668) );
  NAND2X0_LVT U9916 ( .A1(n3615), .A2(n_T_427[1588]), .Y(n8667) );
  NAND2X0_LVT U9917 ( .A1(n3650), .A2(n_T_427[1652]), .Y(n8666) );
  NAND3X0_LVT U9918 ( .A1(n8668), .A2(n8667), .A3(n8666), .Y(n8669) );
  NAND2X0_LVT U9919 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[53]), .Y(n8674) );
  NAND2X0_LVT U9920 ( .A1(n9065), .A2(n_T_1165[53]), .Y(n8673) );
  NAND2X0_LVT U9921 ( .A1(n_T_628[53]), .A2(n2493), .Y(n8672) );
  NAND2X0_LVT U9922 ( .A1(n9066), .A2(n_T_918[53]), .Y(n8671) );
  NAND4X0_LVT U9923 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .Y(
        io_fpu_fromint_data[53]) );
  NAND2X0_LVT U9924 ( .A1(n3607), .A2(n_T_427[1397]), .Y(n8675) );
  NAND2X0_LVT U9925 ( .A1(n3627), .A2(n_T_427[1461]), .Y(n8677) );
  NAND2X0_LVT U9926 ( .A1(n2882), .A2(n_T_427[1933]), .Y(n8676) );
  AND3X1_LVT U9927 ( .A1(n8678), .A2(n8677), .A3(n8676), .Y(n8681) );
  NAND2X0_LVT U9928 ( .A1(n3647), .A2(n_T_427[54]), .Y(n8680) );
  NAND2X0_LVT U9929 ( .A1(n3789), .A2(n_T_427[310]), .Y(n8692) );
  NAND2X0_LVT U9930 ( .A1(n2982), .A2(n4469), .Y(n8691) );
  AO22X1_LVT U9931 ( .A1(n3976), .A2(n_T_427[566]), .A3(n4042), .A4(
        n_T_427[118]), .Y(n8688) );
  AO22X1_LVT U9932 ( .A1(n4022), .A2(n_T_427[694]), .A3(n4036), .A4(
        n_T_427[374]), .Y(n8687) );
  AOI22X1_LVT U9933 ( .A1(n4023), .A2(n_T_427[949]), .A3(n3960), .A4(
        n_T_427[502]), .Y(n8685) );
  AOI22X1_LVT U9934 ( .A1(n3975), .A2(n_T_427[182]), .A3(n3979), .A4(
        n_T_427[821]), .Y(n8684) );
  NAND2X0_LVT U9935 ( .A1(n4031), .A2(n_T_427[630]), .Y(n8683) );
  NAND2X0_LVT U9936 ( .A1(n4030), .A2(n_T_427[885]), .Y(n8682) );
  NAND4X0_LVT U9937 ( .A1(n8685), .A2(n8684), .A3(n8683), .A4(n8682), .Y(n8686) );
  OR3X1_LVT U9938 ( .A1(n8688), .A2(n8687), .A3(n8686), .Y(n8689) );
  NAND2X0_LVT U9939 ( .A1(n4053), .A2(n8689), .Y(n8690) );
  NAND2X0_LVT U9940 ( .A1(n3712), .A2(n_T_427[1013]), .Y(n8693) );
  OA21X1_LVT U9941 ( .A1(n4012), .A2(n3359), .A3(n8693), .Y(n8696) );
  NAND2X0_LVT U9942 ( .A1(n3636), .A2(n_T_427[1269]), .Y(n8695) );
  NAND2X0_LVT U9943 ( .A1(n3668), .A2(n_T_427[1141]), .Y(n8694) );
  OA21X1_LVT U9944 ( .A1(n3471), .A2(n3601), .A3(n8697), .Y(n8700) );
  NAND2X0_LVT U9945 ( .A1(n3999), .A2(n_T_427[1333]), .Y(n8699) );
  NAND2X0_LVT U9946 ( .A1(n4004), .A2(n_T_427[1781]), .Y(n8698) );
  NAND3X0_LVT U9947 ( .A1(n8700), .A2(n8699), .A3(n8698), .Y(n8706) );
  NAND2X0_LVT U9948 ( .A1(n3770), .A2(n_T_427[1525]), .Y(n8701) );
  OA21X1_LVT U9949 ( .A1(n4009), .A2(n3360), .A3(n8701), .Y(n8704) );
  NAND2X0_LVT U9950 ( .A1(n3616), .A2(n_T_427[1589]), .Y(n8703) );
  NAND2X0_LVT U9951 ( .A1(n_T_427[1653]), .A2(n3651), .Y(n8702) );
  NAND3X0_LVT U9952 ( .A1(n8704), .A2(n8703), .A3(n8702), .Y(n8705) );
  NAND2X0_LVT U9953 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[54]), .Y(n8710) );
  NAND2X0_LVT U9954 ( .A1(n9065), .A2(n_T_1165[54]), .Y(n8709) );
  NAND2X0_LVT U9955 ( .A1(n2493), .A2(n_T_628[54]), .Y(n8708) );
  NAND2X0_LVT U9956 ( .A1(n9066), .A2(n_T_918[54]), .Y(n8707) );
  NAND4X0_LVT U9957 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .Y(
        io_fpu_fromint_data[54]) );
  NAND2X0_LVT U9958 ( .A1(n_T_427[503]), .A2(n9052), .Y(n8711) );
  OA21X1_LVT U9959 ( .A1(n3691), .A2(n3301), .A3(n8711), .Y(n8720) );
  AO22X1_LVT U9960 ( .A1(n4024), .A2(n_T_427[950]), .A3(n3976), .A4(
        n_T_427[567]), .Y(n8715) );
  AO22X1_LVT U9961 ( .A1(n3971), .A2(n_T_427[439]), .A3(n4021), .A4(
        n_T_427[695]), .Y(n8714) );
  AO22X1_LVT U9962 ( .A1(n3967), .A2(n_T_427[311]), .A3(n3979), .A4(
        n_T_427[822]), .Y(n8713) );
  AO22X1_LVT U9963 ( .A1(n4034), .A2(n_T_427[631]), .A3(n4027), .A4(
        n_T_427[886]), .Y(n8712) );
  NOR4X1_LVT U9964 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .Y(n8717)
         );
  NAND2X0_LVT U9965 ( .A1(n2982), .A2(n4472), .Y(n8716) );
  OA21X1_LVT U9966 ( .A1(n8717), .A2(n3612), .A3(n8716), .Y(n8719) );
  NAND2X0_LVT U9967 ( .A1(n8939), .A2(n_T_427[375]), .Y(n8718) );
  NAND2X0_LVT U9968 ( .A1(n3624), .A2(n_T_427[247]), .Y(n8722) );
  NAND2X0_LVT U9969 ( .A1(n8994), .A2(n_T_427[119]), .Y(n8721) );
  AND2X1_LVT U9970 ( .A1(n8722), .A2(n8721), .Y(n8725) );
  NAND2X0_LVT U9971 ( .A1(n_T_427[183]), .A2(n3714), .Y(n8724) );
  NAND2X0_LVT U9972 ( .A1(n3647), .A2(n_T_427[55]), .Y(n8723) );
  NAND2X0_LVT U9973 ( .A1(n3608), .A2(n_T_427[1398]), .Y(n8726) );
  OA21X1_LVT U9974 ( .A1(n3160), .A2(n2969), .A3(n8726), .Y(n8729) );
  NAND2X0_LVT U9975 ( .A1(n2967), .A2(n_T_427[1462]), .Y(n8728) );
  NAND2X0_LVT U9976 ( .A1(n2986), .A2(n_T_427[1934]), .Y(n8727) );
  NAND2X0_LVT U9977 ( .A1(n3657), .A2(n_T_427[1718]), .Y(n8730) );
  OA21X1_LVT U9978 ( .A1(n3161), .A2(n3751), .A3(n8730), .Y(n8733) );
  NAND2X0_LVT U9979 ( .A1(n2094), .A2(n_T_427[1334]), .Y(n8732) );
  NAND2X0_LVT U9980 ( .A1(n4001), .A2(n_T_427[1782]), .Y(n8731) );
  NAND2X0_LVT U9981 ( .A1(n3769), .A2(n_T_427[1526]), .Y(n8734) );
  OA21X1_LVT U9982 ( .A1(n4009), .A2(n3361), .A3(n8734), .Y(n8737) );
  NAND2X0_LVT U9983 ( .A1(n3616), .A2(n_T_427[1590]), .Y(n8736) );
  NAND2X0_LVT U9984 ( .A1(n3643), .A2(n_T_427[1654]), .Y(n8735) );
  NAND2X0_LVT U9985 ( .A1(n_T_427[1270]), .A2(n3636), .Y(n8739) );
  NAND2X0_LVT U9986 ( .A1(n3669), .A2(n_T_427[1142]), .Y(n8738) );
  NAND2X0_LVT U9987 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[55]), .Y(n8744) );
  NAND2X0_LVT U9988 ( .A1(n9065), .A2(n_T_1165[55]), .Y(n8743) );
  NAND2X0_LVT U9989 ( .A1(n2493), .A2(n_T_628[55]), .Y(n8742) );
  NAND2X0_LVT U9990 ( .A1(n9066), .A2(n_T_918[55]), .Y(n8741) );
  NAND4X0_LVT U9991 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .Y(
        io_fpu_fromint_data[55]) );
  AO22X1_LVT U9992 ( .A1(n4022), .A2(n_T_427[696]), .A3(n4036), .A4(
        n_T_427[376]), .Y(n8750) );
  AO22X1_LVT U9993 ( .A1(n4044), .A2(n_T_427[120]), .A3(n4048), .A4(
        n_T_427[759]), .Y(n8749) );
  AO22X1_LVT U9994 ( .A1(n3975), .A2(n_T_427[184]), .A3(n3979), .A4(
        n_T_427[823]), .Y(n8747) );
  AO22X1_LVT U9995 ( .A1(n4023), .A2(n_T_427[951]), .A3(n4031), .A4(
        n_T_427[632]), .Y(n8746) );
  AO22X1_LVT U9996 ( .A1(n3971), .A2(n_T_427[440]), .A3(n3976), .A4(
        n_T_427[568]), .Y(n8745) );
  OR3X1_LVT U9997 ( .A1(n8747), .A2(n8746), .A3(n8745), .Y(n8748) );
  OR3X1_LVT U9998 ( .A1(n8750), .A2(n8749), .A3(n8748), .Y(n8751) );
  NAND2X0_LVT U9999 ( .A1(n4053), .A2(n8751), .Y(n8752) );
  NAND2X0_LVT U10000 ( .A1(n3661), .A2(n_T_427[887]), .Y(n8755) );
  NAND2X0_LVT U10001 ( .A1(n_T_427[504]), .A2(n9052), .Y(n8754) );
  NAND2X0_LVT U10002 ( .A1(n3675), .A2(n_T_427[1143]), .Y(n8756) );
  NAND2X0_LVT U10003 ( .A1(n3758), .A2(n_T_427[1015]), .Y(n8758) );
  NAND2X0_LVT U10004 ( .A1(n3716), .A2(n_T_427[1079]), .Y(n8757) );
  NAND2X0_LVT U10005 ( .A1(n_T_427[1399]), .A2(n3609), .Y(n8759) );
  OA21X1_LVT U10006 ( .A1(n3162), .A2(n3989), .A3(n8759), .Y(n8762) );
  NAND2X0_LVT U10007 ( .A1(n3627), .A2(n_T_427[1463]), .Y(n8761) );
  NAND2X0_LVT U10008 ( .A1(n2998), .A2(n_T_427[1935]), .Y(n8760) );
  AND3X1_LVT U10009 ( .A1(n8762), .A2(n8761), .A3(n8760), .Y(n8765) );
  NAND2X0_LVT U10010 ( .A1(n3745), .A2(n_T_427[248]), .Y(n8764) );
  NAND2X0_LVT U10011 ( .A1(n3647), .A2(n_T_427[56]), .Y(n8763) );
  NAND3X0_LVT U10012 ( .A1(n8765), .A2(n8764), .A3(n8763), .Y(n8775) );
  NAND2X0_LVT U10013 ( .A1(n3689), .A2(n_T_427[1719]), .Y(n8766) );
  OA21X1_LVT U10014 ( .A1(n3472), .A2(n3994), .A3(n8766), .Y(n8769) );
  NAND2X0_LVT U10015 ( .A1(n3999), .A2(n_T_427[1335]), .Y(n8768) );
  NAND2X0_LVT U10016 ( .A1(n4004), .A2(n_T_427[1783]), .Y(n8767) );
  NAND2X0_LVT U10017 ( .A1(n3770), .A2(n_T_427[1527]), .Y(n8770) );
  OA21X1_LVT U10018 ( .A1(n3664), .A2(n3362), .A3(n8770), .Y(n8773) );
  NAND2X0_LVT U10019 ( .A1(n3617), .A2(n_T_427[1591]), .Y(n8772) );
  NAND2X0_LVT U10020 ( .A1(n3642), .A2(n_T_427[1655]), .Y(n8771) );
  OR3X1_LVT U10021 ( .A1(n8776), .A2(n8775), .A3(n8774), .Y(N736) );
  NAND2X0_LVT U10022 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[56]), .Y(n8780)
         );
  NAND2X0_LVT U10023 ( .A1(n9065), .A2(n_T_1165[56]), .Y(n8779) );
  NAND2X0_LVT U10024 ( .A1(n2497), .A2(n_T_628[56]), .Y(n8778) );
  NAND2X0_LVT U10025 ( .A1(n9066), .A2(n_T_918[56]), .Y(n8777) );
  NAND4X0_LVT U10026 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .Y(
        io_fpu_fromint_data[56]) );
  NAND2X0_LVT U10027 ( .A1(n3629), .A2(n_T_427[1464]), .Y(n8783) );
  NAND2X0_LVT U10028 ( .A1(n3992), .A2(n_T_427[1936]), .Y(n8782) );
  NAND3X0_LVT U10029 ( .A1(n8784), .A2(n8783), .A3(n8782), .Y(n8790) );
  NAND2X0_LVT U10030 ( .A1(n3689), .A2(n_T_427[1720]), .Y(n8785) );
  OA21X1_LVT U10031 ( .A1(n3751), .A2(n3473), .A3(n8785), .Y(n8788) );
  NAND2X0_LVT U10032 ( .A1(n3997), .A2(n_T_427[1336]), .Y(n8787) );
  NAND2X0_LVT U10033 ( .A1(n4005), .A2(n_T_427[1784]), .Y(n8786) );
  NAND3X0_LVT U10034 ( .A1(n8788), .A2(n8787), .A3(n8786), .Y(n8789) );
  NAND2X0_LVT U10035 ( .A1(n3770), .A2(n_T_427[1528]), .Y(n8791) );
  OA21X1_LVT U10036 ( .A1(n4009), .A2(n3363), .A3(n8791), .Y(n8794) );
  NAND2X0_LVT U10037 ( .A1(n3616), .A2(n_T_427[1592]), .Y(n8793) );
  NAND2X0_LVT U10038 ( .A1(n3649), .A2(n_T_427[1656]), .Y(n8792) );
  NAND3X0_LVT U10039 ( .A1(n8794), .A2(n8793), .A3(n8792), .Y(n8798) );
  NAND2X0_LVT U10040 ( .A1(n_T_427[1272]), .A2(n3638), .Y(n8796) );
  NAND2X0_LVT U10041 ( .A1(n3674), .A2(n_T_427[1144]), .Y(n8795) );
  NAND2X0_LVT U10042 ( .A1(n3787), .A2(n_T_427[569]), .Y(n8806) );
  NAND2X0_LVT U10043 ( .A1(n3665), .A2(n4478), .Y(n8805) );
  AO22X1_LVT U10044 ( .A1(n4023), .A2(n_T_427[952]), .A3(n3960), .A4(
        n_T_427[505]), .Y(n8802) );
  AO22X1_LVT U10045 ( .A1(n4022), .A2(n_T_427[697]), .A3(n4043), .A4(
        n_T_427[121]), .Y(n8801) );
  AO22X1_LVT U10046 ( .A1(n4035), .A2(n_T_427[633]), .A3(n4027), .A4(
        n_T_427[888]), .Y(n8800) );
  AO22X1_LVT U10047 ( .A1(n4039), .A2(n_T_427[377]), .A3(n4052), .A4(
        n_T_427[57]), .Y(n8799) );
  NOR4X1_LVT U10048 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .Y(n8803) );
  NAND3X0_LVT U10049 ( .A1(n8806), .A2(n8805), .A3(n8804), .Y(n8815) );
  NAND2X0_LVT U10050 ( .A1(n3713), .A2(n_T_427[185]), .Y(n8808) );
  NAND2X0_LVT U10051 ( .A1(n3790), .A2(n_T_427[313]), .Y(n8807) );
  NAND2X0_LVT U10052 ( .A1(n8808), .A2(n8807), .Y(n8814) );
  NAND2X0_LVT U10053 ( .A1(n9058), .A2(n_T_427[249]), .Y(n8809) );
  OA21X1_LVT U10054 ( .A1(n3708), .A2(n3302), .A3(n8809), .Y(n8812) );
  NAND2X0_LVT U10055 ( .A1(n9056), .A2(n_T_427[824]), .Y(n8810) );
  NAND3X0_LVT U10056 ( .A1(n8811), .A2(n8812), .A3(n8810), .Y(n8813) );
  NAND2X0_LVT U10057 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[57]), .Y(n8819)
         );
  NAND2X0_LVT U10058 ( .A1(n9065), .A2(n_T_1165[57]), .Y(n8818) );
  NAND2X0_LVT U10059 ( .A1(n2497), .A2(n_T_628[57]), .Y(n8817) );
  NAND2X0_LVT U10060 ( .A1(n9066), .A2(n_T_918[57]), .Y(n8816) );
  NAND4X0_LVT U10061 ( .A1(n8819), .A2(n8818), .A3(n8817), .A4(n8816), .Y(
        io_fpu_fromint_data[57]) );
  NAND2X0_LVT U10062 ( .A1(n3610), .A2(n_T_427[1401]), .Y(n8820) );
  OA21X1_LVT U10063 ( .A1(n3164), .A2(n2969), .A3(n8820), .Y(n8823) );
  NAND2X0_LVT U10064 ( .A1(n3630), .A2(n_T_427[1465]), .Y(n8822) );
  NAND2X0_LVT U10065 ( .A1(n2882), .A2(n_T_427[1937]), .Y(n8821) );
  NAND2X0_LVT U10066 ( .A1(n3689), .A2(n_T_427[1721]), .Y(n8824) );
  OA21X1_LVT U10067 ( .A1(n3474), .A2(n3994), .A3(n8824), .Y(n8827) );
  NAND2X0_LVT U10068 ( .A1(n3999), .A2(n_T_427[1337]), .Y(n8826) );
  NAND2X0_LVT U10069 ( .A1(n4001), .A2(n_T_427[1785]), .Y(n8825) );
  NAND2X0_LVT U10070 ( .A1(n3769), .A2(n_T_427[1529]), .Y(n8828) );
  NAND2X0_LVT U10071 ( .A1(n3619), .A2(n_T_427[1593]), .Y(n8830) );
  NAND3X0_LVT U10072 ( .A1(n8831), .A2(n8830), .A3(n8829), .Y(n8836) );
  NAND2X0_LVT U10073 ( .A1(n3759), .A2(n_T_427[1017]), .Y(n8832) );
  NAND2X0_LVT U10074 ( .A1(n_T_427[1273]), .A2(n3640), .Y(n8834) );
  NAND2X0_LVT U10075 ( .A1(n3675), .A2(n_T_427[1145]), .Y(n8833) );
  NAND2X0_LVT U10076 ( .A1(n8837), .A2(n_T_427[634]), .Y(n8845) );
  NAND2X0_LVT U10077 ( .A1(n3060), .A2(n4481), .Y(n8844) );
  AO22X1_LVT U10078 ( .A1(n4023), .A2(n_T_427[953]), .A3(n4021), .A4(
        n_T_427[698]), .Y(n8841) );
  AO22X1_LVT U10079 ( .A1(n3971), .A2(n_T_427[442]), .A3(n4036), .A4(
        n_T_427[378]), .Y(n8840) );
  AO22X1_LVT U10080 ( .A1(n3986), .A2(n_T_427[250]), .A3(n4028), .A4(
        n_T_427[889]), .Y(n8839) );
  AO22X1_LVT U10081 ( .A1(n4052), .A2(n_T_427[58]), .A3(n4048), .A4(
        n_T_427[761]), .Y(n8838) );
  NOR4X1_LVT U10082 ( .A1(n8841), .A2(n8840), .A3(n8839), .A4(n8838), .Y(n8842) );
  NAND3X0_LVT U10083 ( .A1(n8845), .A2(n8844), .A3(n8843), .Y(n8851) );
  NAND2X0_LVT U10084 ( .A1(n3788), .A2(n_T_427[570]), .Y(n8847) );
  NAND2X0_LVT U10085 ( .A1(n_T_427[506]), .A2(n9052), .Y(n8846) );
  NAND2X0_LVT U10086 ( .A1(n8847), .A2(n8846), .Y(n8850) );
  NAND2X0_LVT U10087 ( .A1(n_T_427[314]), .A2(n9053), .Y(n8848) );
  NAND2X0_LVT U10088 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[58]), .Y(n8855)
         );
  NAND2X0_LVT U10089 ( .A1(n9065), .A2(n_T_1165[58]), .Y(n8854) );
  NAND2X0_LVT U10090 ( .A1(n2497), .A2(n_T_628[58]), .Y(n8853) );
  NAND2X0_LVT U10091 ( .A1(n9066), .A2(n_T_918[58]), .Y(n8852) );
  NAND4X0_LVT U10092 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .Y(
        io_fpu_fromint_data[58]) );
  NAND2X0_LVT U10093 ( .A1(n3609), .A2(n_T_427[1402]), .Y(n8856) );
  OA21X1_LVT U10094 ( .A1(n3165), .A2(n3988), .A3(n8856), .Y(n8859) );
  NAND2X0_LVT U10095 ( .A1(n3628), .A2(n_T_427[1466]), .Y(n8858) );
  NAND2X0_LVT U10096 ( .A1(n2998), .A2(n_T_427[1938]), .Y(n8857) );
  NAND2X0_LVT U10097 ( .A1(n3689), .A2(n_T_427[1722]), .Y(n8860) );
  OA21X1_LVT U10098 ( .A1(n3166), .A2(n3994), .A3(n8860), .Y(n8863) );
  NAND2X0_LVT U10099 ( .A1(n4000), .A2(n_T_427[1338]), .Y(n8862) );
  NAND2X0_LVT U10100 ( .A1(n2092), .A2(n_T_427[1786]), .Y(n8861) );
  NAND2X0_LVT U10101 ( .A1(n3769), .A2(n_T_427[1530]), .Y(n8864) );
  OA21X1_LVT U10102 ( .A1(n3663), .A2(n3367), .A3(n8864), .Y(n8867) );
  NAND2X0_LVT U10103 ( .A1(n3617), .A2(n_T_427[1594]), .Y(n8866) );
  NAND2X0_LVT U10104 ( .A1(n3643), .A2(n_T_427[1658]), .Y(n8865) );
  NAND3X0_LVT U10105 ( .A1(n8867), .A2(n8866), .A3(n8865), .Y(n8872) );
  NAND2X0_LVT U10106 ( .A1(n3757), .A2(n_T_427[1018]), .Y(n8868) );
  NAND2X0_LVT U10107 ( .A1(n3637), .A2(n_T_427[1274]), .Y(n8870) );
  NAND2X0_LVT U10108 ( .A1(n_T_427[1146]), .A2(n3669), .Y(n8869) );
  NAND2X0_LVT U10109 ( .A1(n8873), .A2(n_T_427[954]), .Y(n8881) );
  NAND2X0_LVT U10110 ( .A1(n3060), .A2(n4484), .Y(n8880) );
  AO22X1_LVT U10111 ( .A1(n3971), .A2(n_T_427[443]), .A3(n4021), .A4(
        n_T_427[699]), .Y(n8877) );
  AO22X1_LVT U10112 ( .A1(n2858), .A2(n_T_427[187]), .A3(n4048), .A4(
        n_T_427[762]), .Y(n8876) );
  AO22X1_LVT U10113 ( .A1(n3963), .A2(n_T_427[507]), .A3(n4031), .A4(
        n_T_427[635]), .Y(n8875) );
  AO22X1_LVT U10114 ( .A1(n4041), .A2(n_T_427[123]), .A3(n4036), .A4(
        n_T_427[379]), .Y(n8874) );
  NOR4X1_LVT U10115 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .Y(n8878) );
  NAND3X0_LVT U10116 ( .A1(n8881), .A2(n8880), .A3(n8879), .Y(n8889) );
  NAND2X0_LVT U10117 ( .A1(n3787), .A2(n_T_427[571]), .Y(n8883) );
  NAND2X0_LVT U10118 ( .A1(n3661), .A2(n_T_427[890]), .Y(n8882) );
  NAND2X0_LVT U10119 ( .A1(n8883), .A2(n8882), .Y(n8888) );
  NAND2X0_LVT U10120 ( .A1(n_T_427[251]), .A2(n9058), .Y(n8885) );
  AND2X1_LVT U10121 ( .A1(n8885), .A2(n8884), .Y(n8887) );
  NAND2X0_LVT U10122 ( .A1(n_T_427[315]), .A2(n3790), .Y(n8886) );
  NAND2X0_LVT U10123 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[59]), .Y(n8893)
         );
  NAND2X0_LVT U10124 ( .A1(n9065), .A2(n_T_1165[59]), .Y(n8892) );
  NAND2X0_LVT U10125 ( .A1(n2497), .A2(n_T_628[59]), .Y(n8891) );
  NAND2X0_LVT U10126 ( .A1(n9066), .A2(n_T_918[59]), .Y(n8890) );
  NAND4X0_LVT U10127 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .Y(
        io_fpu_fromint_data[59]) );
  NAND2X0_LVT U10128 ( .A1(n3610), .A2(n_T_427[1403]), .Y(n8894) );
  NAND2X0_LVT U10129 ( .A1(n3628), .A2(n_T_427[1467]), .Y(n8896) );
  NAND2X0_LVT U10130 ( .A1(n2882), .A2(n_T_427[1939]), .Y(n8895) );
  NAND2X0_LVT U10131 ( .A1(n3600), .A2(n_T_427[827]), .Y(n8898) );
  NAND2X0_LVT U10132 ( .A1(n3707), .A2(n_T_427[124]), .Y(n8897) );
  NAND3X0_LVT U10133 ( .A1(n8899), .A2(n8898), .A3(n8897), .Y(n8925) );
  NAND2X0_LVT U10134 ( .A1(n3786), .A2(n_T_427[572]), .Y(n8908) );
  NAND2X0_LVT U10135 ( .A1(n3060), .A2(n4487), .Y(n8907) );
  AO22X1_LVT U10136 ( .A1(n3960), .A2(n_T_427[508]), .A3(n4036), .A4(
        n_T_427[380]), .Y(n8904) );
  AO22X1_LVT U10137 ( .A1(n3970), .A2(n_T_427[444]), .A3(n3964), .A4(
        n_T_427[316]), .Y(n8903) );
  OR3X1_LVT U10138 ( .A1(n8904), .A2(n8903), .A3(n8902), .Y(n8905) );
  NAND2X0_LVT U10139 ( .A1(n4053), .A2(n8905), .Y(n8906) );
  NAND2X0_LVT U10140 ( .A1(n8991), .A2(n_T_427[891]), .Y(n8909) );
  NAND2X0_LVT U10141 ( .A1(n_T_427[1019]), .A2(n3755), .Y(n8911) );
  OA21X1_LVT U10142 ( .A1(n4011), .A2(n3303), .A3(n8911), .Y(n8914) );
  NAND2X0_LVT U10143 ( .A1(n_T_427[1275]), .A2(n3638), .Y(n8913) );
  NAND2X0_LVT U10144 ( .A1(n3668), .A2(n_T_427[1147]), .Y(n8912) );
  NAND2X0_LVT U10145 ( .A1(n3689), .A2(n_T_427[1723]), .Y(n8915) );
  OA21X1_LVT U10146 ( .A1(n3410), .A2(n3747), .A3(n8915), .Y(n8918) );
  NAND2X0_LVT U10147 ( .A1(n3996), .A2(n_T_427[1339]), .Y(n8917) );
  NAND2X0_LVT U10148 ( .A1(n4002), .A2(n_T_427[1787]), .Y(n8916) );
  NAND2X0_LVT U10149 ( .A1(n3769), .A2(n_T_427[1531]), .Y(n8919) );
  OA21X1_LVT U10150 ( .A1(n4009), .A2(n3304), .A3(n8919), .Y(n8922) );
  NAND2X0_LVT U10151 ( .A1(n3618), .A2(n_T_427[1595]), .Y(n8921) );
  NAND2X0_LVT U10152 ( .A1(n3649), .A2(n_T_427[1659]), .Y(n8920) );
  OR3X1_LVT U10153 ( .A1(n8924), .A2(n8925), .A3(n8923), .Y(N740) );
  NAND2X0_LVT U10154 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[60]), .Y(n8929)
         );
  NAND2X0_LVT U10155 ( .A1(n9065), .A2(n_T_1165[60]), .Y(n8928) );
  NAND2X0_LVT U10156 ( .A1(n2493), .A2(n_T_628[60]), .Y(n8927) );
  NAND2X0_LVT U10157 ( .A1(n9066), .A2(n_T_918[60]), .Y(n8926) );
  NAND4X0_LVT U10158 ( .A1(n8929), .A2(n8928), .A3(n8927), .A4(n8926), .Y(
        io_fpu_fromint_data[60]) );
  NAND2X0_LVT U10159 ( .A1(n3789), .A2(n_T_427[317]), .Y(n8930) );
  OA21X1_LVT U10160 ( .A1(n3691), .A2(n3280), .A3(n8930), .Y(n8942) );
  AO22X1_LVT U10161 ( .A1(n4023), .A2(n_T_427[956]), .A3(n3976), .A4(
        n_T_427[573]), .Y(n8936) );
  AO22X1_LVT U10162 ( .A1(n3968), .A2(n_T_427[445]), .A3(n4020), .A4(
        n_T_427[701]), .Y(n8935) );
  AO22X1_LVT U10163 ( .A1(n2858), .A2(n_T_427[189]), .A3(n3979), .A4(
        n_T_427[828]), .Y(n8934) );
  AO22X1_LVT U10164 ( .A1(n4035), .A2(n_T_427[637]), .A3(n4027), .A4(
        n_T_427[892]), .Y(n8933) );
  NOR4X1_LVT U10165 ( .A1(n8936), .A2(n8935), .A3(n8934), .A4(n8933), .Y(n8938) );
  NAND2X0_LVT U10166 ( .A1(n2982), .A2(n4490), .Y(n8937) );
  OA21X1_LVT U10167 ( .A1(n8938), .A2(n3612), .A3(n8937), .Y(n8941) );
  NAND2X0_LVT U10168 ( .A1(n8939), .A2(n_T_427[381]), .Y(n8940) );
  NAND2X0_LVT U10169 ( .A1(n3745), .A2(n_T_427[253]), .Y(n8943) );
  NAND2X0_LVT U10170 ( .A1(n_T_427[509]), .A2(n3614), .Y(n8946) );
  NAND2X0_LVT U10171 ( .A1(n8944), .A2(n_T_427[61]), .Y(n8945) );
  NAND2X0_LVT U10172 ( .A1(n3605), .A2(n_T_427[1404]), .Y(n8947) );
  OA21X1_LVT U10173 ( .A1(n3167), .A2(n3987), .A3(n8947), .Y(n8950) );
  NAND2X0_LVT U10174 ( .A1(n2966), .A2(n_T_427[1468]), .Y(n8949) );
  NAND2X0_LVT U10175 ( .A1(n3991), .A2(n_T_427[1940]), .Y(n8948) );
  NAND2X0_LVT U10176 ( .A1(n3657), .A2(n_T_427[1724]), .Y(n8951) );
  OA21X1_LVT U10177 ( .A1(n3168), .A2(n3751), .A3(n8951), .Y(n8954) );
  NAND2X0_LVT U10178 ( .A1(n2094), .A2(n_T_427[1340]), .Y(n8953) );
  NAND2X0_LVT U10179 ( .A1(n4005), .A2(n_T_427[1788]), .Y(n8952) );
  NAND2X0_LVT U10180 ( .A1(n3770), .A2(n_T_427[1532]), .Y(n8955) );
  NAND2X0_LVT U10181 ( .A1(n3615), .A2(n_T_427[1596]), .Y(n8957) );
  NAND2X0_LVT U10182 ( .A1(n_T_427[1660]), .A2(n3650), .Y(n8956) );
  NAND2X0_LVT U10183 ( .A1(n3712), .A2(n_T_427[1020]), .Y(n8959) );
  OA21X1_LVT U10184 ( .A1(n4011), .A2(n3281), .A3(n8959), .Y(n8962) );
  NAND2X0_LVT U10185 ( .A1(n_T_427[1276]), .A2(n3638), .Y(n8961) );
  NAND2X0_LVT U10186 ( .A1(n3667), .A2(n_T_427[1148]), .Y(n8960) );
  NAND2X0_LVT U10187 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[61]), .Y(n8966)
         );
  NAND2X0_LVT U10188 ( .A1(n9065), .A2(n_T_1165[61]), .Y(n8965) );
  NAND2X0_LVT U10189 ( .A1(n2493), .A2(n_T_628[61]), .Y(n8964) );
  NAND2X0_LVT U10190 ( .A1(n9066), .A2(n_T_918[61]), .Y(n8963) );
  NAND4X0_LVT U10191 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .Y(
        io_fpu_fromint_data[61]) );
  NAND2X0_LVT U10192 ( .A1(n_T_427[1405]), .A2(n3608), .Y(n8967) );
  OA21X1_LVT U10193 ( .A1(n3169), .A2(n3989), .A3(n8967), .Y(n8970) );
  NAND2X0_LVT U10194 ( .A1(n3626), .A2(n_T_427[1469]), .Y(n8969) );
  NAND2X0_LVT U10195 ( .A1(n2986), .A2(n_T_427[1941]), .Y(n8968) );
  NAND2X0_LVT U10196 ( .A1(n3657), .A2(n_T_427[1725]), .Y(n8971) );
  OA21X1_LVT U10197 ( .A1(n3411), .A2(n3751), .A3(n8971), .Y(n8974) );
  NAND2X0_LVT U10198 ( .A1(n3998), .A2(n_T_427[1341]), .Y(n8973) );
  NAND2X0_LVT U10199 ( .A1(n4003), .A2(n_T_427[1789]), .Y(n8972) );
  NAND2X0_LVT U10200 ( .A1(n3770), .A2(n_T_427[1533]), .Y(n8975) );
  NAND2X0_LVT U10201 ( .A1(n3620), .A2(n_T_427[1597]), .Y(n8977) );
  NAND2X0_LVT U10202 ( .A1(n3650), .A2(n_T_427[1661]), .Y(n8976) );
  NAND2X0_LVT U10203 ( .A1(n3756), .A2(n_T_427[1021]), .Y(n8979) );
  NAND2X0_LVT U10204 ( .A1(n_T_427[318]), .A2(n3790), .Y(n8990) );
  NAND2X0_LVT U10205 ( .A1(n3665), .A2(n4493), .Y(n8989) );
  AO22X1_LVT U10206 ( .A1(n4023), .A2(n_T_427[957]), .A3(n3976), .A4(
        n_T_427[574]), .Y(n8986) );
  AO22X1_LVT U10207 ( .A1(n3979), .A2(n_T_427[829]), .A3(n4052), .A4(
        n_T_427[62]), .Y(n8985) );
  AO22X1_LVT U10208 ( .A1(n4034), .A2(n_T_427[638]), .A3(n3983), .A4(
        n_T_427[254]), .Y(n8984) );
  AO22X1_LVT U10209 ( .A1(n4039), .A2(n_T_427[382]), .A3(n4048), .A4(
        n_T_427[765]), .Y(n8983) );
  NOR4X1_LVT U10210 ( .A1(n8986), .A2(n8985), .A3(n8984), .A4(n8983), .Y(n8987) );
  NAND2X0_LVT U10211 ( .A1(n8991), .A2(n_T_427[893]), .Y(n8993) );
  NAND2X0_LVT U10212 ( .A1(n_T_427[510]), .A2(n9052), .Y(n8992) );
  NAND2X0_LVT U10213 ( .A1(n8994), .A2(n_T_427[126]), .Y(n8995) );
  OA21X1_LVT U10214 ( .A1(n3478), .A2(n8996), .A3(n8995), .Y(n8999) );
  NAND2X0_LVT U10215 ( .A1(n3713), .A2(n_T_427[190]), .Y(n8997) );
  NAND2X0_LVT U10216 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[62]), .Y(n9003)
         );
  NAND2X0_LVT U10217 ( .A1(n9065), .A2(n_T_1165[62]), .Y(n9002) );
  NAND2X0_LVT U10218 ( .A1(n2493), .A2(n_T_628[62]), .Y(n9001) );
  NAND2X0_LVT U10219 ( .A1(n9066), .A2(n_T_918[62]), .Y(n9000) );
  NAND4X0_LVT U10220 ( .A1(n9003), .A2(n9002), .A3(n9001), .A4(n9000), .Y(
        io_fpu_fromint_data[62]) );
  NAND2X0_LVT U10221 ( .A1(n3604), .A2(n_T_427[1406]), .Y(n9005) );
  NAND2X0_LVT U10222 ( .A1(n3626), .A2(n_T_427[1470]), .Y(n9010) );
  NAND2X0_LVT U10223 ( .A1(n3992), .A2(n_T_427[1942]), .Y(n9009) );
  NAND2X0_LVT U10224 ( .A1(n2922), .A2(n_T_427[1726]), .Y(n9013) );
  OA21X1_LVT U10225 ( .A1(n3171), .A2(n3747), .A3(n9013), .Y(n9019) );
  NAND2X0_LVT U10226 ( .A1(n3997), .A2(n_T_427[1342]), .Y(n9018) );
  NAND2X0_LVT U10227 ( .A1(n4003), .A2(n_T_427[1790]), .Y(n9017) );
  NAND2X0_LVT U10228 ( .A1(n3769), .A2(n_T_427[1534]), .Y(n9020) );
  OA21X1_LVT U10229 ( .A1(n3663), .A2(n3308), .A3(n9020), .Y(n9025) );
  NAND2X0_LVT U10230 ( .A1(n3620), .A2(n_T_427[1598]), .Y(n9024) );
  NAND3X0_LVT U10231 ( .A1(n9025), .A2(n9024), .A3(n9023), .Y(n9034) );
  NAND2X0_LVT U10232 ( .A1(n_T_427[1022]), .A2(n3761), .Y(n9027) );
  NAND2X0_LVT U10233 ( .A1(n3639), .A2(n_T_427[1278]), .Y(n9032) );
  NAND2X0_LVT U10234 ( .A1(n3674), .A2(n_T_427[1150]), .Y(n9031) );
  NAND2X0_LVT U10235 ( .A1(n3787), .A2(n_T_427[575]), .Y(n9051) );
  NAND2X0_LVT U10236 ( .A1(n3665), .A2(n4496), .Y(n9050) );
  AO22X1_LVT U10237 ( .A1(n4025), .A2(n_T_427[958]), .A3(n4018), .A4(
        n_T_427[703]), .Y(n9046) );
  AO22X1_LVT U10238 ( .A1(n4031), .A2(n_T_427[639]), .A3(n4028), .A4(
        n_T_427[894]), .Y(n9045) );
  AO22X1_LVT U10239 ( .A1(n4044), .A2(n_T_427[127]), .A3(n4038), .A4(
        n_T_427[383]), .Y(n9044) );
  AO22X1_LVT U10240 ( .A1(n4052), .A2(n_T_427[63]), .A3(n4045), .A4(
        n_T_427[766]), .Y(n9043) );
  NOR4X1_LVT U10241 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .Y(n9048) );
  NAND3X0_LVT U10242 ( .A1(n9051), .A2(n9050), .A3(n9049), .Y(n9063) );
  NAND2X0_LVT U10243 ( .A1(n_T_427[511]), .A2(n9052), .Y(n9055) );
  NAND2X0_LVT U10244 ( .A1(n3790), .A2(n_T_427[319]), .Y(n9054) );
  NAND2X0_LVT U10245 ( .A1(n9055), .A2(n9054), .Y(n9062) );
  NAND2X0_LVT U10246 ( .A1(n9056), .A2(n_T_427[830]), .Y(n9057) );
  NAND2X0_LVT U10247 ( .A1(n_T_427[255]), .A2(n3624), .Y(n9061) );
  NAND2X0_LVT U10248 ( .A1(n3714), .A2(n_T_427[191]), .Y(n9060) );
  NAND2X0_LVT U10249 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[63]), .Y(n9070)
         );
  NAND2X0_LVT U10250 ( .A1(n9065), .A2(n_T_1165[63]), .Y(n9069) );
  NAND2X0_LVT U10251 ( .A1(n2493), .A2(n_T_628[63]), .Y(n9068) );
  NAND2X0_LVT U10252 ( .A1(n9066), .A2(n_T_918[63]), .Y(n9067) );
  NAND4X0_LVT U10253 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .Y(
        io_fpu_fromint_data[63]) );
  MUX21X1_LVT U10254 ( .A1(n2553), .A2(io_fpu_inst[14]), .S0(io_fpu_inst[13]), 
        .Y(n9072) );
  NAND2X0_LVT U10255 ( .A1(n9107), .A2(n1891), .Y(n9071) );
  NAND2X0_LVT U10256 ( .A1(n9071), .A2(n9413), .Y(n9078) );
  AO21X1_LVT U10257 ( .A1(n9073), .A2(n9072), .A3(n9078), .Y(n9074) );
  AND2X1_LVT U10258 ( .A1(n2677), .A2(n9074), .Y(n1589) );
  NAND2X0_LVT U10259 ( .A1(n9087), .A2(io_fpu_inst[13]), .Y(n9085) );
  NAND2X0_LVT U10260 ( .A1(n9078), .A2(io_fpu_inst[13]), .Y(n9082) );
  NAND3X0_LVT U10261 ( .A1(n9082), .A2(n9081), .A3(n9080), .Y(n9083) );
  NAND2X0_LVT U10262 ( .A1(n2677), .A2(n9083), .Y(n9084) );
  NAND3X0_LVT U10263 ( .A1(n9084), .A2(n9228), .A3(n9085), .Y(N282) );
  NAND2X0_LVT U10264 ( .A1(n3079), .A2(n2618), .Y(n9086) );
  NAND2X0_LVT U10265 ( .A1(n9086), .A2(n9087), .Y(n9093) );
  NAND3X0_LVT U10266 ( .A1(n9093), .A2(n9233), .A3(n9229), .Y(N283) );
  INVX1_LVT U10267 ( .A(bpu_io_debug_if), .Y(n9242) );
  AO22X1_LVT U10268 ( .A1(io_fpu_inst[6]), .A2(io_fpu_inst[3]), .A3(n9097), 
        .A4(n1863), .Y(n9098) );
  NAND2X0_LVT U10269 ( .A1(n9116), .A2(n9098), .Y(n9100) );
  AO21X1_LVT U10270 ( .A1(n9103), .A2(io_fpu_fromint_data[40]), .A3(n9102), 
        .Y(alu_io_in1[40]) );
  AO21X1_LVT U10271 ( .A1(n9103), .A2(io_fpu_fromint_data[42]), .A3(n9102), 
        .Y(alu_io_in1[42]) );
  AO21X1_LVT U10272 ( .A1(n9103), .A2(io_fpu_fromint_data[44]), .A3(n9102), 
        .Y(alu_io_in1[44]) );
  AO21X1_LVT U10273 ( .A1(n9103), .A2(io_fpu_fromint_data[45]), .A3(n9102), 
        .Y(alu_io_in1[45]) );
  AO21X1_LVT U10274 ( .A1(n9103), .A2(io_fpu_fromint_data[46]), .A3(n9102), 
        .Y(alu_io_in1[46]) );
  AO21X1_LVT U10275 ( .A1(n9103), .A2(io_fpu_fromint_data[47]), .A3(n9102), 
        .Y(alu_io_in1[47]) );
  AO21X1_LVT U10276 ( .A1(n9103), .A2(io_fpu_fromint_data[48]), .A3(n9102), 
        .Y(alu_io_in1[48]) );
  AO21X1_LVT U10277 ( .A1(n9103), .A2(io_fpu_fromint_data[50]), .A3(n9102), 
        .Y(alu_io_in1[50]) );
  AO21X1_LVT U10278 ( .A1(n9103), .A2(io_fpu_fromint_data[52]), .A3(n9102), 
        .Y(alu_io_in1[52]) );
  AO21X1_LVT U10279 ( .A1(n9103), .A2(io_fpu_fromint_data[53]), .A3(n9102), 
        .Y(alu_io_in1[53]) );
  AO21X1_LVT U10280 ( .A1(n9103), .A2(io_fpu_fromint_data[54]), .A3(n9102), 
        .Y(alu_io_in1[54]) );
  AO21X1_LVT U10281 ( .A1(n9103), .A2(io_fpu_fromint_data[56]), .A3(n9102), 
        .Y(alu_io_in1[56]) );
  AO21X1_LVT U10282 ( .A1(n9103), .A2(io_fpu_fromint_data[57]), .A3(n9102), 
        .Y(alu_io_in1[57]) );
  AO21X1_LVT U10283 ( .A1(n9103), .A2(io_fpu_fromint_data[58]), .A3(n9102), 
        .Y(alu_io_in1[58]) );
  AO21X1_LVT U10284 ( .A1(n9103), .A2(io_fpu_fromint_data[59]), .A3(n9102), 
        .Y(alu_io_in1[59]) );
  AO21X1_LVT U10285 ( .A1(n9103), .A2(io_fpu_fromint_data[60]), .A3(n9102), 
        .Y(alu_io_in1[60]) );
  AO21X1_LVT U10286 ( .A1(n9103), .A2(io_fpu_fromint_data[61]), .A3(n9102), 
        .Y(alu_io_in1[61]) );
  AO21X1_LVT U10287 ( .A1(n9103), .A2(io_fpu_fromint_data[62]), .A3(n9102), 
        .Y(alu_io_in1[62]) );
  MUX21X1_LVT U10288 ( .A1(n9105), .A2(n1867), .S0(n1863), .Y(n9106) );
  AO21X1_LVT U10289 ( .A1(n9108), .A2(n9107), .A3(n9106), .Y(
        id_ctrl_sel_imm[2]) );
  NAND2X0_LVT U10290 ( .A1(n9110), .A2(io_fpu_inst[2]), .Y(n9114) );
  NAND2X0_LVT U10291 ( .A1(n9116), .A2(n9115), .Y(n9117) );
  NAND2X0_LVT U10292 ( .A1(n9117), .A2(n9430), .Y(n9119) );
  AND3X1_LVT U10293 ( .A1(n9119), .A2(n9118), .A3(n9244), .Y(N274) );
  AND2X1_LVT U10294 ( .A1(ex_ctrl_sel_alu2[1]), .A2(ex_ctrl_sel_alu2[0]), .Y(
        n9179) );
  NAND3X0_LVT U10295 ( .A1(n546), .A2(ex_ctrl_sel_imm[0]), .A3(
        ex_ctrl_sel_imm[2]), .Y(n9173) );
  AND2X1_LVT U10296 ( .A1(n9120), .A2(n9227), .Y(n9130) );
  AOI22X1_LVT U10297 ( .A1(n9144), .A2(n_T_648[3]), .A3(
        io_fpu_dmem_resp_data[0]), .A4(n9130), .Y(n9129) );
  NAND3X0_LVT U10298 ( .A1(n546), .A2(ex_ctrl_sel_imm[2]), .A3(n_T_642[0]), 
        .Y(n9121) );
  NAND2X0_LVT U10299 ( .A1(n3231), .A2(n546), .Y(n9172) );
  OA22X1_LVT U10300 ( .A1(n9121), .A2(n9201), .A3(n592), .A4(n9163), .Y(n9122)
         );
  OR2X1_LVT U10301 ( .A1(ex_ctrl_sel_imm[0]), .A2(n9122), .Y(n9128) );
  NAND3X0_LVT U10302 ( .A1(n9125), .A2(n9124), .A3(n9123), .Y(n9126) );
  NAND2X0_LVT U10303 ( .A1(n9227), .A2(n9126), .Y(n9127) );
  NAND3X0_LVT U10304 ( .A1(n9129), .A2(n9128), .A3(n9127), .Y(alu_io_in2[0])
         );
  OR2X1_LVT U10305 ( .A1(ex_ctrl_sel_imm[0]), .A2(n9178), .Y(n9200) );
  AND2X1_LVT U10306 ( .A1(n9199), .A2(n9172), .Y(n9158) );
  NAND2X0_LVT U10307 ( .A1(n9158), .A2(n_T_642[1]), .Y(n9141) );
  NAND2X0_LVT U10308 ( .A1(io_fpu_dmem_resp_data[1]), .A2(n9130), .Y(n9134) );
  NAND2X0_LVT U10309 ( .A1(ex_ctrl_sel_alu2[0]), .A2(n3278), .Y(n9142) );
  OR2X1_LVT U10310 ( .A1(n3215), .A2(n9142), .Y(n9131) );
  OA21X1_LVT U10311 ( .A1(n591), .A2(n9163), .A3(n9131), .Y(n9133) );
  NAND2X0_LVT U10312 ( .A1(n_T_648[4]), .A2(n9144), .Y(n9132) );
  AND3X1_LVT U10313 ( .A1(n9134), .A2(n9133), .A3(n9132), .Y(n9140) );
  NAND3X0_LVT U10314 ( .A1(n9137), .A2(n9136), .A3(n9135), .Y(n9138) );
  NAND2X0_LVT U10315 ( .A1(n9227), .A2(n9138), .Y(n9139) );
  NAND3X0_LVT U10316 ( .A1(n9141), .A2(n9140), .A3(n9139), .Y(alu_io_in2[1])
         );
  NAND2X0_LVT U10317 ( .A1(n_T_642[2]), .A2(n9158), .Y(n9154) );
  OR2X1_LVT U10318 ( .A1(ex_reg_rvc), .A2(n9142), .Y(n9143) );
  OA21X1_LVT U10319 ( .A1(n590), .A2(n9163), .A3(n9143), .Y(n9147) );
  NAND3X0_LVT U10320 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[2]), .A3(n9227), 
        .Y(n9146) );
  NAND2X0_LVT U10321 ( .A1(n9144), .A2(n_T_648[5]), .Y(n9145) );
  AND3X1_LVT U10322 ( .A1(n9147), .A2(n9146), .A3(n9145), .Y(n9153) );
  NAND3X0_LVT U10323 ( .A1(n9150), .A2(n9149), .A3(n9148), .Y(n9151) );
  NAND2X0_LVT U10324 ( .A1(n9227), .A2(n9151), .Y(n9152) );
  NAND3X0_LVT U10325 ( .A1(n9154), .A2(n9153), .A3(n9152), .Y(alu_io_in2[2])
         );
  NAND2X0_LVT U10326 ( .A1(n_T_642[4]), .A2(n9158), .Y(n9169) );
  NAND3X0_LVT U10327 ( .A1(n9161), .A2(n9160), .A3(n9159), .Y(n9162) );
  NAND2X0_LVT U10328 ( .A1(n9227), .A2(n9162), .Y(n9168) );
  OA22X1_LVT U10329 ( .A1(n160), .A2(n9164), .A3(n588), .A4(n9163), .Y(n9167)
         );
  NAND3X0_LVT U10330 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[4]), .A3(n9227), 
        .Y(n9166) );
  NAND4X0_LVT U10331 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .Y(
        alu_io_in2[4]) );
  AO22X1_LVT U10332 ( .A1(n_T_642[5]), .A2(n9199), .A3(n_T_702[5]), .A4(n9227), 
        .Y(alu_io_in2[5]) );
  AO22X1_LVT U10333 ( .A1(n_T_642[6]), .A2(n9199), .A3(n_T_702[6]), .A4(n9227), 
        .Y(alu_io_in2[6]) );
  AO22X1_LVT U10334 ( .A1(n_T_642[7]), .A2(n9199), .A3(n_T_702[7]), .A4(n9227), 
        .Y(alu_io_in2[7]) );
  AO22X1_LVT U10335 ( .A1(n_T_642[8]), .A2(n9199), .A3(n_T_702[8]), .A4(n9227), 
        .Y(alu_io_in2[8]) );
  AO22X1_LVT U10336 ( .A1(n_T_642[9]), .A2(n9199), .A3(n_T_702[9]), .A4(n9227), 
        .Y(alu_io_in2[9]) );
  AO22X1_LVT U10337 ( .A1(n_T_642[10]), .A2(n9199), .A3(n_T_702[10]), .A4(
        n9227), .Y(alu_io_in2[10]) );
  NAND2X0_LVT U10338 ( .A1(n9227), .A2(n_T_702[11]), .Y(n9177) );
  AND2X1_LVT U10339 ( .A1(io_dmem_req_bits_tag[1]), .A2(ex_ctrl_sel_imm[0]), 
        .Y(n9170) );
  MUX21X1_LVT U10340 ( .A1(n_T_642[0]), .A2(n9170), .S0(n546), .Y(n9171) );
  NAND3X0_LVT U10341 ( .A1(n9199), .A2(n3231), .A3(n9171), .Y(n9176) );
  NAND2X0_LVT U10342 ( .A1(n9178), .A2(n9226), .Y(n9197) );
  AO21X1_LVT U10343 ( .A1(n9174), .A2(ex_ctrl_sel_imm[0]), .A3(n9197), .Y(
        n9175) );
  NAND3X0_LVT U10344 ( .A1(n9177), .A2(n9176), .A3(n9175), .Y(alu_io_in2[11])
         );
  NAND2X0_LVT U10345 ( .A1(n9227), .A2(n_T_702[12]), .Y(n9182) );
  AND2X1_LVT U10346 ( .A1(n9180), .A2(n9179), .Y(n9195) );
  NAND2X0_LVT U10347 ( .A1(n9195), .A2(n_T_648[0]), .Y(n9181) );
  NAND3X0_LVT U10348 ( .A1(n9182), .A2(n9197), .A3(n9181), .Y(alu_io_in2[12])
         );
  NAND2X0_LVT U10349 ( .A1(n9227), .A2(n_T_702[13]), .Y(n9184) );
  NAND2X0_LVT U10350 ( .A1(n9195), .A2(n_T_648[1]), .Y(n9183) );
  NAND3X0_LVT U10351 ( .A1(n9184), .A2(n9197), .A3(n9183), .Y(alu_io_in2[13])
         );
  NAND2X0_LVT U10352 ( .A1(n9227), .A2(n_T_702[14]), .Y(n9186) );
  NAND2X0_LVT U10353 ( .A1(n9195), .A2(n_T_648[2]), .Y(n9185) );
  NAND3X0_LVT U10354 ( .A1(n9186), .A2(n9197), .A3(n9185), .Y(alu_io_in2[14])
         );
  NAND2X0_LVT U10355 ( .A1(n9227), .A2(n_T_702[15]), .Y(n9188) );
  NAND2X0_LVT U10356 ( .A1(n9195), .A2(n_T_648[3]), .Y(n9187) );
  NAND3X0_LVT U10357 ( .A1(n9188), .A2(n9197), .A3(n9187), .Y(alu_io_in2[15])
         );
  NAND2X0_LVT U10358 ( .A1(n9227), .A2(n_T_702[16]), .Y(n9190) );
  NAND2X0_LVT U10359 ( .A1(n9195), .A2(n_T_648[4]), .Y(n9189) );
  NAND3X0_LVT U10360 ( .A1(n9190), .A2(n9197), .A3(n9189), .Y(alu_io_in2[16])
         );
  NAND2X0_LVT U10361 ( .A1(n9227), .A2(n_T_702[17]), .Y(n9192) );
  NAND2X0_LVT U10362 ( .A1(n9195), .A2(n_T_648[5]), .Y(n9191) );
  NAND3X0_LVT U10363 ( .A1(n9192), .A2(n9197), .A3(n9191), .Y(alu_io_in2[17])
         );
  NAND2X0_LVT U10364 ( .A1(n9227), .A2(n_T_702[18]), .Y(n9194) );
  NAND2X0_LVT U10365 ( .A1(n9195), .A2(n_T_648[6]), .Y(n9193) );
  NAND3X0_LVT U10366 ( .A1(n9194), .A2(n9197), .A3(n9193), .Y(alu_io_in2[18])
         );
  NAND2X0_LVT U10367 ( .A1(n9227), .A2(n_T_702[19]), .Y(n9198) );
  NAND2X0_LVT U10368 ( .A1(n9195), .A2(n_T_648[7]), .Y(n9196) );
  NAND3X0_LVT U10369 ( .A1(n9198), .A2(n9197), .A3(n9196), .Y(alu_io_in2[19])
         );
  NAND2X0_LVT U10370 ( .A1(n9227), .A2(n_T_702[20]), .Y(n9203) );
  NAND2X0_LVT U10371 ( .A1(n9199), .A2(ex_reg_inst_31_), .Y(n9224) );
  NAND2X0_LVT U10372 ( .A1(n9222), .A2(n_T_642[0]), .Y(n9202) );
  NAND3X0_LVT U10373 ( .A1(n9203), .A2(n9224), .A3(n9202), .Y(alu_io_in2[20])
         );
  NAND2X0_LVT U10374 ( .A1(n9227), .A2(n_T_702[21]), .Y(n9205) );
  NAND2X0_LVT U10375 ( .A1(n9222), .A2(n_T_642[1]), .Y(n9204) );
  NAND3X0_LVT U10376 ( .A1(n9205), .A2(n9224), .A3(n9204), .Y(alu_io_in2[21])
         );
  NAND2X0_LVT U10377 ( .A1(n9227), .A2(n_T_702[22]), .Y(n9207) );
  NAND2X0_LVT U10378 ( .A1(n9222), .A2(n_T_642[2]), .Y(n9206) );
  NAND3X0_LVT U10379 ( .A1(n9207), .A2(n9224), .A3(n9206), .Y(alu_io_in2[22])
         );
  NAND2X0_LVT U10380 ( .A1(n9227), .A2(n_T_702[23]), .Y(n9209) );
  NAND2X0_LVT U10381 ( .A1(n9222), .A2(n_T_642[3]), .Y(n9208) );
  NAND3X0_LVT U10382 ( .A1(n9209), .A2(n9224), .A3(n9208), .Y(alu_io_in2[23])
         );
  NAND2X0_LVT U10383 ( .A1(n9227), .A2(n_T_702[24]), .Y(n9211) );
  NAND2X0_LVT U10384 ( .A1(n9222), .A2(n_T_642[4]), .Y(n9210) );
  NAND3X0_LVT U10385 ( .A1(n9211), .A2(n9224), .A3(n9210), .Y(alu_io_in2[24])
         );
  NAND2X0_LVT U10386 ( .A1(n9227), .A2(n_T_702[25]), .Y(n9213) );
  NAND2X0_LVT U10387 ( .A1(n9222), .A2(n_T_642[5]), .Y(n9212) );
  NAND3X0_LVT U10388 ( .A1(n9213), .A2(n9224), .A3(n9212), .Y(alu_io_in2[25])
         );
  NAND2X0_LVT U10389 ( .A1(n9227), .A2(n_T_702[26]), .Y(n9215) );
  NAND2X0_LVT U10390 ( .A1(n9222), .A2(n_T_642[6]), .Y(n9214) );
  NAND3X0_LVT U10391 ( .A1(n9215), .A2(n9224), .A3(n9214), .Y(alu_io_in2[26])
         );
  NAND2X0_LVT U10392 ( .A1(n9227), .A2(n_T_702[27]), .Y(n9217) );
  NAND2X0_LVT U10393 ( .A1(n9222), .A2(n_T_642[7]), .Y(n9216) );
  NAND3X0_LVT U10394 ( .A1(n9217), .A2(n9224), .A3(n9216), .Y(alu_io_in2[27])
         );
  NAND2X0_LVT U10395 ( .A1(n9227), .A2(n_T_702[28]), .Y(n9219) );
  NAND2X0_LVT U10396 ( .A1(n9222), .A2(n_T_642[8]), .Y(n9218) );
  NAND3X0_LVT U10397 ( .A1(n9219), .A2(n9224), .A3(n9218), .Y(alu_io_in2[28])
         );
  NAND2X0_LVT U10398 ( .A1(n9227), .A2(n_T_702[29]), .Y(n9221) );
  NAND2X0_LVT U10399 ( .A1(n9222), .A2(n_T_642[9]), .Y(n9220) );
  NAND3X0_LVT U10400 ( .A1(n9221), .A2(n9224), .A3(n9220), .Y(alu_io_in2[29])
         );
  NAND2X0_LVT U10401 ( .A1(n9227), .A2(n_T_702[30]), .Y(n9225) );
  NAND2X0_LVT U10402 ( .A1(n9222), .A2(n_T_642[10]), .Y(n9223) );
  NAND3X0_LVT U10403 ( .A1(n9225), .A2(n9224), .A3(n9223), .Y(alu_io_in2[30])
         );
  AO21X1_LVT U10404 ( .A1(n9227), .A2(n_T_702[31]), .A3(n9226), .Y(
        alu_io_in2[31]) );
  AO21X1_LVT U10405 ( .A1(n9227), .A2(n_T_702[32]), .A3(n9226), .Y(
        alu_io_in2[32]) );
  AO21X1_LVT U10406 ( .A1(n9227), .A2(n_T_702[33]), .A3(n9226), .Y(
        alu_io_in2[33]) );
  AO21X1_LVT U10407 ( .A1(n9227), .A2(n_T_702[34]), .A3(n9226), .Y(
        alu_io_in2[34]) );
  AO21X1_LVT U10408 ( .A1(n9227), .A2(n_T_702[35]), .A3(n9226), .Y(
        alu_io_in2[35]) );
  AO21X1_LVT U10409 ( .A1(n9227), .A2(n_T_702[36]), .A3(n9226), .Y(
        alu_io_in2[36]) );
  AO21X1_LVT U10410 ( .A1(n9227), .A2(n_T_702[37]), .A3(n9226), .Y(
        alu_io_in2[37]) );
  AO21X1_LVT U10411 ( .A1(n9227), .A2(n_T_702[38]), .A3(n9226), .Y(
        alu_io_in2[38]) );
  AO21X1_LVT U10412 ( .A1(n9227), .A2(n_T_702[39]), .A3(n9226), .Y(
        alu_io_in2[39]) );
  AO21X1_LVT U10413 ( .A1(n9227), .A2(n_T_702[40]), .A3(n9226), .Y(
        alu_io_in2[40]) );
  AO21X1_LVT U10414 ( .A1(n9227), .A2(n_T_702[41]), .A3(n9226), .Y(
        alu_io_in2[41]) );
  AO21X1_LVT U10415 ( .A1(n9227), .A2(n_T_702[42]), .A3(n9226), .Y(
        alu_io_in2[42]) );
  AO21X1_LVT U10416 ( .A1(n9227), .A2(n_T_702[43]), .A3(n9226), .Y(
        alu_io_in2[43]) );
  AO21X1_LVT U10417 ( .A1(n9227), .A2(n_T_702[44]), .A3(n9226), .Y(
        alu_io_in2[44]) );
  AO21X1_LVT U10418 ( .A1(n9227), .A2(n_T_702[45]), .A3(n9226), .Y(
        alu_io_in2[45]) );
  AO21X1_LVT U10419 ( .A1(n9227), .A2(n_T_702[46]), .A3(n9226), .Y(
        alu_io_in2[46]) );
  AO21X1_LVT U10420 ( .A1(n9227), .A2(n_T_702[47]), .A3(n9226), .Y(
        alu_io_in2[47]) );
  AO21X1_LVT U10421 ( .A1(n9227), .A2(n_T_702[48]), .A3(n9226), .Y(
        alu_io_in2[48]) );
  AO21X1_LVT U10422 ( .A1(n9227), .A2(n_T_702[49]), .A3(n9226), .Y(
        alu_io_in2[49]) );
  AO21X1_LVT U10423 ( .A1(n9227), .A2(n_T_702[50]), .A3(n9226), .Y(
        alu_io_in2[50]) );
  AO21X1_LVT U10424 ( .A1(n9227), .A2(n_T_702[51]), .A3(n9226), .Y(
        alu_io_in2[51]) );
  AO21X1_LVT U10425 ( .A1(n9227), .A2(n_T_702[52]), .A3(n9226), .Y(
        alu_io_in2[52]) );
  AO21X1_LVT U10426 ( .A1(n9227), .A2(n_T_702[53]), .A3(n9226), .Y(
        alu_io_in2[53]) );
  AO21X1_LVT U10427 ( .A1(n9227), .A2(n_T_702[54]), .A3(n9226), .Y(
        alu_io_in2[54]) );
  AO21X1_LVT U10428 ( .A1(n9227), .A2(n_T_702[55]), .A3(n9226), .Y(
        alu_io_in2[55]) );
  AO21X1_LVT U10429 ( .A1(n9227), .A2(n_T_702[56]), .A3(n9226), .Y(
        alu_io_in2[56]) );
  AO21X1_LVT U10430 ( .A1(n9227), .A2(n_T_702[57]), .A3(n9226), .Y(
        alu_io_in2[57]) );
  AO21X1_LVT U10431 ( .A1(n9227), .A2(n_T_702[58]), .A3(n9226), .Y(
        alu_io_in2[58]) );
  AO21X1_LVT U10432 ( .A1(n9227), .A2(n_T_702[59]), .A3(n9226), .Y(
        alu_io_in2[59]) );
  AO21X1_LVT U10433 ( .A1(n9227), .A2(n_T_702[60]), .A3(n9226), .Y(
        alu_io_in2[60]) );
  AO21X1_LVT U10434 ( .A1(n9227), .A2(n_T_702[61]), .A3(n9226), .Y(
        alu_io_in2[61]) );
  AO21X1_LVT U10435 ( .A1(n9227), .A2(n_T_702[62]), .A3(n9226), .Y(
        alu_io_in2[62]) );
  AO21X1_LVT U10436 ( .A1(n9227), .A2(n_T_702[63]), .A3(n9226), .Y(
        alu_io_in2[63]) );
  OA21X1_LVT U10437 ( .A1(io_fpu_inst[14]), .A2(n9229), .A3(n9228), .Y(n9234)
         );
  NAND3X0_LVT U10438 ( .A1(n9234), .A2(n9233), .A3(n9232), .Y(N284) );
  INVX1_LVT U10439 ( .A(n9237), .Y(n9235) );
  AO22X1_LVT U10440 ( .A1(n9235), .A2(n9425), .A3(mem_reg_cause[0]), .A4(n1279), .Y(N533) );
  NAND2X0_LVT U10441 ( .A1(n3262), .A2(wb_reg_cause[0]), .Y(n9236) );
  NAND2X0_LVT U10442 ( .A1(n9240), .A2(n9236), .Y(wb_cause[0]) );
  AND2X1_LVT U10443 ( .A1(n9425), .A2(n9237), .Y(n9238) );
  AO21X1_LVT U10444 ( .A1(mem_reg_cause[2]), .A2(n1279), .A3(n9238), .Y(N535)
         );
  OR2X1_LVT U10445 ( .A1(wb_reg_cause[2]), .A2(n576), .Y(wb_cause[2]) );
  AO21X1_LVT U10446 ( .A1(mem_reg_cause[3]), .A2(n1279), .A3(n9238), .Y(N536)
         );
  NAND2X0_LVT U10447 ( .A1(n9249), .A2(n9239), .Y(n9241) );
  OAI22X1_LVT U10448 ( .A1(n576), .A2(n3565), .A3(n9241), .A4(n9240), .Y(
        wb_cause[3]) );
  MUX21X1_LVT U10449 ( .A1(csr_io_interrupt_cause[1]), .A2(n9245), .S0(n9448), 
        .Y(N304) );
  AND2X1_LVT U10450 ( .A1(io_dmem_s2_xcpt_ae_st), .A2(n9246), .Y(n9248) );
  OA21X1_LVT U10451 ( .A1(io_dmem_s2_xcpt_pf_st), .A2(n9248), .A3(n9247), .Y(
        n9250) );
  OA21X1_LVT U10452 ( .A1(io_dmem_s2_xcpt_ma_st), .A2(n9250), .A3(n9249), .Y(
        n9251) );
  INVX1_LVT U10453 ( .A(wb_cause[2]), .Y(n9252) );
  AND2X1_LVT U10454 ( .A1(n3262), .A2(wb_reg_cause[63]), .Y(wb_cause[63]) );
  AND2X1_LVT U10455 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[0]), .Y(
        csr_io_tval[0]) );
  AND2X1_LVT U10456 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[1]), .Y(
        csr_io_tval[1]) );
  AND2X1_LVT U10457 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[2]), .Y(
        csr_io_tval[2]) );
  AND2X1_LVT U10458 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[3]), .Y(
        csr_io_tval[3]) );
  AND2X1_LVT U10459 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[4]), .Y(
        csr_io_tval[4]) );
  AND2X1_LVT U10460 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[5]), .Y(
        csr_io_tval[5]) );
  AND2X1_LVT U10461 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[6]), .Y(
        csr_io_tval[6]) );
  AND2X1_LVT U10462 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[7]), .Y(
        csr_io_tval[7]) );
  AND2X1_LVT U10463 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[8]), .Y(
        csr_io_tval[8]) );
  AND2X1_LVT U10464 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[9]), .Y(
        csr_io_tval[9]) );
  AND2X1_LVT U10465 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[10]), .Y(
        csr_io_tval[10]) );
  AND2X1_LVT U10466 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[11]), .Y(
        csr_io_tval[11]) );
  AND2X1_LVT U10467 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[12]), .Y(
        csr_io_tval[12]) );
  AND2X1_LVT U10468 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[13]), .Y(
        csr_io_tval[13]) );
  AND2X1_LVT U10469 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[14]), .Y(
        csr_io_tval[14]) );
  AND2X1_LVT U10470 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[15]), .Y(
        csr_io_tval[15]) );
  AND2X1_LVT U10471 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[16]), .Y(
        csr_io_tval[16]) );
  AND2X1_LVT U10472 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[17]), .Y(
        csr_io_tval[17]) );
  AND2X1_LVT U10473 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[18]), .Y(
        csr_io_tval[18]) );
  AND2X1_LVT U10474 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[19]), .Y(
        csr_io_tval[19]) );
  AND2X1_LVT U10475 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[20]), .Y(
        csr_io_tval[20]) );
  AND2X1_LVT U10476 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[21]), .Y(
        csr_io_tval[21]) );
  AND2X1_LVT U10477 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[22]), .Y(
        csr_io_tval[22]) );
  AND2X1_LVT U10478 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[23]), .Y(
        csr_io_tval[23]) );
  AND2X1_LVT U10479 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[24]), .Y(
        csr_io_tval[24]) );
  AND2X1_LVT U10480 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[25]), .Y(
        csr_io_tval[25]) );
  AND2X1_LVT U10481 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[26]), .Y(
        csr_io_tval[26]) );
  AND2X1_LVT U10482 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[27]), .Y(
        csr_io_tval[27]) );
  AND2X1_LVT U10483 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[28]), .Y(
        csr_io_tval[28]) );
  AND2X1_LVT U10484 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[29]), .Y(
        csr_io_tval[29]) );
  AND2X1_LVT U10485 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[30]), .Y(
        csr_io_tval[30]) );
  AND2X1_LVT U10486 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[31]), .Y(
        csr_io_tval[31]) );
  AND2X1_LVT U10487 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[32]), .Y(
        csr_io_tval[32]) );
  AND2X1_LVT U10488 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[33]), .Y(
        csr_io_tval[33]) );
  AND2X1_LVT U10489 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[34]), .Y(
        csr_io_tval[34]) );
  AND2X1_LVT U10490 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[35]), .Y(
        csr_io_tval[35]) );
  AND2X1_LVT U10491 ( .A1(n9276), .A2(io_imem_sfence_bits_addr[36]), .Y(
        csr_io_tval[36]) );
  AND2X1_LVT U10492 ( .A1(n9276), .A2(io_imem_sfence_bits_addr[37]), .Y(
        csr_io_tval[37]) );
  AND2X1_LVT U10493 ( .A1(n9276), .A2(io_imem_sfence_bits_addr[38]), .Y(
        csr_io_tval[38]) );
  NOR4X1_LVT U10494 ( .A1(n_T_1165[45]), .A2(n_T_1165[44]), .A3(n_T_1165[46]), 
        .A4(n_T_1165[47]), .Y(n9258) );
  NOR4X1_LVT U10495 ( .A1(n_T_1165[40]), .A2(n_T_1165[42]), .A3(n_T_1165[41]), 
        .A4(n_T_1165[43]), .Y(n9257) );
  NAND2X0_LVT U10496 ( .A1(n9258), .A2(n9257), .Y(n9264) );
  NOR4X1_LVT U10497 ( .A1(n_T_1165[57]), .A2(n_T_1165[56]), .A3(n_T_1165[58]), 
        .A4(n_T_1165[60]), .Y(n9262) );
  NOR4X1_LVT U10498 ( .A1(n_T_1165[52]), .A2(n_T_1165[54]), .A3(n_T_1165[53]), 
        .A4(n_T_1165[55]), .Y(n9261) );
  NOR4X1_LVT U10499 ( .A1(n_T_1165[48]), .A2(n_T_1165[49]), .A3(n_T_1165[51]), 
        .A4(n_T_1165[50]), .Y(n9260) );
  NOR4X1_LVT U10500 ( .A1(n_T_1165[59]), .A2(n_T_1165[61]), .A3(n_T_1165[63]), 
        .A4(n_T_1165[62]), .Y(n9259) );
  NAND4X0_LVT U10501 ( .A1(n9262), .A2(n9261), .A3(n9260), .A4(n9259), .Y(
        n9263) );
  OR2X1_LVT U10502 ( .A1(n9264), .A2(n9263), .Y(n9273) );
  NAND4X0_LVT U10503 ( .A1(n_T_1165[61]), .A2(n_T_1165[63]), .A3(n_T_1165[62]), 
        .A4(n_T_1165[59]), .Y(n9268) );
  NAND4X0_LVT U10504 ( .A1(n_T_1165[57]), .A2(n_T_1165[56]), .A3(n_T_1165[58]), 
        .A4(n_T_1165[60]), .Y(n9267) );
  NAND4X0_LVT U10505 ( .A1(n_T_1165[52]), .A2(n_T_1165[54]), .A3(n_T_1165[53]), 
        .A4(n_T_1165[55]), .Y(n9266) );
  NAND4X0_LVT U10506 ( .A1(n_T_1165[48]), .A2(n_T_1165[49]), .A3(n_T_1165[51]), 
        .A4(n_T_1165[50]), .Y(n9265) );
  NOR4X1_LVT U10507 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .Y(n9271) );
  AND4X1_LVT U10508 ( .A1(n_T_1165[45]), .A2(n_T_1165[44]), .A3(n_T_1165[46]), 
        .A4(n_T_1165[47]), .Y(n9270) );
  AND4X1_LVT U10509 ( .A1(n_T_1165[40]), .A2(n_T_1165[42]), .A3(n_T_1165[41]), 
        .A4(n_T_1165[43]), .Y(n9269) );
  NAND3X0_LVT U10510 ( .A1(n9271), .A2(n9270), .A3(n9269), .Y(n9272) );
  MUX21X1_LVT U10511 ( .A1(n9273), .A2(n9272), .S0(n_T_1165[39]), .Y(n9274) );
  MUX21X1_LVT U10512 ( .A1(n_T_1165[39]), .A2(n3228), .S0(n9274), .Y(n9275) );
  AND2X1_LVT U10513 ( .A1(n9276), .A2(n9275), .Y(csr_io_tval[39]) );
  AND2X1_LVT U10514 ( .A1(wb_reg_valid), .A2(wb_ctrl_csr[2]), .Y(
        csr_io_rw_cmd_2_) );
  NAND3X0_LVT U10515 ( .A1(n9279), .A2(n9278), .A3(n9277), .Y(n9284) );
  NOR3X0_LVT U10516 ( .A1(mem_reg_valid), .A2(mem_reg_xcpt_interrupt), .A3(
        mem_reg_replay), .Y(n9449) );
  INVX1_LVT U10517 ( .A(n9449), .Y(mem_pc_valid) );
  AND2X1_LVT U10518 ( .A1(wb_reg_valid), .A2(wb_reg_sfence), .Y(
        io_imem_sfence_valid) );
  MUX21X1_LVT U10519 ( .A1(mem_reg_rs2[0]), .A2(io_fpu_store_data[0]), .S0(
        n2498), .Y(io_dmem_s1_data_data[0]) );
  MUX21X1_LVT U10520 ( .A1(mem_reg_rs2[1]), .A2(io_fpu_store_data[1]), .S0(
        n2498), .Y(io_dmem_s1_data_data[1]) );
  MUX21X1_LVT U10521 ( .A1(mem_reg_rs2[2]), .A2(io_fpu_store_data[2]), .S0(
        n2498), .Y(io_dmem_s1_data_data[2]) );
  MUX21X1_LVT U10522 ( .A1(mem_reg_rs2[3]), .A2(io_fpu_store_data[3]), .S0(
        n2498), .Y(io_dmem_s1_data_data[3]) );
  MUX21X1_LVT U10523 ( .A1(mem_reg_rs2[4]), .A2(io_fpu_store_data[4]), .S0(
        n2492), .Y(io_dmem_s1_data_data[4]) );
  MUX21X1_LVT U10524 ( .A1(mem_reg_rs2[5]), .A2(io_fpu_store_data[5]), .S0(
        n2498), .Y(io_dmem_s1_data_data[5]) );
  MUX21X1_LVT U10525 ( .A1(mem_reg_rs2[6]), .A2(io_fpu_store_data[6]), .S0(
        n2498), .Y(io_dmem_s1_data_data[6]) );
  MUX21X1_LVT U10526 ( .A1(mem_reg_rs2[7]), .A2(io_fpu_store_data[7]), .S0(
        n2498), .Y(io_dmem_s1_data_data[7]) );
  NAND2X0_LVT U10527 ( .A1(n313), .A2(io_dmem_req_bits_size[1]), .Y(n9292) );
  NAND2X0_LVT U10528 ( .A1(n586), .A2(io_dmem_req_bits_size[0]), .Y(n9289) );
  NAND2X0_LVT U10529 ( .A1(n9292), .A2(n9289), .Y(n9290) );
  AO22X1_LVT U10530 ( .A1(n_T_702[8]), .A2(n9290), .A3(n9291), .A4(n_T_702[0]), 
        .Y(n9293) );
  AO21X1_LVT U10531 ( .A1(n4058), .A2(n_T_702[8]), .A3(n9293), .Y(N469) );
  MUX21X1_LVT U10532 ( .A1(mem_reg_rs2[8]), .A2(io_fpu_store_data[8]), .S0(
        n2492), .Y(io_dmem_s1_data_data[8]) );
  AO22X1_LVT U10533 ( .A1(n_T_702[9]), .A2(n9290), .A3(n9291), .A4(n_T_702[1]), 
        .Y(n9295) );
  AO21X1_LVT U10534 ( .A1(n4058), .A2(n_T_702[9]), .A3(n9295), .Y(N470) );
  MUX21X1_LVT U10535 ( .A1(mem_reg_rs2[9]), .A2(io_fpu_store_data[9]), .S0(
        n2498), .Y(io_dmem_s1_data_data[9]) );
  AO22X1_LVT U10536 ( .A1(n_T_702[10]), .A2(n9290), .A3(n9291), .A4(n_T_702[2]), .Y(n9296) );
  AO21X1_LVT U10537 ( .A1(n4058), .A2(n_T_702[10]), .A3(n9296), .Y(N471) );
  MUX21X1_LVT U10538 ( .A1(mem_reg_rs2[10]), .A2(io_fpu_store_data[10]), .S0(
        n2498), .Y(io_dmem_s1_data_data[10]) );
  AO22X1_LVT U10539 ( .A1(n_T_702[11]), .A2(n9290), .A3(n9291), .A4(n_T_702[3]), .Y(n9297) );
  AO21X1_LVT U10540 ( .A1(n4058), .A2(n_T_702[11]), .A3(n9297), .Y(N472) );
  MUX21X1_LVT U10541 ( .A1(mem_reg_rs2[11]), .A2(io_fpu_store_data[11]), .S0(
        n2498), .Y(io_dmem_s1_data_data[11]) );
  AO22X1_LVT U10542 ( .A1(n_T_702[12]), .A2(n9290), .A3(n9291), .A4(n_T_702[4]), .Y(n9298) );
  AO21X1_LVT U10543 ( .A1(n4058), .A2(n_T_702[12]), .A3(n9298), .Y(N473) );
  MUX21X1_LVT U10544 ( .A1(mem_reg_rs2[12]), .A2(io_fpu_store_data[12]), .S0(
        n2498), .Y(io_dmem_s1_data_data[12]) );
  AO22X1_LVT U10545 ( .A1(n_T_702[5]), .A2(n9291), .A3(n9290), .A4(n_T_702[13]), .Y(n9299) );
  AO21X1_LVT U10546 ( .A1(n4058), .A2(n_T_702[13]), .A3(n9299), .Y(N474) );
  MUX21X1_LVT U10547 ( .A1(mem_reg_rs2[13]), .A2(io_fpu_store_data[13]), .S0(
        n2498), .Y(io_dmem_s1_data_data[13]) );
  AO22X1_LVT U10548 ( .A1(n_T_702[6]), .A2(n9291), .A3(n9290), .A4(n_T_702[14]), .Y(n9300) );
  AO21X1_LVT U10549 ( .A1(n4058), .A2(n_T_702[14]), .A3(n9300), .Y(N475) );
  MUX21X1_LVT U10550 ( .A1(mem_reg_rs2[14]), .A2(io_fpu_store_data[14]), .S0(
        n2498), .Y(io_dmem_s1_data_data[14]) );
  AO22X1_LVT U10551 ( .A1(n_T_702[7]), .A2(n9291), .A3(n9290), .A4(n_T_702[15]), .Y(n9302) );
  AO21X1_LVT U10552 ( .A1(n4058), .A2(n_T_702[15]), .A3(n9302), .Y(N476) );
  MUX21X1_LVT U10553 ( .A1(mem_reg_rs2[15]), .A2(io_fpu_store_data[15]), .S0(
        n2498), .Y(io_dmem_s1_data_data[15]) );
  MUX21X1_LVT U10554 ( .A1(n_T_702[16]), .A2(n_T_702[0]), .S0(n586), .Y(N477)
         );
  MUX21X1_LVT U10555 ( .A1(mem_reg_rs2[16]), .A2(io_fpu_store_data[16]), .S0(
        n2492), .Y(io_dmem_s1_data_data[16]) );
  MUX21X1_LVT U10556 ( .A1(n_T_702[17]), .A2(n_T_702[1]), .S0(n2515), .Y(N478)
         );
  MUX21X1_LVT U10557 ( .A1(mem_reg_rs2[17]), .A2(io_fpu_store_data[17]), .S0(
        n2498), .Y(io_dmem_s1_data_data[17]) );
  MUX21X1_LVT U10558 ( .A1(n_T_702[18]), .A2(n_T_702[2]), .S0(n586), .Y(N479)
         );
  MUX21X1_LVT U10559 ( .A1(mem_reg_rs2[18]), .A2(io_fpu_store_data[18]), .S0(
        n2498), .Y(io_dmem_s1_data_data[18]) );
  MUX21X1_LVT U10560 ( .A1(n_T_702[19]), .A2(n_T_702[3]), .S0(n2515), .Y(N480)
         );
  MUX21X1_LVT U10561 ( .A1(mem_reg_rs2[19]), .A2(io_fpu_store_data[19]), .S0(
        n2498), .Y(io_dmem_s1_data_data[19]) );
  MUX21X1_LVT U10562 ( .A1(n_T_702[20]), .A2(n_T_702[4]), .S0(n586), .Y(N481)
         );
  MUX21X1_LVT U10563 ( .A1(mem_reg_rs2[20]), .A2(io_fpu_store_data[20]), .S0(
        n2498), .Y(io_dmem_s1_data_data[20]) );
  MUX21X1_LVT U10564 ( .A1(n_T_702[5]), .A2(n_T_702[21]), .S0(
        io_dmem_req_bits_size[1]), .Y(N482) );
  MUX21X1_LVT U10565 ( .A1(mem_reg_rs2[21]), .A2(io_fpu_store_data[21]), .S0(
        n2498), .Y(io_dmem_s1_data_data[21]) );
  MUX21X1_LVT U10566 ( .A1(n_T_702[6]), .A2(n_T_702[22]), .S0(
        io_dmem_req_bits_size[1]), .Y(N483) );
  MUX21X1_LVT U10567 ( .A1(mem_reg_rs2[22]), .A2(io_fpu_store_data[22]), .S0(
        n2498), .Y(io_dmem_s1_data_data[22]) );
  MUX21X1_LVT U10568 ( .A1(n_T_702[7]), .A2(n_T_702[23]), .S0(
        io_dmem_req_bits_size[1]), .Y(N484) );
  MUX21X1_LVT U10569 ( .A1(mem_reg_rs2[23]), .A2(io_fpu_store_data[23]), .S0(
        n2498), .Y(io_dmem_s1_data_data[23]) );
  MUX21X1_LVT U10570 ( .A1(n_T_702[24]), .A2(n9293), .S0(n586), .Y(N485) );
  MUX21X1_LVT U10571 ( .A1(mem_reg_rs2[24]), .A2(io_fpu_store_data[24]), .S0(
        n2498), .Y(io_dmem_s1_data_data[24]) );
  MUX21X1_LVT U10572 ( .A1(n_T_702[25]), .A2(n9295), .S0(n586), .Y(N486) );
  MUX21X1_LVT U10573 ( .A1(mem_reg_rs2[25]), .A2(io_fpu_store_data[25]), .S0(
        n2498), .Y(io_dmem_s1_data_data[25]) );
  MUX21X1_LVT U10574 ( .A1(n_T_702[26]), .A2(n9296), .S0(n586), .Y(N487) );
  MUX21X1_LVT U10575 ( .A1(mem_reg_rs2[26]), .A2(io_fpu_store_data[26]), .S0(
        n2498), .Y(io_dmem_s1_data_data[26]) );
  MUX21X1_LVT U10576 ( .A1(n_T_702[27]), .A2(n9297), .S0(n586), .Y(N488) );
  MUX21X1_LVT U10577 ( .A1(mem_reg_rs2[27]), .A2(io_fpu_store_data[27]), .S0(
        n2498), .Y(io_dmem_s1_data_data[27]) );
  MUX21X1_LVT U10578 ( .A1(n_T_702[28]), .A2(n9298), .S0(n586), .Y(N489) );
  MUX21X1_LVT U10579 ( .A1(mem_reg_rs2[28]), .A2(io_fpu_store_data[28]), .S0(
        n2498), .Y(io_dmem_s1_data_data[28]) );
  MUX21X1_LVT U10580 ( .A1(n_T_702[29]), .A2(n9299), .S0(n586), .Y(N490) );
  MUX21X1_LVT U10581 ( .A1(mem_reg_rs2[29]), .A2(io_fpu_store_data[29]), .S0(
        n2498), .Y(io_dmem_s1_data_data[29]) );
  MUX21X1_LVT U10582 ( .A1(n_T_702[30]), .A2(n9300), .S0(n586), .Y(N491) );
  MUX21X1_LVT U10583 ( .A1(mem_reg_rs2[30]), .A2(io_fpu_store_data[30]), .S0(
        n2498), .Y(io_dmem_s1_data_data[30]) );
  MUX21X1_LVT U10584 ( .A1(n_T_702[31]), .A2(n9302), .S0(n2515), .Y(N492) );
  MUX21X1_LVT U10585 ( .A1(mem_reg_rs2[31]), .A2(io_fpu_store_data[31]), .S0(
        n2492), .Y(io_dmem_s1_data_data[31]) );
  MUX21X1_LVT U10586 ( .A1(n_T_702[32]), .A2(n_T_702[0]), .S0(n3234), .Y(N493)
         );
  MUX21X1_LVT U10587 ( .A1(mem_reg_rs2[32]), .A2(io_fpu_store_data[32]), .S0(
        n2498), .Y(io_dmem_s1_data_data[32]) );
  MUX21X1_LVT U10588 ( .A1(n_T_702[33]), .A2(n_T_702[1]), .S0(n3234), .Y(N494)
         );
  MUX21X1_LVT U10589 ( .A1(mem_reg_rs2[33]), .A2(io_fpu_store_data[33]), .S0(
        n2498), .Y(io_dmem_s1_data_data[33]) );
  MUX21X1_LVT U10590 ( .A1(n_T_702[34]), .A2(n_T_702[2]), .S0(n3234), .Y(N495)
         );
  MUX21X1_LVT U10591 ( .A1(mem_reg_rs2[34]), .A2(io_fpu_store_data[34]), .S0(
        n2498), .Y(io_dmem_s1_data_data[34]) );
  MUX21X1_LVT U10592 ( .A1(n_T_702[35]), .A2(n_T_702[3]), .S0(n3234), .Y(N496)
         );
  MUX21X1_LVT U10593 ( .A1(mem_reg_rs2[35]), .A2(io_fpu_store_data[35]), .S0(
        n2492), .Y(io_dmem_s1_data_data[35]) );
  MUX21X1_LVT U10594 ( .A1(n_T_702[36]), .A2(n_T_702[4]), .S0(n3234), .Y(N497)
         );
  MUX21X1_LVT U10595 ( .A1(mem_reg_rs2[36]), .A2(io_fpu_store_data[36]), .S0(
        n2498), .Y(io_dmem_s1_data_data[36]) );
  MUX21X1_LVT U10596 ( .A1(n_T_702[37]), .A2(n_T_702[5]), .S0(n3234), .Y(N498)
         );
  MUX21X1_LVT U10597 ( .A1(mem_reg_rs2[37]), .A2(io_fpu_store_data[37]), .S0(
        n2498), .Y(io_dmem_s1_data_data[37]) );
  MUX21X1_LVT U10598 ( .A1(n_T_702[38]), .A2(n_T_702[6]), .S0(n3234), .Y(N499)
         );
  MUX21X1_LVT U10599 ( .A1(mem_reg_rs2[38]), .A2(io_fpu_store_data[38]), .S0(
        n2498), .Y(io_dmem_s1_data_data[38]) );
  MUX21X1_LVT U10600 ( .A1(n_T_702[39]), .A2(n_T_702[7]), .S0(n3234), .Y(N500)
         );
  MUX21X1_LVT U10601 ( .A1(mem_reg_rs2[39]), .A2(io_fpu_store_data[39]), .S0(
        n2492), .Y(io_dmem_s1_data_data[39]) );
  AO21X1_LVT U10602 ( .A1(n4058), .A2(n_T_702[40]), .A3(n9293), .Y(N501) );
  MUX21X1_LVT U10603 ( .A1(mem_reg_rs2[40]), .A2(io_fpu_store_data[40]), .S0(
        n2498), .Y(io_dmem_s1_data_data[40]) );
  AO21X1_LVT U10604 ( .A1(n4058), .A2(n_T_702[41]), .A3(n9295), .Y(N502) );
  MUX21X1_LVT U10605 ( .A1(mem_reg_rs2[41]), .A2(io_fpu_store_data[41]), .S0(
        n2498), .Y(io_dmem_s1_data_data[41]) );
  AO21X1_LVT U10606 ( .A1(n4058), .A2(n_T_702[42]), .A3(n9296), .Y(N503) );
  MUX21X1_LVT U10607 ( .A1(mem_reg_rs2[42]), .A2(io_fpu_store_data[42]), .S0(
        n2498), .Y(io_dmem_s1_data_data[42]) );
  AO21X1_LVT U10608 ( .A1(n4058), .A2(n_T_702[43]), .A3(n9297), .Y(N504) );
  MUX21X1_LVT U10609 ( .A1(mem_reg_rs2[43]), .A2(io_fpu_store_data[43]), .S0(
        n2492), .Y(io_dmem_s1_data_data[43]) );
  AO21X1_LVT U10610 ( .A1(n4058), .A2(n_T_702[44]), .A3(n9298), .Y(N505) );
  MUX21X1_LVT U10611 ( .A1(mem_reg_rs2[44]), .A2(io_fpu_store_data[44]), .S0(
        n2498), .Y(io_dmem_s1_data_data[44]) );
  AO21X1_LVT U10612 ( .A1(n4058), .A2(n_T_702[45]), .A3(n9299), .Y(N506) );
  MUX21X1_LVT U10613 ( .A1(mem_reg_rs2[45]), .A2(io_fpu_store_data[45]), .S0(
        n2498), .Y(io_dmem_s1_data_data[45]) );
  AO21X1_LVT U10614 ( .A1(n4058), .A2(n_T_702[46]), .A3(n9300), .Y(N507) );
  MUX21X1_LVT U10615 ( .A1(mem_reg_rs2[46]), .A2(io_fpu_store_data[46]), .S0(
        n2498), .Y(io_dmem_s1_data_data[46]) );
  AO21X1_LVT U10616 ( .A1(n4058), .A2(n_T_702[47]), .A3(n9302), .Y(N508) );
  MUX21X1_LVT U10617 ( .A1(mem_reg_rs2[47]), .A2(io_fpu_store_data[47]), .S0(
        n2492), .Y(io_dmem_s1_data_data[47]) );
  MUX21X1_LVT U10618 ( .A1(mem_reg_rs2[48]), .A2(io_fpu_store_data[48]), .S0(
        n2498), .Y(io_dmem_s1_data_data[48]) );
  MUX21X1_LVT U10619 ( .A1(mem_reg_rs2[49]), .A2(io_fpu_store_data[49]), .S0(
        n2498), .Y(io_dmem_s1_data_data[49]) );
  MUX21X1_LVT U10620 ( .A1(mem_reg_rs2[50]), .A2(io_fpu_store_data[50]), .S0(
        n2498), .Y(io_dmem_s1_data_data[50]) );
  MUX21X1_LVT U10621 ( .A1(mem_reg_rs2[51]), .A2(io_fpu_store_data[51]), .S0(
        n2492), .Y(io_dmem_s1_data_data[51]) );
  MUX21X1_LVT U10622 ( .A1(mem_reg_rs2[52]), .A2(io_fpu_store_data[52]), .S0(
        n2492), .Y(io_dmem_s1_data_data[52]) );
  MUX21X1_LVT U10623 ( .A1(mem_reg_rs2[53]), .A2(io_fpu_store_data[53]), .S0(
        n2498), .Y(io_dmem_s1_data_data[53]) );
  MUX21X1_LVT U10624 ( .A1(mem_reg_rs2[54]), .A2(io_fpu_store_data[54]), .S0(
        n2498), .Y(io_dmem_s1_data_data[54]) );
  MUX21X1_LVT U10625 ( .A1(mem_reg_rs2[55]), .A2(io_fpu_store_data[55]), .S0(
        n2498), .Y(io_dmem_s1_data_data[55]) );
  MUX21X1_LVT U10626 ( .A1(mem_reg_rs2[56]), .A2(io_fpu_store_data[56]), .S0(
        n2492), .Y(io_dmem_s1_data_data[56]) );
  AO22X1_LVT U10627 ( .A1(n_T_702[57]), .A2(n4058), .A3(n9301), .A4(
        n_T_702[25]), .Y(n9294) );
  AO21X1_LVT U10628 ( .A1(n2515), .A2(n9295), .A3(n9294), .Y(N518) );
  MUX21X1_LVT U10629 ( .A1(mem_reg_rs2[57]), .A2(io_fpu_store_data[57]), .S0(
        n2498), .Y(io_dmem_s1_data_data[57]) );
  MUX21X1_LVT U10630 ( .A1(mem_reg_rs2[58]), .A2(io_fpu_store_data[58]), .S0(
        n2498), .Y(io_dmem_s1_data_data[58]) );
  MUX21X1_LVT U10631 ( .A1(mem_reg_rs2[59]), .A2(io_fpu_store_data[59]), .S0(
        n2498), .Y(io_dmem_s1_data_data[59]) );
  MUX21X1_LVT U10632 ( .A1(mem_reg_rs2[60]), .A2(io_fpu_store_data[60]), .S0(
        n2492), .Y(io_dmem_s1_data_data[60]) );
  MUX21X1_LVT U10633 ( .A1(mem_reg_rs2[61]), .A2(io_fpu_store_data[61]), .S0(
        n2498), .Y(io_dmem_s1_data_data[61]) );
  MUX21X1_LVT U10634 ( .A1(mem_reg_rs2[62]), .A2(io_fpu_store_data[62]), .S0(
        n2498), .Y(io_dmem_s1_data_data[62]) );
  MUX21X1_LVT U10635 ( .A1(mem_reg_rs2[63]), .A2(io_fpu_store_data[63]), .S0(
        n2498), .Y(io_dmem_s1_data_data[63]) );
  NAND4X0_LVT U10636 ( .A1(n9306), .A2(n9305), .A3(n9304), .A4(n9303), .Y(
        n9317) );
  NAND4X0_LVT U10637 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .Y(
        n9316) );
  NOR4X1_LVT U10638 ( .A1(io_fpu_fromint_data[40]), .A2(
        io_fpu_fromint_data[42]), .A3(io_fpu_fromint_data[41]), .A4(
        io_fpu_fromint_data[43]), .Y(n9314) );
  NOR4X1_LVT U10639 ( .A1(io_fpu_fromint_data[45]), .A2(
        io_fpu_fromint_data[44]), .A3(io_fpu_fromint_data[46]), .A4(
        io_fpu_fromint_data[48]), .Y(n9313) );
  NOR4X1_LVT U10640 ( .A1(io_fpu_fromint_data[47]), .A2(
        io_fpu_fromint_data[49]), .A3(io_fpu_fromint_data[51]), .A4(
        io_fpu_fromint_data[50]), .Y(n9312) );
  NOR4X1_LVT U10641 ( .A1(io_fpu_fromint_data[52]), .A2(
        io_fpu_fromint_data[54]), .A3(io_fpu_fromint_data[53]), .A4(
        io_fpu_fromint_data[55]), .Y(n9311) );
  NAND4X0_LVT U10642 ( .A1(n9314), .A2(n9313), .A3(n9312), .A4(n9311), .Y(
        n9315) );
  OR3X1_LVT U10643 ( .A1(n9317), .A2(n9316), .A3(n9315), .Y(n9326) );
  NAND4X0_LVT U10644 ( .A1(io_fpu_fromint_data[57]), .A2(
        io_fpu_fromint_data[56]), .A3(io_fpu_fromint_data[58]), .A4(
        io_fpu_fromint_data[60]), .Y(n9324) );
  NAND4X0_LVT U10645 ( .A1(io_fpu_fromint_data[59]), .A2(
        io_fpu_fromint_data[61]), .A3(io_fpu_fromint_data[63]), .A4(
        io_fpu_fromint_data[62]), .Y(n9323) );
  AND4X1_LVT U10646 ( .A1(io_fpu_fromint_data[40]), .A2(
        io_fpu_fromint_data[42]), .A3(io_fpu_fromint_data[41]), .A4(
        io_fpu_fromint_data[43]), .Y(n9321) );
  AND4X1_LVT U10647 ( .A1(io_fpu_fromint_data[45]), .A2(
        io_fpu_fromint_data[44]), .A3(io_fpu_fromint_data[46]), .A4(
        io_fpu_fromint_data[48]), .Y(n9320) );
  AND4X1_LVT U10648 ( .A1(io_fpu_fromint_data[47]), .A2(
        io_fpu_fromint_data[49]), .A3(io_fpu_fromint_data[51]), .A4(
        io_fpu_fromint_data[50]), .Y(n9319) );
  AND4X1_LVT U10649 ( .A1(io_fpu_fromint_data[52]), .A2(
        io_fpu_fromint_data[54]), .A3(io_fpu_fromint_data[53]), .A4(
        io_fpu_fromint_data[55]), .Y(n9318) );
  NAND4X0_LVT U10650 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .Y(
        n9322) );
  OR3X1_LVT U10651 ( .A1(n9324), .A2(n9323), .A3(n9322), .Y(n9325) );
  MUX21X1_LVT U10652 ( .A1(n9326), .A2(n9325), .S0(io_fpu_fromint_data[39]), 
        .Y(n9327) );
  MUX21X1_LVT U10653 ( .A1(alu_io_adder_out_39_), .A2(n9328), .S0(n9327), .Y(
        io_dmem_req_bits_addr[39]) );
  NAND4X0_LVT U10654 ( .A1(n3310), .A2(n3104), .A3(
        io_imem_bht_update_bits_branch), .A4(n555), .Y(n9329) );
  INVX1_LVT U10655 ( .A(n9512), .Y(n9333) );
  AO222X1_LVT U10656 ( .A1(n4065), .A2(csr_io_evec[1]), .A3(n4062), .A4(
        csr_io_pc[1]), .A5(n9333), .A6(n4060), .Y(io_imem_req_bits_pc[1]) );
  AO22X1_LVT U10657 ( .A1(n4063), .A2(csr_io_pc[2]), .A3(n9334), .A4(n4060), 
        .Y(n9335) );
  AO21X1_LVT U10658 ( .A1(n4067), .A2(csr_io_evec[2]), .A3(n9335), .Y(
        io_imem_req_bits_pc[2]) );
  AO22X1_LVT U10659 ( .A1(n4064), .A2(csr_io_pc[3]), .A3(n9336), .A4(n4061), 
        .Y(n9337) );
  AO21X1_LVT U10660 ( .A1(n4067), .A2(csr_io_evec[3]), .A3(n9337), .Y(
        io_imem_req_bits_pc[3]) );
  AO22X1_LVT U10661 ( .A1(n4064), .A2(csr_io_pc[4]), .A3(n9338), .A4(n4061), 
        .Y(n9339) );
  AO21X1_LVT U10662 ( .A1(n4067), .A2(csr_io_evec[4]), .A3(n9339), .Y(
        io_imem_req_bits_pc[4]) );
  AO22X1_LVT U10663 ( .A1(n4064), .A2(csr_io_pc[5]), .A3(n9340), .A4(n4061), 
        .Y(n9341) );
  AO21X1_LVT U10664 ( .A1(n4067), .A2(csr_io_evec[5]), .A3(n9341), .Y(
        io_imem_req_bits_pc[5]) );
  AO22X1_LVT U10665 ( .A1(n4064), .A2(csr_io_pc[6]), .A3(n9342), .A4(n4061), 
        .Y(n9343) );
  AO21X1_LVT U10666 ( .A1(n4067), .A2(csr_io_evec[6]), .A3(n9343), .Y(
        io_imem_req_bits_pc[6]) );
  AO22X1_LVT U10667 ( .A1(n4064), .A2(csr_io_pc[7]), .A3(n9344), .A4(n4061), 
        .Y(n9345) );
  AO21X1_LVT U10668 ( .A1(n4067), .A2(csr_io_evec[7]), .A3(n9345), .Y(
        io_imem_req_bits_pc[7]) );
  AO22X1_LVT U10669 ( .A1(n4064), .A2(csr_io_pc[8]), .A3(n9346), .A4(n4061), 
        .Y(n9347) );
  AO21X1_LVT U10670 ( .A1(n4067), .A2(csr_io_evec[8]), .A3(n9347), .Y(
        io_imem_req_bits_pc[8]) );
  AO22X1_LVT U10671 ( .A1(n4064), .A2(csr_io_pc[9]), .A3(n9348), .A4(n4061), 
        .Y(n9349) );
  AO21X1_LVT U10672 ( .A1(n4067), .A2(csr_io_evec[9]), .A3(n9349), .Y(
        io_imem_req_bits_pc[9]) );
  INVX1_LVT U10673 ( .A(n9509), .Y(n9350) );
  AO222X1_LVT U10674 ( .A1(n4065), .A2(csr_io_evec[10]), .A3(n4064), .A4(
        csr_io_pc[10]), .A5(n9350), .A6(n4059), .Y(io_imem_req_bits_pc[10]) );
  INVX1_LVT U10675 ( .A(n9490), .Y(n9351) );
  AO222X1_LVT U10676 ( .A1(n4065), .A2(csr_io_evec[11]), .A3(n4064), .A4(
        csr_io_pc[11]), .A5(n9351), .A6(n4059), .Y(io_imem_req_bits_pc[11]) );
  INVX1_LVT U10677 ( .A(n9491), .Y(n9352) );
  AO222X1_LVT U10678 ( .A1(n4065), .A2(csr_io_evec[12]), .A3(n4064), .A4(
        csr_io_pc[12]), .A5(n9352), .A6(n4059), .Y(io_imem_req_bits_pc[12]) );
  INVX1_LVT U10679 ( .A(n9500), .Y(n9353) );
  AO222X1_LVT U10680 ( .A1(n4065), .A2(csr_io_evec[13]), .A3(n4064), .A4(
        csr_io_pc[13]), .A5(n9353), .A6(n4059), .Y(io_imem_req_bits_pc[13]) );
  INVX1_LVT U10681 ( .A(n9506), .Y(n9354) );
  AO222X1_LVT U10682 ( .A1(n4065), .A2(csr_io_evec[14]), .A3(n4064), .A4(
        csr_io_pc[14]), .A5(n9354), .A6(n4059), .Y(io_imem_req_bits_pc[14]) );
  AO222X1_LVT U10683 ( .A1(n4065), .A2(csr_io_evec[15]), .A3(n4064), .A4(
        csr_io_pc[15]), .A5(n9355), .A6(n4059), .Y(io_imem_req_bits_pc[15]) );
  AO222X1_LVT U10684 ( .A1(n4065), .A2(csr_io_evec[16]), .A3(n4063), .A4(
        csr_io_pc[16]), .A5(n9356), .A6(n4059), .Y(io_imem_req_bits_pc[16]) );
  INVX1_LVT U10685 ( .A(n9487), .Y(n9357) );
  AO222X1_LVT U10686 ( .A1(n4065), .A2(csr_io_evec[17]), .A3(n4063), .A4(
        csr_io_pc[17]), .A5(n9357), .A6(n4059), .Y(io_imem_req_bits_pc[17]) );
  INVX1_LVT U10687 ( .A(n9496), .Y(n9358) );
  AO222X1_LVT U10688 ( .A1(n4065), .A2(csr_io_evec[18]), .A3(n4063), .A4(
        csr_io_pc[18]), .A5(n9358), .A6(n4059), .Y(io_imem_req_bits_pc[18]) );
  INVX1_LVT U10689 ( .A(n9510), .Y(n9359) );
  AO222X1_LVT U10690 ( .A1(n4065), .A2(csr_io_evec[19]), .A3(n4063), .A4(
        csr_io_pc[19]), .A5(n9359), .A6(n4059), .Y(io_imem_req_bits_pc[19]) );
  INVX1_LVT U10691 ( .A(n9486), .Y(n9360) );
  AO222X1_LVT U10692 ( .A1(n4066), .A2(csr_io_evec[20]), .A3(n4063), .A4(
        csr_io_pc[20]), .A5(n9360), .A6(n4059), .Y(io_imem_req_bits_pc[20]) );
  AO222X1_LVT U10693 ( .A1(n4066), .A2(csr_io_evec[21]), .A3(n4063), .A4(
        csr_io_pc[21]), .A5(n9361), .A6(n4059), .Y(io_imem_req_bits_pc[21]) );
  INVX1_LVT U10694 ( .A(n9501), .Y(n9362) );
  AO222X1_LVT U10695 ( .A1(n4066), .A2(csr_io_evec[22]), .A3(n4063), .A4(
        csr_io_pc[22]), .A5(n9362), .A6(n4060), .Y(io_imem_req_bits_pc[22]) );
  INVX1_LVT U10696 ( .A(n9488), .Y(n9363) );
  AO222X1_LVT U10697 ( .A1(n4066), .A2(csr_io_evec[23]), .A3(n4063), .A4(
        csr_io_pc[23]), .A5(n9363), .A6(n4060), .Y(io_imem_req_bits_pc[23]) );
  AO222X1_LVT U10698 ( .A1(n4066), .A2(csr_io_evec[24]), .A3(n4063), .A4(
        csr_io_pc[24]), .A5(n9364), .A6(n4060), .Y(io_imem_req_bits_pc[24]) );
  INVX1_LVT U10699 ( .A(n9497), .Y(n9365) );
  AO222X1_LVT U10700 ( .A1(n4066), .A2(csr_io_evec[25]), .A3(n4063), .A4(
        csr_io_pc[25]), .A5(n9365), .A6(n4060), .Y(io_imem_req_bits_pc[25]) );
  INVX1_LVT U10701 ( .A(n9483), .Y(n9366) );
  AO222X1_LVT U10702 ( .A1(n4066), .A2(csr_io_evec[26]), .A3(n4063), .A4(
        csr_io_pc[26]), .A5(n9366), .A6(n4060), .Y(io_imem_req_bits_pc[26]) );
  INVX1_LVT U10703 ( .A(n9489), .Y(n9367) );
  AO222X1_LVT U10704 ( .A1(n4066), .A2(csr_io_evec[27]), .A3(n4063), .A4(
        csr_io_pc[27]), .A5(n9367), .A6(n4060), .Y(io_imem_req_bits_pc[27]) );
  AO222X1_LVT U10705 ( .A1(n4066), .A2(csr_io_evec[28]), .A3(n4062), .A4(
        csr_io_pc[28]), .A5(n9368), .A6(n4060), .Y(io_imem_req_bits_pc[28]) );
  INVX1_LVT U10706 ( .A(n9504), .Y(n9369) );
  AO222X1_LVT U10707 ( .A1(n4066), .A2(csr_io_evec[29]), .A3(n4062), .A4(
        csr_io_pc[29]), .A5(n9369), .A6(n4060), .Y(io_imem_req_bits_pc[29]) );
  INVX1_LVT U10708 ( .A(n9502), .Y(n9370) );
  AO222X1_LVT U10709 ( .A1(n4066), .A2(csr_io_evec[31]), .A3(n4062), .A4(
        csr_io_pc[31]), .A5(n9370), .A6(n4060), .Y(io_imem_req_bits_pc[31]) );
  INVX1_LVT U10710 ( .A(n9505), .Y(n9371) );
  AO222X1_LVT U10711 ( .A1(n4066), .A2(csr_io_evec[32]), .A3(n4062), .A4(
        csr_io_pc[32]), .A5(n9371), .A6(n4060), .Y(io_imem_req_bits_pc[32]) );
  INVX1_LVT U10712 ( .A(n9493), .Y(n9372) );
  AO222X1_LVT U10713 ( .A1(n4066), .A2(csr_io_evec[33]), .A3(n4062), .A4(
        csr_io_pc[33]), .A5(n9372), .A6(n4061), .Y(io_imem_req_bits_pc[33]) );
  AO222X1_LVT U10714 ( .A1(n4066), .A2(csr_io_evec[35]), .A3(n4062), .A4(
        csr_io_pc[35]), .A5(n9374), .A6(n4061), .Y(io_imem_req_bits_pc[35]) );
  INVX1_LVT U10715 ( .A(n9494), .Y(n9375) );
  AO222X1_LVT U10716 ( .A1(n4066), .A2(csr_io_evec[37]), .A3(n4062), .A4(
        csr_io_pc[37]), .A5(n9375), .A6(n4061), .Y(io_imem_req_bits_pc[37]) );
  INVX1_LVT U10717 ( .A(n9498), .Y(n9376) );
  AO222X1_LVT U10718 ( .A1(n4065), .A2(csr_io_evec[38]), .A3(n4062), .A4(
        csr_io_pc[38]), .A5(n9376), .A6(n4061), .Y(io_imem_req_bits_pc[38]) );
  OR2X1_LVT U10719 ( .A1(reset), .A2(n9379), .Y(N778) );
  AND3X1_LVT U10720 ( .A1(ex_ctrl_mem), .A2(N290), .A3(ex_ctrl_rxs2), .Y(N526)
         );
  NAND2X0_LVT U10721 ( .A1(n9417), .A2(n1822), .Y(n9384) );
  NAND2X0_LVT U10722 ( .A1(n9385), .A2(n9384), .Y(n_T_760) );
  AND2X1_LVT U10723 ( .A1(n9389), .A2(n2133), .Y(n9404) );
  AND2X1_LVT U10724 ( .A1(n9394), .A2(n9404), .Y(N238) );
  AND2X1_LVT U10725 ( .A1(n9394), .A2(n9405), .Y(N239) );
  AND2X1_LVT U10726 ( .A1(n9389), .A2(n9392), .Y(n9406) );
  AND2X1_LVT U10727 ( .A1(n9394), .A2(n9406), .Y(N240) );
  AND2X1_LVT U10728 ( .A1(n3042), .A2(n2574), .Y(n9391) );
  AND2X1_LVT U10729 ( .A1(n9391), .A2(n2133), .Y(n9407) );
  AND2X1_LVT U10730 ( .A1(n9394), .A2(n9407), .Y(N241) );
  AND2X1_LVT U10731 ( .A1(n9393), .A2(n2133), .Y(n9408) );
  AND2X1_LVT U10732 ( .A1(n9394), .A2(n9408), .Y(N242) );
  AND2X1_LVT U10733 ( .A1(n9391), .A2(n9392), .Y(n9409) );
  AND2X1_LVT U10734 ( .A1(n9394), .A2(n9409), .Y(N243) );
  AND2X1_LVT U10735 ( .A1(n9393), .A2(n9392), .Y(n9411) );
  AND2X1_LVT U10736 ( .A1(n9394), .A2(n9411), .Y(N244) );
  AND2X1_LVT U10737 ( .A1(n9396), .A2(n2150), .Y(N245) );
  AND2X1_LVT U10738 ( .A1(n9404), .A2(n9396), .Y(N246) );
  AND2X1_LVT U10739 ( .A1(n9405), .A2(n9396), .Y(N247) );
  AND2X1_LVT U10740 ( .A1(n9406), .A2(n9396), .Y(N248) );
  AND2X1_LVT U10741 ( .A1(n9407), .A2(n9396), .Y(N249) );
  AND2X1_LVT U10742 ( .A1(n9408), .A2(n9396), .Y(N250) );
  AND2X1_LVT U10743 ( .A1(n9409), .A2(n9396), .Y(N251) );
  AND2X1_LVT U10744 ( .A1(n9411), .A2(n9396), .Y(N252) );
  AND2X1_LVT U10745 ( .A1(n9401), .A2(n2150), .Y(N253) );
  AND2X1_LVT U10746 ( .A1(n9404), .A2(n9401), .Y(N254) );
  AND2X1_LVT U10747 ( .A1(n9401), .A2(n9405), .Y(N255) );
  AND2X1_LVT U10748 ( .A1(n9406), .A2(n9401), .Y(N256) );
  AND2X1_LVT U10749 ( .A1(n9407), .A2(n9401), .Y(N257) );
  AND2X1_LVT U10750 ( .A1(n9408), .A2(n9401), .Y(N258) );
  AND2X1_LVT U10751 ( .A1(n9409), .A2(n9401), .Y(N259) );
  AND2X1_LVT U10752 ( .A1(n9411), .A2(n9401), .Y(N260) );
  AND2X1_LVT U10753 ( .A1(n9410), .A2(n2150), .Y(N261) );
  AND2X1_LVT U10754 ( .A1(n9404), .A2(n9410), .Y(N262) );
  AND2X1_LVT U10755 ( .A1(n9410), .A2(n9405), .Y(N263) );
  AND2X1_LVT U10756 ( .A1(n9406), .A2(n9410), .Y(N264) );
  AND2X1_LVT U10757 ( .A1(n9407), .A2(n9410), .Y(N265) );
  AND2X1_LVT U10758 ( .A1(n9408), .A2(n9410), .Y(N266) );
  AND2X1_LVT U10759 ( .A1(n9409), .A2(n9410), .Y(N267) );
  AND2X1_LVT U10760 ( .A1(n9411), .A2(n9410), .Y(N268) );
  NAND2X0_LVT U10761 ( .A1(n9426), .A2(n9449), .Y(N271) );
  AOI22X1_LVT U10764 ( .A1(n_T_698[14]), .A2(n9506), .A3(n_T_698[8]), .A4(
        n9511), .Y(n9450) );
  AOI22X1_LVT U10765 ( .A1(n_T_698[12]), .A2(n9491), .A3(n_T_698[29]), .A4(
        n9504), .Y(n9451) );
  AOI22X1_LVT U10766 ( .A1(n_T_698[32]), .A2(n9505), .A3(n_T_698[27]), .A4(
        n9489), .Y(n9452) );
  AOI22X1_LVT U10767 ( .A1(n_T_698[6]), .A2(n9485), .A3(n_T_698[9]), .A4(n9507), .Y(n9453) );
  NAND4X0_LVT U10768 ( .A1(n_T_918[59]), .A2(n_T_918[48]), .A3(n_T_918[62]), 
        .A4(n_T_918[56]), .Y(n9469) );
  AND4X1_LVT U10769 ( .A1(n_T_918[39]), .A2(n_T_918[40]), .A3(n_T_918[47]), 
        .A4(n_T_918[60]), .Y(n9459) );
  NAND4X0_LVT U10770 ( .A1(n_T_918[55]), .A2(n_T_918[58]), .A3(n_T_918[44]), 
        .A4(n_T_918[43]), .Y(n9457) );
  NAND4X0_LVT U10771 ( .A1(n_T_918[49]), .A2(n_T_918[45]), .A3(n_T_918[61]), 
        .A4(n_T_918[57]), .Y(n9456) );
  NAND4X0_LVT U10772 ( .A1(n_T_918[41]), .A2(n_T_918[53]), .A3(n_T_918[54]), 
        .A4(n_T_918[50]), .Y(n9455) );
  NAND4X0_LVT U10773 ( .A1(n_T_918[63]), .A2(n_T_918[46]), .A3(n_T_918[42]), 
        .A4(n_T_918[52]), .Y(n9454) );
  NAND3X0_LVT U10774 ( .A1(n_T_918[51]), .A2(n9459), .A3(n9458), .Y(n9468) );
  NAND4X0_LVT U10775 ( .A1(n9463), .A2(n9462), .A3(n9461), .A4(n9460), .Y(
        n9467) );
  NAND3X0_LVT U10776 ( .A1(n9465), .A2(n9464), .A3(n3249), .Y(n9466) );
  OA22X1_LVT U10777 ( .A1(n9469), .A2(n9468), .A3(n9467), .A4(n9466), .Y(n9470) );
  AOI22X1_LVT U10778 ( .A1(n_T_698[3]), .A2(n9503), .A3(n_T_698[18]), .A4(
        n9496), .Y(n9471) );
  AOI22X1_LVT U10779 ( .A1(n_T_698[10]), .A2(n9509), .A3(n_T_698[13]), .A4(
        n9500), .Y(n9472) );
  OAI22X1_LVT U10780 ( .A1(n_T_698[38]), .A2(n9498), .A3(n_T_698[36]), .A4(
        n9508), .Y(n9473) );
  AO221X1_LVT U10781 ( .A1(n9498), .A2(n_T_698[38]), .A3(n_T_698[36]), .A4(
        n9508), .A5(n9473), .Y(n9482) );
  AOI22X1_LVT U10782 ( .A1(n_T_698[33]), .A2(n9493), .A3(n_T_698[5]), .A4(
        n9484), .Y(n9474) );
  OA221X1_LVT U10783 ( .A1(n_T_698[33]), .A2(n9493), .A3(n_T_698[5]), .A4(
        n9484), .A5(n9474), .Y(n9481) );
  AOI22X1_LVT U10784 ( .A1(n_T_698[37]), .A2(n9494), .A3(n_T_698[30]), .A4(
        n9492), .Y(n9475) );
  OA221X1_LVT U10785 ( .A1(n_T_698[37]), .A2(n9494), .A3(n_T_698[30]), .A4(
        n9492), .A5(n9475), .Y(n9480) );
  AOI22X1_LVT U10786 ( .A1(n_T_698[26]), .A2(n9483), .A3(n_T_698[20]), .A4(
        n9486), .Y(n9476) );
  OA221X1_LVT U10787 ( .A1(n_T_698[26]), .A2(n9483), .A3(n_T_698[20]), .A4(
        n9486), .A5(n9476), .Y(n9479) );
  AOI22X1_LVT U10788 ( .A1(n_T_698[11]), .A2(n9490), .A3(n_T_698[17]), .A4(
        n9487), .Y(n9477) );
  OA221X1_LVT U10789 ( .A1(n_T_698[11]), .A2(n9490), .A3(n_T_698[17]), .A4(
        n9487), .A5(n9477), .Y(n9478) );
  NAND2X0_LVT U10790 ( .A1(n555), .A2(n3104), .Y(n9514) );
  AND2X1_LVT U10791 ( .A1(n3202), .A2(n9514), .Y(
        io_imem_btb_update_bits_cfiType[0]) );
  AO22X1_LVT U10792 ( .A1(n_T_849[11]), .A2(n9514), .A3(n_T_904[3]), .A4(n9513), .Y(io_imem_btb_update_bits_cfiType[1]) );
  OR2X1_LVT U10793 ( .A1(io_imem_bht_update_bits_branch), .A2(n9514), .Y(
        io_imem_btb_update_bits_isValid) );
  AND3X1_LVT ibuf_U231 ( .A1(ibuf_n120), .A2(ibuf_n121), .A3(n1822), .Y(
        io_imem_resp_ready) );
  NAND3X0_LVT ibuf_U230 ( .A1(ibuf_n119), .A2(ibuf_n118), .A3(ibuf_n117), .Y(
        ibuf_n120) );
  AND2X1_LVT ibuf_U229 ( .A1(ibuf_n112), .A2(ibuf_n111), .Y(
        ibuf_io_inst_0_valid) );
  NAND2X0_LVT ibuf_U228 ( .A1(ibuf_n110), .A2(ibuf_n12), .Y(ibuf_n111) );
  MUX21X1_LVT ibuf_U227 ( .A1(ibuf_buf__xcpt_pf_inst), .A2(
        io_imem_resp_bits_xcpt_pf_inst), .S0(ibuf_n12), .Y(n_T_728[1]) );
  MUX21X1_LVT ibuf_U226 ( .A1(ibuf_buf__xcpt_ae_inst), .A2(
        io_imem_resp_bits_xcpt_ae_inst), .S0(ibuf_n12), .Y(n_T_728[0]) );
  AND2X1_LVT ibuf_U225 ( .A1(io_imem_resp_bits_xcpt_pf_inst), .A2(ibuf_n122), 
        .Y(n_T_726[1]) );
  AND2X1_LVT ibuf_U224 ( .A1(io_imem_resp_bits_xcpt_ae_inst), .A2(ibuf_n122), 
        .Y(n_T_726[0]) );
  NAND2X0_LVT ibuf_U223 ( .A1(ibuf_n109), .A2(ibuf_n108), .Y(
        ibuf_io_inst_0_bits_replay) );
  NAND4X0_LVT ibuf_U222 ( .A1(ibuf_n113), .A2(io_imem_resp_valid), .A3(
        io_imem_resp_bits_replay), .A4(ibuf_n107), .Y(ibuf_n109) );
  MUX21X1_LVT ibuf_U221 ( .A1(io_imem_resp_bits_data[3]), .A2(
        io_imem_resp_bits_data[19]), .S0(ibuf_n29), .Y(
        ibuf_io_inst_0_bits_raw[19]) );
  MUX21X1_LVT ibuf_U220 ( .A1(io_imem_resp_bits_data[2]), .A2(
        io_imem_resp_bits_data[18]), .S0(ibuf_n23), .Y(
        ibuf_io_inst_0_bits_raw[18]) );
  MUX21X1_LVT ibuf_U219 ( .A1(io_imem_resp_bits_data[0]), .A2(
        io_imem_resp_bits_data[16]), .S0(ibuf_n29), .Y(
        ibuf_io_inst_0_bits_raw[16]) );
  NAND2X0_LVT ibuf_U218 ( .A1(ibuf_n34), .A2(ibuf_buf__data[15]), .Y(ibuf_n104) );
  NAND2X0_LVT ibuf_U217 ( .A1(ibuf_n101), .A2(ibuf_n20), .Y(ibuf_n103) );
  NAND2X0_LVT ibuf_U216 ( .A1(ibuf_buf__data[14]), .A2(ibuf_n34), .Y(ibuf_n99)
         );
  NAND2X0_LVT ibuf_U215 ( .A1(io_imem_resp_bits_data[28]), .A2(ibuf_n18), .Y(
        ibuf_n93) );
  NAND2X0_LVT ibuf_U214 ( .A1(ibuf_buf__data[12]), .A2(ibuf_n34), .Y(ibuf_n94)
         );
  NAND2X0_LVT ibuf_U213 ( .A1(io_imem_resp_bits_data[12]), .A2(ibuf_n28), .Y(
        ibuf_n95) );
  NAND2X0_LVT ibuf_U212 ( .A1(io_imem_resp_bits_data[27]), .A2(ibuf_n115), .Y(
        ibuf_n90) );
  NAND2X0_LVT ibuf_U211 ( .A1(ibuf_buf__data[11]), .A2(ibuf_n34), .Y(ibuf_n91)
         );
  NAND2X0_LVT ibuf_U210 ( .A1(io_imem_resp_bits_data[26]), .A2(ibuf_n18), .Y(
        ibuf_n87) );
  NAND2X0_LVT ibuf_U209 ( .A1(ibuf_buf__data[10]), .A2(ibuf_n34), .Y(ibuf_n88)
         );
  NAND2X0_LVT ibuf_U208 ( .A1(io_imem_resp_bits_data[25]), .A2(ibuf_n115), .Y(
        ibuf_n84) );
  NAND2X0_LVT ibuf_U207 ( .A1(ibuf_buf__data[9]), .A2(ibuf_n34), .Y(ibuf_n85)
         );
  NAND2X0_LVT ibuf_U206 ( .A1(io_imem_resp_bits_data[9]), .A2(ibuf_n28), .Y(
        ibuf_n86) );
  NAND2X0_LVT ibuf_U205 ( .A1(io_imem_resp_bits_data[24]), .A2(ibuf_n18), .Y(
        ibuf_n81) );
  NAND2X0_LVT ibuf_U204 ( .A1(ibuf_buf__data[8]), .A2(ibuf_n34), .Y(ibuf_n82)
         );
  NAND2X0_LVT ibuf_U203 ( .A1(ibuf_n5), .A2(ibuf_n114), .Y(ibuf_n83) );
  NAND2X0_LVT ibuf_U202 ( .A1(io_imem_resp_bits_data[23]), .A2(ibuf_n115), .Y(
        ibuf_n78) );
  NAND2X0_LVT ibuf_U201 ( .A1(ibuf_buf__data[7]), .A2(ibuf_n34), .Y(ibuf_n79)
         );
  NAND2X0_LVT ibuf_U200 ( .A1(io_imem_resp_bits_data[22]), .A2(ibuf_n115), .Y(
        ibuf_n75) );
  NAND2X0_LVT ibuf_U199 ( .A1(ibuf_buf__data[6]), .A2(ibuf_n34), .Y(ibuf_n76)
         );
  NAND2X0_LVT ibuf_U198 ( .A1(io_imem_resp_bits_data[21]), .A2(ibuf_n18), .Y(
        ibuf_n72) );
  NAND2X0_LVT ibuf_U197 ( .A1(ibuf_buf__data[5]), .A2(ibuf_n34), .Y(ibuf_n73)
         );
  NAND2X0_LVT ibuf_U196 ( .A1(ibuf_n28), .A2(io_imem_resp_bits_data[5]), .Y(
        ibuf_n74) );
  NAND2X0_LVT ibuf_U195 ( .A1(io_imem_resp_bits_data[20]), .A2(ibuf_n115), .Y(
        ibuf_n69) );
  NAND2X0_LVT ibuf_U194 ( .A1(ibuf_n34), .A2(ibuf_buf__data[4]), .Y(ibuf_n70)
         );
  NAND2X0_LVT ibuf_U193 ( .A1(io_imem_resp_bits_data[19]), .A2(ibuf_n18), .Y(
        ibuf_n66) );
  NAND2X0_LVT ibuf_U192 ( .A1(ibuf_buf__data[3]), .A2(ibuf_n34), .Y(ibuf_n67)
         );
  NAND2X0_LVT ibuf_U191 ( .A1(io_imem_resp_bits_data[3]), .A2(ibuf_n28), .Y(
        ibuf_n68) );
  NAND3X0_LVT ibuf_U190 ( .A1(ibuf_n65), .A2(ibuf_n64), .A3(ibuf_n63), .Y(
        ibuf_io_inst_0_bits_raw[2]) );
  NAND2X0_LVT ibuf_U189 ( .A1(io_imem_resp_bits_data[18]), .A2(ibuf_n115), .Y(
        ibuf_n63) );
  NAND2X0_LVT ibuf_U188 ( .A1(ibuf_buf__data[2]), .A2(ibuf_n34), .Y(ibuf_n64)
         );
  NAND2X0_LVT ibuf_U187 ( .A1(io_imem_resp_bits_data[2]), .A2(ibuf_n28), .Y(
        ibuf_n65) );
  NAND2X0_LVT ibuf_U186 ( .A1(ibuf_n117), .A2(ibuf_n19), .Y(ibuf_n55) );
  OA21X1_LVT ibuf_U185 ( .A1(ibuf_n54), .A2(ibuf_n34), .A3(ibuf_n121), .Y(
        ibuf_n119) );
  NOR2X0_LVT ibuf_U184 ( .A1(ibuf_n53), .A2(io_imem_req_valid), .Y(ibuf_n40)
         );
  AO21X1_LVT ibuf_U183 ( .A1(ibuf_n51), .A2(ibuf_n52), .A3(reset), .Y(ibuf_n53) );
  AND3X1_LVT ibuf_U182 ( .A1(ibuf_n50), .A2(io_imem_resp_valid), .A3(n1822), 
        .Y(ibuf_N51) );
  MUX21X1_LVT ibuf_U181 ( .A1(ibuf_n49), .A2(ibuf_n48), .S0(ibuf_n116), .Y(
        ibuf_n50) );
  AND2X1_LVT ibuf_U180 ( .A1(ibuf_n107), .A2(ibuf_n117), .Y(ibuf_n48) );
  OR2X1_LVT ibuf_U179 ( .A1(ibuf_n34), .A2(ibuf_io_inst_0_bits_rvc), .Y(
        ibuf_n47) );
  OA21X1_LVT ibuf_U178 ( .A1(ibuf_n12), .A2(n1822), .A3(ibuf_n121), .Y(
        ibuf_n52) );
  OR2X1_LVT ibuf_U177 ( .A1(ibuf_n12), .A2(ibuf_n112), .Y(ibuf_n121) );
  OR2X1_LVT ibuf_U176 ( .A1(ibuf_n46), .A2(ibuf_io_inst_0_bits_rvc), .Y(
        ibuf_n112) );
  NAND2X0_LVT ibuf_U175 ( .A1(ibuf_n54), .A2(ibuf_n108), .Y(ibuf_n46) );
  NAND2X0_LVT ibuf_U174 ( .A1(ibuf_n34), .A2(ibuf_buf__replay), .Y(ibuf_n108)
         );
  AO21X1_LVT ibuf_U173 ( .A1(ibuf_n12), .A2(ibuf_n116), .A3(ibuf_n110), .Y(
        ibuf_n54) );
  NAND2X0_LVT ibuf_U172 ( .A1(io_imem_resp_valid), .A2(ibuf_n107), .Y(
        ibuf_n110) );
  NAND3X0_LVT ibuf_U171 ( .A1(ibuf_n45), .A2(io_imem_resp_bits_btb_taken), 
        .A3(ibuf_n19), .Y(ibuf_n107) );
  NAND2X0_LVT ibuf_U170 ( .A1(ibuf_buf__data[0]), .A2(ibuf_n34), .Y(ibuf_n59)
         );
  NAND3X0_LVT ibuf_U169 ( .A1(ibuf_n58), .A2(ibuf_n59), .A3(ibuf_n57), .Y(
        ibuf_n131) );
  NAND2X0_LVT ibuf_U168 ( .A1(ibuf_buf__data[1]), .A2(ibuf_n34), .Y(ibuf_n62)
         );
  NAND3X0_LVT ibuf_U167 ( .A1(ibuf_n102), .A2(ibuf_n12), .A3(ibuf_n103), .Y(
        ibuf_n105) );
  NAND2X4_LVT ibuf_U166 ( .A1(ibuf_io_inst_0_bits_rvc), .A2(ibuf_n34), .Y(
        ibuf_n113) );
  INVX1_LVT ibuf_U165 ( .A(ibuf_n34), .Y(ibuf_n36) );
  MUX21X1_LVT ibuf_U164 ( .A1(ibuf_n19), .A2(ibuf_n117), .S0(ibuf_n119), .Y(
        ibuf_n56) );
  XOR2X1_LVT ibuf_U163 ( .A1(ibuf_n117), .A2(ibuf_n25), .Y(ibuf_n_T_27_0_) );
  MUX21X1_LVT ibuf_U162 ( .A1(ibuf_ibufBTBResp_bht_history[6]), .A2(
        io_imem_resp_bits_btb_bht_history[6]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[6]) );
  MUX21X1_LVT ibuf_U161 ( .A1(ibuf_ibufBTBResp_bht_history[3]), .A2(
        io_imem_resp_bits_btb_bht_history[3]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[3]) );
  MUX21X1_LVT ibuf_U160 ( .A1(ibuf_ibufBTBResp_bht_history[5]), .A2(
        io_imem_resp_bits_btb_bht_history[5]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[5]) );
  MUX21X1_LVT ibuf_U159 ( .A1(ibuf_ibufBTBResp_entry[4]), .A2(
        io_imem_resp_bits_btb_entry[4]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_entry[4]) );
  MUX21X1_LVT ibuf_U158 ( .A1(ibuf_ibufBTBResp_bht_history[0]), .A2(
        io_imem_resp_bits_btb_bht_history[0]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[0]) );
  MUX21X1_LVT ibuf_U157 ( .A1(ibuf_ibufBTBResp_bht_history[4]), .A2(
        io_imem_resp_bits_btb_bht_history[4]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[4]) );
  MUX21X1_LVT ibuf_U156 ( .A1(ibuf_ibufBTBResp_bht_history[2]), .A2(
        io_imem_resp_bits_btb_bht_history[2]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[2]) );
  MUX21X1_LVT ibuf_U155 ( .A1(ibuf_ibufBTBResp_entry[3]), .A2(
        io_imem_resp_bits_btb_entry[3]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_entry[3]) );
  MUX21X1_LVT ibuf_U154 ( .A1(ibuf_ibufBTBResp_entry[2]), .A2(
        io_imem_resp_bits_btb_entry[2]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_entry[2]) );
  MUX21X1_LVT ibuf_U153 ( .A1(ibuf_ibufBTBResp_bht_history[1]), .A2(
        io_imem_resp_bits_btb_bht_history[1]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[1]) );
  MUX21X1_LVT ibuf_U152 ( .A1(ibuf_ibufBTBResp_entry[0]), .A2(
        io_imem_resp_bits_btb_entry[0]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_entry[0]) );
  MUX21X1_LVT ibuf_U151 ( .A1(ibuf_ibufBTBResp_entry[1]), .A2(
        io_imem_resp_bits_btb_entry[1]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_entry[1]) );
  MUX21X1_LVT ibuf_U150 ( .A1(ibuf_ibufBTBResp_bht_history[7]), .A2(
        io_imem_resp_bits_btb_bht_history[7]), .S0(ibuf_n113), .Y(
        ibuf_io_btb_resp_bht_history[7]) );
  NAND3X0_LVT ibuf_U149 ( .A1(ibuf_n68), .A2(ibuf_n67), .A3(ibuf_n66), .Y(
        ibuf_n129) );
  MUX21X1_LVT ibuf_U148 ( .A1(io_imem_resp_bits_data[9]), .A2(
        io_imem_resp_bits_data[25]), .S0(ibuf_n29), .Y(
        ibuf_io_inst_0_bits_raw[25]) );
  MUX21X1_LVT ibuf_U147 ( .A1(ibuf_buf__pc[3]), .A2(io_imem_resp_bits_pc[3]), 
        .S0(ibuf_n12), .Y(ibuf_io_pc[3]) );
  MUX21X1_LVT ibuf_U146 ( .A1(ibuf_buf__pc[0]), .A2(io_imem_resp_bits_pc[0]), 
        .S0(ibuf_n12), .Y(ibuf_io_pc[0]) );
  MUX21X1_LVT ibuf_U145 ( .A1(ibuf_buf__pc[2]), .A2(io_imem_resp_bits_pc[2]), 
        .S0(ibuf_n12), .Y(ibuf_io_pc[2]) );
  MUX21X1_LVT ibuf_U144 ( .A1(io_imem_resp_bits_data[13]), .A2(
        io_imem_resp_bits_data[29]), .S0(ibuf_n100), .Y(ibuf_n_T_34[13]) );
  MUX21X1_LVT ibuf_U143 ( .A1(io_imem_resp_bits_data[0]), .A2(
        io_imem_resp_bits_data[16]), .S0(ibuf_n100), .Y(ibuf_n_T_34[0]) );
  MUX21X1_LVT ibuf_U142 ( .A1(io_imem_resp_bits_data[10]), .A2(
        io_imem_resp_bits_data[26]), .S0(ibuf_n100), .Y(ibuf_n_T_34[10]) );
  MUX21X1_LVT ibuf_U141 ( .A1(io_imem_resp_bits_data[9]), .A2(
        io_imem_resp_bits_data[25]), .S0(ibuf_n100), .Y(ibuf_n_T_34[9]) );
  MUX21X1_LVT ibuf_U140 ( .A1(io_imem_resp_bits_data[4]), .A2(
        io_imem_resp_bits_data[20]), .S0(ibuf_n100), .Y(ibuf_n_T_34[4]) );
  MUX21X1_LVT ibuf_U139 ( .A1(io_imem_resp_bits_data[8]), .A2(
        io_imem_resp_bits_data[24]), .S0(ibuf_n100), .Y(ibuf_n_T_34[8]) );
  MUX21X1_LVT ibuf_U138 ( .A1(io_imem_resp_bits_data[11]), .A2(
        io_imem_resp_bits_data[27]), .S0(ibuf_n100), .Y(ibuf_n_T_34[11]) );
  MUX21X1_LVT ibuf_U137 ( .A1(io_imem_resp_bits_data[2]), .A2(
        io_imem_resp_bits_data[18]), .S0(ibuf_n100), .Y(ibuf_n_T_34[2]) );
  MUX21X1_LVT ibuf_U136 ( .A1(io_imem_resp_bits_data[14]), .A2(
        io_imem_resp_bits_data[30]), .S0(ibuf_n100), .Y(ibuf_n_T_34[14]) );
  MUX21X1_LVT ibuf_U135 ( .A1(io_imem_resp_bits_data[7]), .A2(
        io_imem_resp_bits_data[23]), .S0(ibuf_n100), .Y(ibuf_n_T_34[7]) );
  MUX21X1_LVT ibuf_U134 ( .A1(io_imem_resp_bits_data[1]), .A2(
        io_imem_resp_bits_data[17]), .S0(ibuf_n100), .Y(ibuf_n_T_34[1]) );
  MUX21X1_LVT ibuf_U133 ( .A1(io_imem_resp_bits_data[6]), .A2(
        io_imem_resp_bits_data[22]), .S0(ibuf_n100), .Y(ibuf_n_T_34[6]) );
  MUX21X1_LVT ibuf_U132 ( .A1(io_imem_resp_bits_data[15]), .A2(
        io_imem_resp_bits_data[31]), .S0(ibuf_n100), .Y(ibuf_n_T_34[15]) );
  MUX21X1_LVT ibuf_U131 ( .A1(io_imem_resp_bits_data[3]), .A2(
        io_imem_resp_bits_data[19]), .S0(ibuf_n100), .Y(ibuf_n_T_34[3]) );
  MUX21X1_LVT ibuf_U130 ( .A1(io_imem_resp_bits_data[12]), .A2(
        io_imem_resp_bits_data[28]), .S0(ibuf_n100), .Y(ibuf_n_T_34[12]) );
  MUX21X1_LVT ibuf_U129 ( .A1(io_imem_resp_bits_data[5]), .A2(
        io_imem_resp_bits_data[21]), .S0(ibuf_n100), .Y(ibuf_n_T_34[5]) );
  NBUFFX2_LVT ibuf_U128 ( .A(ibuf_net35341), .Y(ibuf_n37) );
  NBUFFX2_LVT ibuf_U127 ( .A(ibuf_net35341), .Y(ibuf_n38) );
  NBUFFX2_LVT ibuf_U126 ( .A(ibuf_net35341), .Y(ibuf_n39) );
  NBUFFX2_LVT ibuf_U125 ( .A(ibuf_net35341), .Y(ibuf_n41) );
  NBUFFX2_LVT ibuf_U124 ( .A(ibuf_net35341), .Y(ibuf_n42) );
  NBUFFX2_LVT ibuf_U123 ( .A(ibuf_net35341), .Y(ibuf_n43) );
  IBUFFX2_LVT ibuf_U122 ( .A(io_imem_resp_bits_pc[1]), .Y(ibuf_n114) );
  INVX1_LVT ibuf_U121 ( .A(io_imem_resp_bits_data[13]), .Y(ibuf_n35) );
  INVX1_LVT ibuf_U120 ( .A(io_imem_resp_bits_data[29]), .Y(ibuf_n96) );
  AO21X2_LVT ibuf_U119 ( .A1(ibuf_buf__pc[1]), .A2(ibuf_n34), .A3(ibuf_n18), 
        .Y(ibuf_io_pc[1]) );
  AND2X1_LVT ibuf_U118 ( .A1(ibuf_n85), .A2(ibuf_n84), .Y(ibuf_n33) );
  NAND2X0_LVT ibuf_U117 ( .A1(ibuf_n12), .A2(io_imem_resp_bits_pc[1]), .Y(
        ibuf_n32) );
  NAND2X0_LVT ibuf_U116 ( .A1(ibuf_n31), .A2(ibuf_n114), .Y(ibuf_n80) );
  NAND2X0_LVT ibuf_U115 ( .A1(ibuf_n25), .A2(ibuf_n30), .Y(ibuf_n89) );
  MUX21X1_LVT ibuf_U114 ( .A1(io_imem_resp_bits_data[5]), .A2(
        io_imem_resp_bits_data[21]), .S0(ibuf_n11), .Y(ibuf_n_T_55_85_) );
  MUX21X1_LVT ibuf_U113 ( .A1(io_imem_resp_bits_data[8]), .A2(
        io_imem_resp_bits_data[24]), .S0(ibuf_n11), .Y(
        ibuf_io_inst_0_bits_raw[24]) );
  MUX21X1_LVT ibuf_U112 ( .A1(io_imem_resp_bits_data[7]), .A2(
        io_imem_resp_bits_data[23]), .S0(ibuf_n10), .Y(
        ibuf_io_inst_0_bits_raw[23]) );
  MUX21X1_LVT ibuf_U111 ( .A1(io_imem_resp_bits_data[6]), .A2(
        io_imem_resp_bits_data[22]), .S0(ibuf_n10), .Y(
        ibuf_io_inst_0_bits_raw[22]) );
  MUX21X1_LVT ibuf_U110 ( .A1(io_imem_resp_bits_data[10]), .A2(
        io_imem_resp_bits_data[26]), .S0(ibuf_n29), .Y(
        ibuf_io_inst_0_bits_raw[26]) );
  MUX21X1_LVT ibuf_U109 ( .A1(io_imem_resp_bits_data[1]), .A2(
        io_imem_resp_bits_data[17]), .S0(ibuf_n29), .Y(
        ibuf_io_inst_0_bits_raw[17]) );
  NBUFFX2_LVT ibuf_U108 ( .A(ibuf_n11), .Y(ibuf_n29) );
  NAND2X0_LVT ibuf_U107 ( .A1(ibuf_n27), .A2(ibuf_n114), .Y(ibuf_n92) );
  NAND2X0_LVT ibuf_U106 ( .A1(ibuf_n25), .A2(ibuf_n26), .Y(ibuf_n77) );
  NAND3X0_LVT ibuf_U105 ( .A1(ibuf_n62), .A2(ibuf_n61), .A3(ibuf_n60), .Y(
        ibuf_n130) );
  NBUFFX2_LVT ibuf_U104 ( .A(ibuf_n114), .Y(ibuf_n25) );
  NAND2X0_LVT ibuf_U103 ( .A1(ibuf_n24), .A2(ibuf_n114), .Y(ibuf_n71) );
  INVX1_LVT ibuf_U102 ( .A(ibuf_n32), .Y(ibuf_n115) );
  NBUFFX2_LVT ibuf_U101 ( .A(ibuf_n10), .Y(ibuf_n23) );
  NBUFFX2_LVT ibuf_U100 ( .A(ibuf_n127), .Y(ibuf_io_inst_0_bits_raw[10]) );
  AND2X1_LVT ibuf_U99 ( .A1(ibuf_n114), .A2(ibuf_n12), .Y(ibuf_n28) );
  MUX21X1_LVT ibuf_U98 ( .A1(io_imem_resp_bits_data[11]), .A2(
        io_imem_resp_bits_data[27]), .S0(ibuf_n11), .Y(ibuf_n_T_55_91_) );
  NBUFFX2_LVT ibuf_U97 ( .A(ibuf_n_T_55_91_), .Y(ibuf_io_inst_0_bits_raw[27])
         );
  NAND2X0_LVT ibuf_U96 ( .A1(ibuf_n33), .A2(ibuf_n86), .Y(
        ibuf_io_inst_0_bits_raw[9]) );
  NBUFFX2_LVT ibuf_U95 ( .A(io_imem_resp_bits_pc[1]), .Y(ibuf_n20) );
  AO21X1_LVT ibuf_U94 ( .A1(io_imem_resp_bits_btb_taken), .A2(ibuf_n45), .A3(
        ibuf_n19), .Y(ibuf_n116) );
  OR2X1_LVT ibuf_U93 ( .A1(ibuf_n20), .A2(io_imem_resp_bits_data[15]), .Y(
        ibuf_n102) );
  NAND3X0_LVT ibuf_U92 ( .A1(ibuf_n12), .A2(ibuf_n20), .A3(
        io_imem_resp_bits_data[16]), .Y(ibuf_n57) );
  IBUFFX2_LVT ibuf_U91 ( .A(io_imem_resp_bits_data[31]), .Y(ibuf_n101) );
  INVX1_LVT ibuf_U90 ( .A(ibuf_n32), .Y(ibuf_n18) );
  NBUFFX2_LVT ibuf_U89 ( .A(ibuf_n125), .Y(ibuf_io_inst_0_bits_raw[13]) );
  NAND3X0_LVT ibuf_U88 ( .A1(ibuf_n62), .A2(ibuf_n61), .A3(ibuf_n60), .Y(
        ibuf_io_inst_0_bits_raw[1]) );
  NBUFFX2_LVT ibuf_U87 ( .A(ibuf_n_T_55_85_), .Y(ibuf_io_inst_0_bits_raw[21])
         );
  NAND3X0_LVT ibuf_U86 ( .A1(ibuf_n98), .A2(ibuf_n99), .A3(ibuf_n97), .Y(
        ibuf_n124) );
  INVX0_LVT ibuf_U85 ( .A(io_imem_resp_bits_btb_bridx), .Y(ibuf_n45) );
  INVX0_LVT ibuf_U84 ( .A(ibuf_n25), .Y(ibuf_n19) );
  INVX0_LVT ibuf_U83 ( .A(ibuf_n116), .Y(ibuf_n118) );
  MUX21X1_LVT ibuf_U82 ( .A1(io_imem_resp_bits_data[14]), .A2(
        io_imem_resp_bits_data[30]), .S0(ibuf_n11), .Y(
        ibuf_io_inst_0_bits_raw[30]) );
  MUX21X1_LVT ibuf_U81 ( .A1(io_imem_resp_bits_data[13]), .A2(
        io_imem_resp_bits_data[29]), .S0(ibuf_n23), .Y(
        ibuf_io_inst_0_bits_raw[29]) );
  NAND3X0_LVT ibuf_U80 ( .A1(ibuf_n69), .A2(ibuf_n70), .A3(ibuf_n71), .Y(
        ibuf_io_inst_0_bits_raw[4]) );
  NAND3X0_LVT ibuf_U79 ( .A1(ibuf_n74), .A2(ibuf_n73), .A3(ibuf_n72), .Y(
        ibuf_io_inst_0_bits_raw[5]) );
  NAND3X0_LVT ibuf_U78 ( .A1(ibuf_n77), .A2(ibuf_n76), .A3(ibuf_n75), .Y(
        ibuf_n128) );
  NAND3X0_LVT ibuf_U77 ( .A1(ibuf_n80), .A2(ibuf_n79), .A3(ibuf_n78), .Y(
        ibuf_io_inst_0_bits_raw[7]) );
  NAND2X0_LVT ibuf_U76 ( .A1(ibuf_n47), .A2(ibuf_n113), .Y(ibuf_n117) );
  INVX0_LVT ibuf_U75 ( .A(ibuf_n117), .Y(ibuf_n49) );
  INVX0_LVT ibuf_U74 ( .A(ibuf_N51), .Y(ibuf_n51) );
  INVX1_LVT ibuf_U73 ( .A(ibuf_n122), .Y(ibuf_io_inst_0_bits_rvc) );
  NAND2X0_LVT ibuf_U72 ( .A1(ibuf_n56), .A2(ibuf_n55), .Y(ibuf_n100) );
  NAND3X0_LVT ibuf_U71 ( .A1(ibuf_n90), .A2(ibuf_n91), .A3(ibuf_n92), .Y(
        ibuf_io_inst_0_bits_raw[11]) );
  NAND3X1_LVT ibuf_U70 ( .A1(ibuf_n114), .A2(ibuf_n12), .A3(
        io_imem_resp_bits_data[1]), .Y(ibuf_n61) );
  NBUFFX2_LVT ibuf_U69 ( .A(ibuf_n123), .Y(ibuf_io_inst_0_bits_raw[15]) );
  MUX21X2_LVT ibuf_U68 ( .A1(io_imem_resp_bits_data[12]), .A2(
        io_imem_resp_bits_data[28]), .S0(ibuf_n10), .Y(
        ibuf_io_inst_0_bits_raw[28]) );
  NAND3X0_LVT ibuf_U67 ( .A1(ibuf_n95), .A2(ibuf_n94), .A3(ibuf_n93), .Y(
        ibuf_n126) );
  NAND3X0_LVT ibuf_U66 ( .A1(ibuf_n95), .A2(ibuf_n94), .A3(ibuf_n93), .Y(
        ibuf_io_inst_0_bits_raw[12]) );
  NAND3X2_LVT ibuf_U65 ( .A1(ibuf_n89), .A2(ibuf_n88), .A3(ibuf_n87), .Y(
        ibuf_n127) );
  NAND3X1_LVT ibuf_U64 ( .A1(ibuf_n12), .A2(ibuf_n20), .A3(
        io_imem_resp_bits_data[17]), .Y(ibuf_n60) );
  MUX21X2_LVT ibuf_U63 ( .A1(io_imem_resp_bits_data[15]), .A2(
        io_imem_resp_bits_data[31]), .S0(ibuf_n106), .Y(n2576) );
  OR2X1_LVT ibuf_U62 ( .A1(ibuf_n20), .A2(ibuf_n12), .Y(ibuf_n106) );
  OR2X2_LVT ibuf_U61 ( .A1(ibuf_n20), .A2(ibuf_n12), .Y(ibuf_n11) );
  OR2X2_LVT ibuf_U60 ( .A1(ibuf_n20), .A2(ibuf_n12), .Y(ibuf_n10) );
  NAND2X4_LVT ibuf_U59 ( .A1(ibuf_n105), .A2(ibuf_n104), .Y(ibuf_n123) );
  AO22X2_LVT ibuf_U58 ( .A1(ibuf_buf__data[13]), .A2(ibuf_n34), .A3(ibuf_n8), 
        .A4(ibuf_n9), .Y(ibuf_n125) );
  NAND2X0_LVT ibuf_U57 ( .A1(ibuf_n20), .A2(ibuf_n96), .Y(ibuf_n9) );
  AND2X1_LVT ibuf_U56 ( .A1(ibuf_n12), .A2(ibuf_n7), .Y(ibuf_n8) );
  NAND2X0_LVT ibuf_U55 ( .A1(ibuf_n35), .A2(ibuf_n114), .Y(ibuf_n7) );
  MUX21X1_LVT ibuf_U54 ( .A1(ibuf_buf__pc[4]), .A2(io_imem_resp_bits_pc[4]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[4]) );
  MUX21X1_LVT ibuf_U53 ( .A1(ibuf_buf__pc[5]), .A2(io_imem_resp_bits_pc[5]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[5]) );
  MUX21X1_LVT ibuf_U52 ( .A1(ibuf_buf__pc[6]), .A2(io_imem_resp_bits_pc[6]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[6]) );
  MUX21X1_LVT ibuf_U51 ( .A1(ibuf_buf__pc[7]), .A2(io_imem_resp_bits_pc[7]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[7]) );
  MUX21X1_LVT ibuf_U50 ( .A1(ibuf_buf__pc[8]), .A2(io_imem_resp_bits_pc[8]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[8]) );
  MUX21X1_LVT ibuf_U49 ( .A1(ibuf_buf__pc[9]), .A2(io_imem_resp_bits_pc[9]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[9]) );
  MUX21X1_LVT ibuf_U48 ( .A1(ibuf_buf__pc[10]), .A2(io_imem_resp_bits_pc[10]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[10]) );
  MUX21X1_LVT ibuf_U47 ( .A1(ibuf_buf__pc[11]), .A2(io_imem_resp_bits_pc[11]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[11]) );
  MUX21X1_LVT ibuf_U46 ( .A1(ibuf_buf__pc[12]), .A2(io_imem_resp_bits_pc[12]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[12]) );
  MUX21X1_LVT ibuf_U45 ( .A1(ibuf_buf__pc[13]), .A2(io_imem_resp_bits_pc[13]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[13]) );
  MUX21X1_LVT ibuf_U44 ( .A1(ibuf_buf__pc[14]), .A2(io_imem_resp_bits_pc[14]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[14]) );
  MUX21X1_LVT ibuf_U43 ( .A1(ibuf_buf__pc[15]), .A2(io_imem_resp_bits_pc[15]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[15]) );
  MUX21X1_LVT ibuf_U42 ( .A1(ibuf_buf__pc[16]), .A2(io_imem_resp_bits_pc[16]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[16]) );
  MUX21X1_LVT ibuf_U41 ( .A1(ibuf_buf__pc[17]), .A2(io_imem_resp_bits_pc[17]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[17]) );
  MUX21X1_LVT ibuf_U40 ( .A1(ibuf_buf__pc[18]), .A2(io_imem_resp_bits_pc[18]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[18]) );
  MUX21X1_LVT ibuf_U39 ( .A1(ibuf_buf__pc[19]), .A2(io_imem_resp_bits_pc[19]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[19]) );
  MUX21X1_LVT ibuf_U38 ( .A1(ibuf_buf__pc[20]), .A2(io_imem_resp_bits_pc[20]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[20]) );
  MUX21X1_LVT ibuf_U37 ( .A1(ibuf_buf__pc[21]), .A2(io_imem_resp_bits_pc[21]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[21]) );
  MUX21X1_LVT ibuf_U36 ( .A1(ibuf_buf__pc[22]), .A2(io_imem_resp_bits_pc[22]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[22]) );
  MUX21X1_LVT ibuf_U35 ( .A1(ibuf_buf__pc[23]), .A2(io_imem_resp_bits_pc[23]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[23]) );
  MUX21X1_LVT ibuf_U34 ( .A1(ibuf_buf__pc[24]), .A2(io_imem_resp_bits_pc[24]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[24]) );
  MUX21X1_LVT ibuf_U33 ( .A1(ibuf_buf__pc[25]), .A2(io_imem_resp_bits_pc[25]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[25]) );
  MUX21X1_LVT ibuf_U32 ( .A1(ibuf_buf__pc[26]), .A2(io_imem_resp_bits_pc[26]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[26]) );
  MUX21X1_LVT ibuf_U31 ( .A1(ibuf_buf__pc[27]), .A2(io_imem_resp_bits_pc[27]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[27]) );
  MUX21X1_LVT ibuf_U30 ( .A1(ibuf_buf__pc[28]), .A2(io_imem_resp_bits_pc[28]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[28]) );
  MUX21X1_LVT ibuf_U29 ( .A1(ibuf_buf__pc[29]), .A2(io_imem_resp_bits_pc[29]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[29]) );
  MUX21X1_LVT ibuf_U28 ( .A1(ibuf_buf__pc[30]), .A2(io_imem_resp_bits_pc[30]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[30]) );
  MUX21X1_LVT ibuf_U27 ( .A1(ibuf_buf__pc[31]), .A2(io_imem_resp_bits_pc[31]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[31]) );
  MUX21X1_LVT ibuf_U26 ( .A1(ibuf_buf__pc[32]), .A2(io_imem_resp_bits_pc[32]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[32]) );
  MUX21X1_LVT ibuf_U25 ( .A1(ibuf_buf__pc[33]), .A2(io_imem_resp_bits_pc[33]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[33]) );
  MUX21X1_LVT ibuf_U24 ( .A1(ibuf_buf__pc[34]), .A2(io_imem_resp_bits_pc[34]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[34]) );
  MUX21X1_LVT ibuf_U23 ( .A1(ibuf_buf__pc[35]), .A2(io_imem_resp_bits_pc[35]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[35]) );
  MUX21X1_LVT ibuf_U22 ( .A1(ibuf_buf__pc[36]), .A2(io_imem_resp_bits_pc[36]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[36]) );
  MUX21X1_LVT ibuf_U21 ( .A1(ibuf_buf__pc[37]), .A2(io_imem_resp_bits_pc[37]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[37]) );
  MUX21X1_LVT ibuf_U20 ( .A1(ibuf_buf__pc[38]), .A2(io_imem_resp_bits_pc[38]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[38]) );
  MUX21X1_LVT ibuf_U19 ( .A1(ibuf_buf__pc[39]), .A2(io_imem_resp_bits_pc[39]), 
        .S0(ibuf_n36), .Y(ibuf_io_pc[39]) );
  AND2X1_LVT ibuf_U18 ( .A1(ibuf_n12), .A2(io_imem_resp_bits_data[4]), .Y(
        ibuf_n24) );
  AND2X1_LVT ibuf_U17 ( .A1(ibuf_n12), .A2(io_imem_resp_bits_data[6]), .Y(
        ibuf_n26) );
  AND2X1_LVT ibuf_U16 ( .A1(ibuf_n12), .A2(io_imem_resp_bits_data[7]), .Y(
        ibuf_n31) );
  AND2X1_LVT ibuf_U15 ( .A1(ibuf_n12), .A2(io_imem_resp_bits_data[10]), .Y(
        ibuf_n30) );
  AND2X1_LVT ibuf_U14 ( .A1(ibuf_n12), .A2(io_imem_resp_bits_data[11]), .Y(
        ibuf_n27) );
  NAND3X0_LVT ibuf_U13 ( .A1(ibuf_n12), .A2(ibuf_n20), .A3(
        io_imem_resp_bits_data[30]), .Y(ibuf_n97) );
  NAND3X2_LVT ibuf_U12 ( .A1(ibuf_n83), .A2(ibuf_n82), .A3(ibuf_n81), .Y(
        ibuf_io_inst_0_bits_raw[8]) );
  NAND3X0_LVT ibuf_U11 ( .A1(ibuf_n58), .A2(ibuf_n59), .A3(ibuf_n57), .Y(
        ibuf_io_inst_0_bits_raw[0]) );
  AND2X1_LVT ibuf_U10 ( .A1(io_imem_resp_bits_data[8]), .A2(ibuf_n12), .Y(
        ibuf_n5) );
  NAND3X0_LVT ibuf_U9 ( .A1(ibuf_n98), .A2(ibuf_n99), .A3(ibuf_n97), .Y(
        ibuf_io_inst_0_bits_raw[14]) );
  NAND3X1_LVT ibuf_U8 ( .A1(ibuf_n114), .A2(ibuf_n36), .A3(
        io_imem_resp_bits_data[0]), .Y(ibuf_n58) );
  NAND3X1_LVT ibuf_U7 ( .A1(ibuf_n114), .A2(ibuf_n12), .A3(
        io_imem_resp_bits_data[14]), .Y(ibuf_n98) );
  NAND3X2_LVT ibuf_U6 ( .A1(ibuf_n77), .A2(ibuf_n76), .A3(ibuf_n75), .Y(
        ibuf_io_inst_0_bits_raw[6]) );
  NAND3X0_LVT ibuf_U5 ( .A1(ibuf_n68), .A2(ibuf_n67), .A3(ibuf_n66), .Y(
        ibuf_io_inst_0_bits_raw[3]) );
  MUX21X1_LVT ibuf_U4 ( .A1(io_imem_resp_bits_data[4]), .A2(
        io_imem_resp_bits_data[20]), .S0(ibuf_n23), .Y(ibuf_n_T_55_84_) );
  MUX21X2_LVT ibuf_U3 ( .A1(io_imem_resp_bits_data[4]), .A2(
        io_imem_resp_bits_data[20]), .S0(ibuf_n23), .Y(
        ibuf_io_inst_0_bits_raw[20]) );
  DFFX2_LVT ibuf_nBufValid_reg ( .D(ibuf_n40), .CLK(n3595), .Q(ibuf_n34), .QN(
        ibuf_n12) );
  DFFX1_LVT ibuf_buf__xcpt_ae_inst_reg ( .D(io_imem_resp_bits_xcpt_ae_inst), 
        .CLK(ibuf_n37), .Q(ibuf_buf__xcpt_ae_inst) );
  DFFX1_LVT ibuf_buf__xcpt_pf_inst_reg ( .D(io_imem_resp_bits_xcpt_pf_inst), 
        .CLK(ibuf_n37), .Q(ibuf_buf__xcpt_pf_inst) );
  DFFX1_LVT ibuf_buf__data_reg_1_ ( .D(ibuf_n_T_34[1]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[1]) );
  DFFX1_LVT ibuf_buf__data_reg_2_ ( .D(ibuf_n_T_34[2]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[2]) );
  DFFX1_LVT ibuf_buf__data_reg_3_ ( .D(ibuf_n_T_34[3]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[3]) );
  DFFX1_LVT ibuf_buf__data_reg_4_ ( .D(ibuf_n_T_34[4]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[4]) );
  DFFX1_LVT ibuf_buf__data_reg_5_ ( .D(ibuf_n_T_34[5]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[5]) );
  DFFX1_LVT ibuf_buf__data_reg_6_ ( .D(ibuf_n_T_34[6]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[6]) );
  DFFX1_LVT ibuf_buf__data_reg_7_ ( .D(ibuf_n_T_34[7]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[7]) );
  DFFX1_LVT ibuf_buf__data_reg_8_ ( .D(ibuf_n_T_34[8]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[8]) );
  DFFX1_LVT ibuf_buf__data_reg_9_ ( .D(ibuf_n_T_34[9]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[9]) );
  DFFX1_LVT ibuf_buf__data_reg_10_ ( .D(ibuf_n_T_34[10]), .CLK(ibuf_n37), .Q(
        ibuf_buf__data[10]) );
  DFFX1_LVT ibuf_buf__data_reg_11_ ( .D(ibuf_n_T_34[11]), .CLK(ibuf_n38), .Q(
        ibuf_buf__data[11]) );
  DFFX1_LVT ibuf_buf__data_reg_12_ ( .D(ibuf_n_T_34[12]), .CLK(ibuf_n38), .Q(
        ibuf_buf__data[12]) );
  DFFX1_LVT ibuf_buf__data_reg_13_ ( .D(ibuf_n_T_34[13]), .CLK(ibuf_n38), .Q(
        ibuf_buf__data[13]) );
  DFFX1_LVT ibuf_buf__data_reg_14_ ( .D(ibuf_n_T_34[14]), .CLK(ibuf_n38), .Q(
        ibuf_buf__data[14]) );
  DFFX1_LVT ibuf_buf__data_reg_15_ ( .D(ibuf_n_T_34[15]), .CLK(ibuf_n38), .Q(
        ibuf_buf__data[15]) );
  DFFX1_LVT ibuf_buf__pc_reg_0_ ( .D(io_imem_resp_bits_pc[0]), .CLK(ibuf_n38), 
        .Q(ibuf_buf__pc[0]) );
  DFFX1_LVT ibuf_buf__pc_reg_1_ ( .D(ibuf_n_T_27_0_), .CLK(ibuf_n38), .Q(
        ibuf_buf__pc[1]) );
  DFFX1_LVT ibuf_buf__pc_reg_2_ ( .D(io_imem_resp_bits_pc[2]), .CLK(ibuf_n38), 
        .Q(ibuf_buf__pc[2]) );
  DFFX1_LVT ibuf_buf__pc_reg_3_ ( .D(io_imem_resp_bits_pc[3]), .CLK(ibuf_n38), 
        .Q(ibuf_buf__pc[3]) );
  DFFX1_LVT ibuf_buf__pc_reg_4_ ( .D(io_imem_resp_bits_pc[4]), .CLK(ibuf_n38), 
        .Q(ibuf_buf__pc[4]) );
  DFFX1_LVT ibuf_buf__pc_reg_5_ ( .D(io_imem_resp_bits_pc[5]), .CLK(ibuf_n38), 
        .Q(ibuf_buf__pc[5]) );
  DFFX1_LVT ibuf_buf__pc_reg_6_ ( .D(io_imem_resp_bits_pc[6]), .CLK(ibuf_n38), 
        .Q(ibuf_buf__pc[6]) );
  DFFX1_LVT ibuf_buf__pc_reg_7_ ( .D(io_imem_resp_bits_pc[7]), .CLK(ibuf_n39), 
        .Q(ibuf_buf__pc[7]) );
  DFFX1_LVT ibuf_buf__pc_reg_8_ ( .D(io_imem_resp_bits_pc[8]), .CLK(ibuf_n39), 
        .Q(ibuf_buf__pc[8]) );
  DFFX1_LVT ibuf_buf__pc_reg_9_ ( .D(io_imem_resp_bits_pc[9]), .CLK(ibuf_n39), 
        .Q(ibuf_buf__pc[9]) );
  DFFX1_LVT ibuf_buf__pc_reg_10_ ( .D(io_imem_resp_bits_pc[10]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[10]) );
  DFFX1_LVT ibuf_buf__pc_reg_11_ ( .D(io_imem_resp_bits_pc[11]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[11]) );
  DFFX1_LVT ibuf_buf__pc_reg_12_ ( .D(io_imem_resp_bits_pc[12]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[12]) );
  DFFX1_LVT ibuf_buf__pc_reg_13_ ( .D(io_imem_resp_bits_pc[13]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[13]) );
  DFFX1_LVT ibuf_buf__pc_reg_14_ ( .D(io_imem_resp_bits_pc[14]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[14]) );
  DFFX1_LVT ibuf_buf__pc_reg_15_ ( .D(io_imem_resp_bits_pc[15]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[15]) );
  DFFX1_LVT ibuf_buf__pc_reg_16_ ( .D(io_imem_resp_bits_pc[16]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[16]) );
  DFFX1_LVT ibuf_buf__pc_reg_17_ ( .D(io_imem_resp_bits_pc[17]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[17]) );
  DFFX1_LVT ibuf_buf__pc_reg_18_ ( .D(io_imem_resp_bits_pc[18]), .CLK(ibuf_n39), .Q(ibuf_buf__pc[18]) );
  DFFX1_LVT ibuf_buf__pc_reg_19_ ( .D(io_imem_resp_bits_pc[19]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[19]) );
  DFFX1_LVT ibuf_buf__pc_reg_20_ ( .D(io_imem_resp_bits_pc[20]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[20]) );
  DFFX1_LVT ibuf_buf__pc_reg_21_ ( .D(io_imem_resp_bits_pc[21]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[21]) );
  DFFX1_LVT ibuf_buf__pc_reg_22_ ( .D(io_imem_resp_bits_pc[22]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[22]) );
  DFFX1_LVT ibuf_buf__pc_reg_23_ ( .D(io_imem_resp_bits_pc[23]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[23]) );
  DFFX1_LVT ibuf_buf__pc_reg_24_ ( .D(io_imem_resp_bits_pc[24]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[24]) );
  DFFX1_LVT ibuf_buf__pc_reg_25_ ( .D(io_imem_resp_bits_pc[25]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[25]) );
  DFFX1_LVT ibuf_buf__pc_reg_26_ ( .D(io_imem_resp_bits_pc[26]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[26]) );
  DFFX1_LVT ibuf_buf__pc_reg_27_ ( .D(io_imem_resp_bits_pc[27]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[27]) );
  DFFX1_LVT ibuf_buf__pc_reg_28_ ( .D(io_imem_resp_bits_pc[28]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[28]) );
  DFFX1_LVT ibuf_buf__pc_reg_29_ ( .D(io_imem_resp_bits_pc[29]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[29]) );
  DFFX1_LVT ibuf_buf__pc_reg_30_ ( .D(io_imem_resp_bits_pc[30]), .CLK(ibuf_n41), .Q(ibuf_buf__pc[30]) );
  DFFX1_LVT ibuf_buf__pc_reg_31_ ( .D(io_imem_resp_bits_pc[31]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[31]) );
  DFFX1_LVT ibuf_buf__pc_reg_32_ ( .D(io_imem_resp_bits_pc[32]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[32]) );
  DFFX1_LVT ibuf_buf__pc_reg_33_ ( .D(io_imem_resp_bits_pc[33]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[33]) );
  DFFX1_LVT ibuf_buf__pc_reg_34_ ( .D(io_imem_resp_bits_pc[34]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[34]) );
  DFFX1_LVT ibuf_buf__pc_reg_35_ ( .D(io_imem_resp_bits_pc[35]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[35]) );
  DFFX1_LVT ibuf_buf__pc_reg_36_ ( .D(io_imem_resp_bits_pc[36]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[36]) );
  DFFX1_LVT ibuf_buf__pc_reg_37_ ( .D(io_imem_resp_bits_pc[37]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[37]) );
  DFFX1_LVT ibuf_buf__pc_reg_38_ ( .D(io_imem_resp_bits_pc[38]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[38]) );
  DFFX1_LVT ibuf_buf__pc_reg_39_ ( .D(io_imem_resp_bits_pc[39]), .CLK(ibuf_n42), .Q(ibuf_buf__pc[39]) );
  DFFX1_LVT ibuf_buf__replay_reg ( .D(io_imem_resp_bits_replay), .CLK(ibuf_n42), .Q(ibuf_buf__replay) );
  DFFX1_LVT ibuf_ibufBTBResp_entry_reg_0_ ( .D(io_imem_resp_bits_btb_entry[0]), 
        .CLK(ibuf_n42), .Q(ibuf_ibufBTBResp_entry[0]) );
  DFFX1_LVT ibuf_ibufBTBResp_entry_reg_1_ ( .D(io_imem_resp_bits_btb_entry[1]), 
        .CLK(ibuf_n42), .Q(ibuf_ibufBTBResp_entry[1]) );
  DFFX1_LVT ibuf_ibufBTBResp_entry_reg_2_ ( .D(io_imem_resp_bits_btb_entry[2]), 
        .CLK(ibuf_n43), .Q(ibuf_ibufBTBResp_entry[2]) );
  DFFX1_LVT ibuf_ibufBTBResp_entry_reg_3_ ( .D(io_imem_resp_bits_btb_entry[3]), 
        .CLK(ibuf_n43), .Q(ibuf_ibufBTBResp_entry[3]) );
  DFFX1_LVT ibuf_ibufBTBResp_entry_reg_4_ ( .D(io_imem_resp_bits_btb_entry[4]), 
        .CLK(ibuf_n43), .Q(ibuf_ibufBTBResp_entry[4]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_0_ ( .D(
        io_imem_resp_bits_btb_bht_history[0]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[0]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_1_ ( .D(
        io_imem_resp_bits_btb_bht_history[1]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[1]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_2_ ( .D(
        io_imem_resp_bits_btb_bht_history[2]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[2]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_3_ ( .D(
        io_imem_resp_bits_btb_bht_history[3]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[3]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_4_ ( .D(
        io_imem_resp_bits_btb_bht_history[4]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[4]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_5_ ( .D(
        io_imem_resp_bits_btb_bht_history[5]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[5]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_6_ ( .D(
        io_imem_resp_bits_btb_bht_history[6]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[6]) );
  DFFX1_LVT ibuf_ibufBTBResp_bht_history_reg_7_ ( .D(
        io_imem_resp_bits_btb_bht_history[7]), .CLK(ibuf_n43), .Q(
        ibuf_ibufBTBResp_bht_history[7]) );
  DFFX1_LVT ibuf_buf__data_reg_0_ ( .D(ibuf_n_T_34[0]), .CLK(ibuf_n43), .Q(
        ibuf_buf__data[0]) );
  SNPS_CLOCK_GATE_HIGH_IBuf ibuf_clk_gate_ibufBTBResp_bht_history_reg ( .CLK(
        n3595), .EN(ibuf_N51), .ENCLK(ibuf_net35341), .TE(1'b0) );
  OA22X1_LVT ibuf_RVCExpander_U395 ( .A1(ibuf_RVCExpander_n40), .A2(
        ibuf_RVCExpander_n351), .A3(ibuf_RVCExpander_n350), .A4(
        ibuf_RVCExpander_n349), .Y(ibuf_RVCExpander_n352) );
  INVX1_LVT ibuf_RVCExpander_U394 ( .A(n2576), .Y(ibuf_RVCExpander_n351) );
  NAND2X0_LVT ibuf_RVCExpander_U393 ( .A1(ibuf_RVCExpander_n342), .A2(
        ibuf_RVCExpander_n341), .Y(ibuf_RVCExpander_n346) );
  NAND3X0_LVT ibuf_RVCExpander_U392 ( .A1(ibuf_RVCExpander_n337), .A2(
        ibuf_n127), .A3(ibuf_RVCExpander_n336), .Y(ibuf_RVCExpander_n338) );
  NAND2X0_LVT ibuf_RVCExpander_U391 ( .A1(ibuf_io_inst_0_bits_raw[29]), .A2(
        ibuf_n122), .Y(ibuf_RVCExpander_n339) );
  AND2X1_LVT ibuf_RVCExpander_U390 ( .A1(ibuf_RVCExpander_n353), .A2(
        ibuf_RVCExpander_n335), .Y(ibuf_RVCExpander_n348) );
  AO21X1_LVT ibuf_RVCExpander_U389 ( .A1(ibuf_RVCExpander_n333), .A2(
        ibuf_RVCExpander_n334), .A3(ibuf_RVCExpander_n350), .Y(
        ibuf_RVCExpander_n353) );
  NAND2X0_LVT ibuf_RVCExpander_U388 ( .A1(ibuf_RVCExpander_n327), .A2(
        ibuf_RVCExpander_n326), .Y(ibuf_RVCExpander_n330) );
  NAND2X0_LVT ibuf_RVCExpander_U387 ( .A1(ibuf_RVCExpander_n66), .A2(
        ibuf_RVCExpander_n337), .Y(ibuf_RVCExpander_n326) );
  NAND2X0_LVT ibuf_RVCExpander_U386 ( .A1(ibuf_RVCExpander_n52), .A2(
        ibuf_RVCExpander_n325), .Y(ibuf_RVCExpander_n327) );
  AND3X1_LVT ibuf_RVCExpander_U385 ( .A1(ibuf_RVCExpander_n324), .A2(
        ibuf_RVCExpander_n323), .A3(ibuf_RVCExpander_n322), .Y(
        ibuf_RVCExpander_n332) );
  NAND2X0_LVT ibuf_RVCExpander_U384 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(
        ibuf_n122), .Y(ibuf_RVCExpander_n322) );
  MUX21X1_LVT ibuf_RVCExpander_U383 ( .A1(ibuf_RVCExpander_n52), .A2(
        ibuf_RVCExpander_n66), .S0(ibuf_n123), .Y(ibuf_RVCExpander_n321) );
  NAND2X0_LVT ibuf_RVCExpander_U382 ( .A1(ibuf_RVCExpander_n70), .A2(
        ibuf_RVCExpander_n319), .Y(ibuf_RVCExpander_n324) );
  AND2X1_LVT ibuf_RVCExpander_U381 ( .A1(ibuf_RVCExpander_n54), .A2(
        ibuf_RVCExpander_n328), .Y(ibuf_RVCExpander_n318) );
  NAND2X0_LVT ibuf_RVCExpander_U380 ( .A1(ibuf_RVCExpander_n313), .A2(
        ibuf_RVCExpander_n312), .Y(ibuf_RVCExpander_n314) );
  AO21X1_LVT ibuf_RVCExpander_U379 ( .A1(ibuf_RVCExpander_n311), .A2(
        ibuf_RVCExpander_n310), .A3(ibuf_RVCExpander_n309), .Y(
        ibuf_RVCExpander_n313) );
  NAND3X0_LVT ibuf_RVCExpander_U378 ( .A1(ibuf_RVCExpander_n308), .A2(
        ibuf_RVCExpander_n307), .A3(ibuf_RVCExpander_n306), .Y(
        ibuf_RVCExpander_n315) );
  NAND2X0_LVT ibuf_RVCExpander_U377 ( .A1(ibuf_RVCExpander_n337), .A2(
        ibuf_io_inst_0_bits_raw[8]), .Y(ibuf_RVCExpander_n306) );
  AND3X1_LVT ibuf_RVCExpander_U376 ( .A1(ibuf_RVCExpander_n305), .A2(
        ibuf_RVCExpander_n312), .A3(ibuf_RVCExpander_n304), .Y(
        ibuf_RVCExpander_n308) );
  NAND2X0_LVT ibuf_RVCExpander_U375 ( .A1(ibuf_RVCExpander_n325), .A2(
        ibuf_RVCExpander_n55), .Y(ibuf_RVCExpander_n304) );
  OA222X1_LVT ibuf_RVCExpander_U374 ( .A1(ibuf_RVCExpander_n40), .A2(
        ibuf_RVCExpander_n303), .A3(ibuf_RVCExpander_n302), .A4(
        ibuf_RVCExpander_n301), .A5(ibuf_RVCExpander_n300), .A6(
        ibuf_RVCExpander_n299), .Y(ibuf_RVCExpander_n312) );
  OA21X1_LVT ibuf_RVCExpander_U373 ( .A1(ibuf_RVCExpander_n298), .A2(
        ibuf_RVCExpander_n297), .A3(ibuf_RVCExpander_n311), .Y(
        ibuf_RVCExpander_n305) );
  NAND2X0_LVT ibuf_RVCExpander_U372 ( .A1(ibuf_RVCExpander_n296), .A2(
        ibuf_RVCExpander_n9), .Y(ibuf_RVCExpander_n311) );
  NAND4X0_LVT ibuf_RVCExpander_U371 ( .A1(ibuf_RVCExpander_n295), .A2(
        ibuf_RVCExpander_n294), .A3(ibuf_RVCExpander_n293), .A4(
        ibuf_RVCExpander_n292), .Y(io_fpu_inst[26]) );
  NAND2X0_LVT ibuf_RVCExpander_U370 ( .A1(ibuf_io_inst_0_bits_raw[26]), .A2(
        ibuf_n122), .Y(ibuf_RVCExpander_n292) );
  NAND2X0_LVT ibuf_RVCExpander_U369 ( .A1(ibuf_RVCExpander_n62), .A2(
        ibuf_RVCExpander_n291), .Y(ibuf_RVCExpander_n293) );
  NAND4X0_LVT ibuf_RVCExpander_U368 ( .A1(ibuf_RVCExpander_n287), .A2(
        ibuf_RVCExpander_n286), .A3(ibuf_RVCExpander_n285), .A4(
        ibuf_RVCExpander_n284), .Y(ibuf_RVCExpander_n295) );
  NAND2X0_LVT ibuf_RVCExpander_U367 ( .A1(ibuf_RVCExpander_n283), .A2(
        ibuf_RVCExpander_n282), .Y(ibuf_RVCExpander_n284) );
  NAND3X0_LVT ibuf_RVCExpander_U366 ( .A1(ibuf_RVCExpander_n307), .A2(
        ibuf_RVCExpander_n282), .A3(ibuf_RVCExpander_n281), .Y(
        ibuf_RVCExpander_n287) );
  NAND2X0_LVT ibuf_RVCExpander_U365 ( .A1(ibuf_RVCExpander_n62), .A2(
        ibuf_RVCExpander_n337), .Y(ibuf_RVCExpander_n281) );
  NAND2X0_LVT ibuf_RVCExpander_U364 ( .A1(ibuf_RVCExpander_n38), .A2(
        ibuf_RVCExpander_n278), .Y(ibuf_RVCExpander_n282) );
  NAND3X0_LVT ibuf_RVCExpander_U363 ( .A1(ibuf_RVCExpander_n277), .A2(
        ibuf_RVCExpander_n68), .A3(ibuf_RVCExpander_n328), .Y(
        ibuf_RVCExpander_n278) );
  OA21X1_LVT ibuf_RVCExpander_U362 ( .A1(ibuf_RVCExpander_n350), .A2(
        ibuf_RVCExpander_n276), .A3(ibuf_RVCExpander_n275), .Y(
        ibuf_RVCExpander_n307) );
  OR3X1_LVT ibuf_RVCExpander_U361 ( .A1(ibuf_RVCExpander_n272), .A2(
        ibuf_RVCExpander_n271), .A3(ibuf_RVCExpander_n309), .Y(
        ibuf_RVCExpander_n273) );
  OR2X1_LVT ibuf_RVCExpander_U360 ( .A1(ibuf_RVCExpander_n350), .A2(
        ibuf_RVCExpander_n296), .Y(ibuf_RVCExpander_n272) );
  AND3X1_LVT ibuf_RVCExpander_U359 ( .A1(ibuf_RVCExpander_n269), .A2(
        ibuf_RVCExpander_n268), .A3(ibuf_RVCExpander_n267), .Y(
        ibuf_RVCExpander_n274) );
  NAND2X0_LVT ibuf_RVCExpander_U358 ( .A1(ibuf_io_inst_0_bits_raw[25]), .A2(
        ibuf_n122), .Y(ibuf_RVCExpander_n267) );
  AO21X1_LVT ibuf_RVCExpander_U357 ( .A1(ibuf_RVCExpander_n266), .A2(
        ibuf_RVCExpander_n277), .A3(ibuf_RVCExpander_n290), .Y(
        ibuf_RVCExpander_n269) );
  AO21X1_LVT ibuf_RVCExpander_U356 ( .A1(ibuf_RVCExpander_n262), .A2(
        ibuf_RVCExpander_n336), .A3(ibuf_RVCExpander_n261), .Y(io_fpu_inst[23]) );
  NAND4X0_LVT ibuf_RVCExpander_U355 ( .A1(ibuf_RVCExpander_n260), .A2(
        ibuf_RVCExpander_n259), .A3(ibuf_RVCExpander_n275), .A4(
        ibuf_RVCExpander_n258), .Y(ibuf_RVCExpander_n262) );
  NAND2X0_LVT ibuf_RVCExpander_U354 ( .A1(ibuf_RVCExpander_n257), .A2(
        ibuf_RVCExpander_n38), .Y(ibuf_RVCExpander_n258) );
  OA21X1_LVT ibuf_RVCExpander_U353 ( .A1(ibuf_RVCExpander_n344), .A2(
        ibuf_RVCExpander_n256), .A3(ibuf_RVCExpander_n255), .Y(
        ibuf_RVCExpander_n259) );
  NAND3X0_LVT ibuf_RVCExpander_U352 ( .A1(ibuf_RVCExpander_n254), .A2(
        ibuf_RVCExpander_n253), .A3(ibuf_RVCExpander_n252), .Y(io_fpu_inst[22]) );
  NAND2X0_LVT ibuf_RVCExpander_U351 ( .A1(ibuf_RVCExpander_n52), .A2(
        ibuf_RVCExpander_n251), .Y(ibuf_RVCExpander_n252) );
  NAND3X0_LVT ibuf_RVCExpander_U350 ( .A1(ibuf_RVCExpander_n250), .A2(
        ibuf_RVCExpander_n317), .A3(ibuf_RVCExpander_n249), .Y(
        ibuf_RVCExpander_n251) );
  OA21X1_LVT ibuf_RVCExpander_U349 ( .A1(ibuf_n125), .A2(ibuf_RVCExpander_n248), .A3(ibuf_RVCExpander_n65), .Y(ibuf_RVCExpander_n249) );
  AND3X1_LVT ibuf_RVCExpander_U348 ( .A1(ibuf_RVCExpander_n247), .A2(
        ibuf_RVCExpander_n275), .A3(ibuf_RVCExpander_n246), .Y(
        ibuf_RVCExpander_n253) );
  OR2X1_LVT ibuf_RVCExpander_U347 ( .A1(ibuf_RVCExpander_n245), .A2(
        ibuf_RVCExpander_n299), .Y(ibuf_RVCExpander_n247) );
  NAND2X0_LVT ibuf_RVCExpander_U346 ( .A1(ibuf_n125), .A2(
        ibuf_RVCExpander_n241), .Y(ibuf_RVCExpander_n297) );
  OA22X1_LVT ibuf_RVCExpander_U345 ( .A1(ibuf_RVCExpander_n240), .A2(
        ibuf_RVCExpander_n263), .A3(ibuf_RVCExpander_n239), .A4(
        ibuf_RVCExpander_n238), .Y(io_fpu_inst[21]) );
  NAND2X0_LVT ibuf_RVCExpander_U344 ( .A1(ibuf_RVCExpander_n275), .A2(
        ibuf_RVCExpander_n250), .Y(ibuf_RVCExpander_n238) );
  NAND4X0_LVT ibuf_RVCExpander_U343 ( .A1(ibuf_RVCExpander_n299), .A2(
        ibuf_RVCExpander_n317), .A3(ibuf_RVCExpander_n65), .A4(
        ibuf_RVCExpander_n237), .Y(ibuf_RVCExpander_n239) );
  INVX1_LVT ibuf_RVCExpander_U342 ( .A(ibuf_RVCExpander_n275), .Y(
        ibuf_RVCExpander_n263) );
  NAND2X0_LVT ibuf_RVCExpander_U341 ( .A1(ibuf_RVCExpander_n237), .A2(
        ibuf_RVCExpander_n301), .Y(ibuf_RVCExpander_n240) );
  NAND3X0_LVT ibuf_RVCExpander_U340 ( .A1(ibuf_RVCExpander_n236), .A2(
        ibuf_RVCExpander_n235), .A3(ibuf_RVCExpander_n234), .Y(io_fpu_inst[20]) );
  OA21X1_LVT ibuf_RVCExpander_U339 ( .A1(ibuf_RVCExpander_n233), .A2(
        ibuf_RVCExpander_n232), .A3(ibuf_RVCExpander_n231), .Y(
        ibuf_RVCExpander_n236) );
  NAND2X0_LVT ibuf_RVCExpander_U338 ( .A1(ibuf_RVCExpander_n1), .A2(
        ibuf_RVCExpander_n230), .Y(ibuf_RVCExpander_n231) );
  NAND3X0_LVT ibuf_RVCExpander_U337 ( .A1(ibuf_RVCExpander_n250), .A2(
        ibuf_RVCExpander_n317), .A3(ibuf_RVCExpander_n299), .Y(
        ibuf_RVCExpander_n230) );
  NAND2X0_LVT ibuf_RVCExpander_U336 ( .A1(ibuf_RVCExpander_n227), .A2(
        ibuf_RVCExpander_n235), .Y(io_fpu_inst[19]) );
  AND2X1_LVT ibuf_RVCExpander_U335 ( .A1(ibuf_RVCExpander_n275), .A2(
        ibuf_RVCExpander_n222), .Y(ibuf_RVCExpander_n235) );
  AND2X1_LVT ibuf_RVCExpander_U334 ( .A1(ibuf_RVCExpander_n220), .A2(
        ibuf_RVCExpander_n219), .Y(io_fpu_inst[16]) );
  NAND3X0_LVT ibuf_RVCExpander_U333 ( .A1(ibuf_RVCExpander_n218), .A2(
        ibuf_RVCExpander_n222), .A3(ibuf_RVCExpander_n217), .Y(
        ibuf_RVCExpander_n219) );
  OA222X1_LVT ibuf_RVCExpander_U332 ( .A1(ibuf_RVCExpander_n298), .A2(
        ibuf_RVCExpander_n53), .A3(ibuf_RVCExpander_n300), .A4(
        ibuf_RVCExpander_n214), .A5(ibuf_RVCExpander_n213), .A6(
        ibuf_RVCExpander_n212), .Y(ibuf_RVCExpander_n215) );
  AND2X1_LVT ibuf_RVCExpander_U331 ( .A1(ibuf_RVCExpander_n211), .A2(
        ibuf_RVCExpander_n277), .Y(ibuf_RVCExpander_n214) );
  NAND3X0_LVT ibuf_RVCExpander_U330 ( .A1(ibuf_RVCExpander_n208), .A2(
        ibuf_RVCExpander_n207), .A3(ibuf_RVCExpander_n206), .Y(
        ibuf_RVCExpander_n220) );
  AO21X1_LVT ibuf_RVCExpander_U329 ( .A1(ibuf_RVCExpander_n205), .A2(
        ibuf_RVCExpander_n328), .A3(ibuf_RVCExpander_n300), .Y(
        ibuf_RVCExpander_n208) );
  AND2X1_LVT ibuf_RVCExpander_U328 ( .A1(ibuf_RVCExpander_n201), .A2(
        ibuf_RVCExpander_n328), .Y(ibuf_RVCExpander_n202) );
  NAND3X0_LVT ibuf_RVCExpander_U327 ( .A1(ibuf_RVCExpander_n270), .A2(
        ibuf_RVCExpander_n196), .A3(ibuf_RVCExpander_n350), .Y(
        ibuf_RVCExpander_n197) );
  NAND2X0_LVT ibuf_RVCExpander_U326 ( .A1(ibuf_RVCExpander_n52), .A2(
        ibuf_RVCExpander_n64), .Y(ibuf_RVCExpander_n198) );
  OR2X1_LVT ibuf_RVCExpander_U325 ( .A1(ibuf_RVCExpander_n195), .A2(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n199) );
  NAND2X0_LVT ibuf_RVCExpander_U324 ( .A1(ibuf_RVCExpander_n63), .A2(
        ibuf_RVCExpander_n341), .Y(ibuf_RVCExpander_n192) );
  AND3X1_LVT ibuf_RVCExpander_U323 ( .A1(ibuf_RVCExpander_n68), .A2(
        ibuf_RVCExpander_n191), .A3(ibuf_RVCExpander_n222), .Y(
        ibuf_RVCExpander_n193) );
  OA21X1_LVT ibuf_RVCExpander_U322 ( .A1(ibuf_RVCExpander_n190), .A2(
        ibuf_RVCExpander_n285), .A3(ibuf_RVCExpander_n189), .Y(
        ibuf_RVCExpander_n191) );
  OR2X1_LVT ibuf_RVCExpander_U321 ( .A1(ibuf_RVCExpander_n216), .A2(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n189) );
  NAND2X0_LVT ibuf_RVCExpander_U320 ( .A1(ibuf_io_inst_0_bits_raw[11]), .A2(
        ibuf_RVCExpander_n187), .Y(ibuf_RVCExpander_n188) );
  AND3X1_LVT ibuf_RVCExpander_U319 ( .A1(ibuf_RVCExpander_n328), .A2(
        ibuf_RVCExpander_n285), .A3(ibuf_RVCExpander_n182), .Y(
        ibuf_RVCExpander_n184) );
  OA21X1_LVT ibuf_RVCExpander_U318 ( .A1(ibuf_RVCExpander_n316), .A2(
        ibuf_RVCExpander_n290), .A3(ibuf_RVCExpander_n181), .Y(
        ibuf_RVCExpander_n186) );
  AND2X1_LVT ibuf_RVCExpander_U317 ( .A1(ibuf_RVCExpander_n222), .A2(
        ibuf_RVCExpander_n343), .Y(ibuf_RVCExpander_n200) );
  NAND2X0_LVT ibuf_RVCExpander_U316 ( .A1(ibuf_RVCExpander_n340), .A2(
        ibuf_RVCExpander_n70), .Y(ibuf_RVCExpander_n222) );
  OAI22X1_LVT ibuf_RVCExpander_U315 ( .A1(ibuf_RVCExpander_n176), .A2(
        ibuf_RVCExpander_n344), .A3(ibuf_RVCExpander_n309), .A4(
        ibuf_RVCExpander_n175), .Y(io_fpu_inst[10]) );
  OR3X1_LVT ibuf_RVCExpander_U314 ( .A1(ibuf_RVCExpander_n174), .A2(
        ibuf_RVCExpander_n47), .A3(ibuf_RVCExpander_n310), .Y(
        ibuf_RVCExpander_n175) );
  NAND2X0_LVT ibuf_RVCExpander_U313 ( .A1(ibuf_RVCExpander_n349), .A2(
        ibuf_RVCExpander_n173), .Y(ibuf_RVCExpander_n310) );
  NAND3X0_LVT ibuf_RVCExpander_U312 ( .A1(ibuf_RVCExpander_n167), .A2(
        ibuf_RVCExpander_n166), .A3(ibuf_RVCExpander_n165), .Y(io_fpu_inst[8])
         );
  NAND2X0_LVT ibuf_RVCExpander_U311 ( .A1(ibuf_RVCExpander_n279), .A2(
        ibuf_io_inst_0_bits_raw[8]), .Y(ibuf_RVCExpander_n166) );
  NAND2X0_LVT ibuf_RVCExpander_U310 ( .A1(ibuf_RVCExpander_n164), .A2(
        ibuf_io_inst_0_bits_raw[8]), .Y(ibuf_RVCExpander_n167) );
  NAND2X0_LVT ibuf_RVCExpander_U309 ( .A1(ibuf_RVCExpander_n169), .A2(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n164) );
  NAND2X0_LVT ibuf_RVCExpander_U308 ( .A1(ibuf_RVCExpander_n283), .A2(
        ibuf_RVCExpander_n70), .Y(ibuf_RVCExpander_n335) );
  NAND2X0_LVT ibuf_RVCExpander_U307 ( .A1(ibuf_RVCExpander_n63), .A2(ibuf_n122), .Y(ibuf_RVCExpander_n159) );
  NAND2X0_LVT ibuf_RVCExpander_U306 ( .A1(ibuf_RVCExpander_n158), .A2(
        ibuf_RVCExpander_n3), .Y(ibuf_RVCExpander_n160) );
  NAND2X0_LVT ibuf_RVCExpander_U305 ( .A1(ibuf_RVCExpander_n8), .A2(
        ibuf_RVCExpander_n172), .Y(ibuf_RVCExpander_n155) );
  OA21X1_LVT ibuf_RVCExpander_U304 ( .A1(ibuf_RVCExpander_n71), .A2(
        ibuf_RVCExpander_n151), .A3(ibuf_RVCExpander_n299), .Y(
        ibuf_RVCExpander_n156) );
  AND2X1_LVT ibuf_RVCExpander_U303 ( .A1(ibuf_RVCExpander_n37), .A2(
        ibuf_RVCExpander_n288), .Y(ibuf_RVCExpander_n299) );
  AND3X1_LVT ibuf_RVCExpander_U302 ( .A1(ibuf_RVCExpander_n170), .A2(
        ibuf_RVCExpander_n266), .A3(ibuf_RVCExpander_n54), .Y(
        ibuf_RVCExpander_n157) );
  NOR2X0_LVT ibuf_RVCExpander_U301 ( .A1(ibuf_RVCExpander_n174), .A2(
        ibuf_RVCExpander_n341), .Y(ibuf_RVCExpander_n260) );
  NAND3X0_LVT ibuf_RVCExpander_U300 ( .A1(ibuf_RVCExpander_n150), .A2(
        ibuf_RVCExpander_n149), .A3(ibuf_RVCExpander_n148), .Y(n9527) );
  NAND2X0_LVT ibuf_RVCExpander_U299 ( .A1(ibuf_RVCExpander_n163), .A2(
        ibuf_RVCExpander_n147), .Y(ibuf_RVCExpander_n148) );
  NAND2X0_LVT ibuf_RVCExpander_U298 ( .A1(ibuf_RVCExpander_n61), .A2(
        ibuf_RVCExpander_n248), .Y(ibuf_RVCExpander_n147) );
  OA21X1_LVT ibuf_RVCExpander_U297 ( .A1(ibuf_RVCExpander_n40), .A2(
        ibuf_RVCExpander_n245), .A3(ibuf_RVCExpander_n170), .Y(
        ibuf_RVCExpander_n149) );
  NAND2X0_LVT ibuf_RVCExpander_U296 ( .A1(ibuf_RVCExpander_n61), .A2(
        ibuf_RVCExpander_n349), .Y(ibuf_RVCExpander_n145) );
  NAND2X0_LVT ibuf_RVCExpander_U295 ( .A1(ibuf_RVCExpander_n302), .A2(
        ibuf_RVCExpander_n67), .Y(ibuf_RVCExpander_n146) );
  NAND2X0_LVT ibuf_RVCExpander_U294 ( .A1(ibuf_n122), .A2(ibuf_RVCExpander_n55), .Y(ibuf_RVCExpander_n142) );
  OR2X1_LVT ibuf_RVCExpander_U293 ( .A1(ibuf_RVCExpander_n233), .A2(
        ibuf_RVCExpander_n141), .Y(ibuf_RVCExpander_n143) );
  NAND3X0_LVT ibuf_RVCExpander_U292 ( .A1(ibuf_RVCExpander_n139), .A2(
        ibuf_RVCExpander_n138), .A3(ibuf_RVCExpander_n137), .Y(
        ibuf_RVCExpander_n140) );
  AO21X1_LVT ibuf_RVCExpander_U291 ( .A1(ibuf_RVCExpander_n135), .A2(
        ibuf_RVCExpander_n136), .A3(ibuf_RVCExpander_n134), .Y(
        ibuf_RVCExpander_n137) );
  NAND3X0_LVT ibuf_RVCExpander_U290 ( .A1(ibuf_RVCExpander_n201), .A2(
        ibuf_RVCExpander_n210), .A3(ibuf_RVCExpander_n177), .Y(
        ibuf_RVCExpander_n134) );
  NAND3X0_LVT ibuf_RVCExpander_U289 ( .A1(ibuf_RVCExpander_n133), .A2(
        ibuf_RVCExpander_n132), .A3(ibuf_RVCExpander_n256), .Y(
        ibuf_RVCExpander_n135) );
  NAND2X0_LVT ibuf_RVCExpander_U288 ( .A1(ibuf_RVCExpander_n190), .A2(
        ibuf_n123), .Y(ibuf_RVCExpander_n136) );
  OA21X1_LVT ibuf_RVCExpander_U287 ( .A1(ibuf_RVCExpander_n211), .A2(
        ibuf_RVCExpander_n216), .A3(ibuf_RVCExpander_n131), .Y(
        ibuf_RVCExpander_n139) );
  NAND2X0_LVT ibuf_RVCExpander_U286 ( .A1(ibuf_RVCExpander_n341), .A2(
        ibuf_RVCExpander_n70), .Y(ibuf_RVCExpander_n131) );
  AND2X1_LVT ibuf_RVCExpander_U285 ( .A1(ibuf_RVCExpander_n270), .A2(
        ibuf_RVCExpander_n179), .Y(ibuf_RVCExpander_n341) );
  INVX1_LVT ibuf_RVCExpander_U284 ( .A(ibuf_RVCExpander_n187), .Y(
        ibuf_RVCExpander_n179) );
  NAND2X0_LVT ibuf_RVCExpander_U283 ( .A1(ibuf_io_inst_0_bits_raw[11]), .A2(
        ibuf_n127), .Y(ibuf_RVCExpander_n187) );
  NAND2X0_LVT ibuf_RVCExpander_U282 ( .A1(ibuf_RVCExpander_n127), .A2(
        ibuf_RVCExpander_n126), .Y(ibuf_RVCExpander_n128) );
  NAND3X0_LVT ibuf_RVCExpander_U281 ( .A1(ibuf_RVCExpander_n125), .A2(
        ibuf_RVCExpander_n124), .A3(ibuf_RVCExpander_n123), .Y(
        ibuf_RVCExpander_n130) );
  NAND3X0_LVT ibuf_RVCExpander_U280 ( .A1(ibuf_RVCExpander_n122), .A2(
        ibuf_RVCExpander_n161), .A3(ibuf_RVCExpander_n195), .Y(
        ibuf_RVCExpander_n123) );
  AND2X1_LVT ibuf_RVCExpander_U279 ( .A1(ibuf_RVCExpander_n300), .A2(
        ibuf_RVCExpander_n350), .Y(ibuf_RVCExpander_n152) );
  NOR2X0_LVT ibuf_RVCExpander_U278 ( .A1(ibuf_n127), .A2(ibuf_RVCExpander_n62), 
        .Y(ibuf_RVCExpander_n154) );
  INVX1_LVT ibuf_RVCExpander_U277 ( .A(ibuf_RVCExpander_n5), .Y(
        ibuf_RVCExpander_n168) );
  AND3X1_LVT ibuf_RVCExpander_U276 ( .A1(ibuf_RVCExpander_n119), .A2(
        ibuf_RVCExpander_n71), .A3(ibuf_RVCExpander_n54), .Y(
        ibuf_RVCExpander_n124) );
  INVX1_LVT ibuf_RVCExpander_U275 ( .A(ibuf_RVCExpander_n117), .Y(
        ibuf_RVCExpander_n118) );
  INVX1_LVT ibuf_RVCExpander_U274 ( .A(ibuf_io_inst_0_bits_raw[7]), .Y(
        ibuf_RVCExpander_n289) );
  NAND2X0_LVT ibuf_RVCExpander_U273 ( .A1(ibuf_RVCExpander_n113), .A2(
        ibuf_RVCExpander_n112), .Y(ibuf_RVCExpander_n173) );
  INVX1_LVT ibuf_RVCExpander_U272 ( .A(ibuf_RVCExpander_n57), .Y(
        ibuf_RVCExpander_n195) );
  AND2X1_LVT ibuf_RVCExpander_U271 ( .A1(ibuf_RVCExpander_n127), .A2(
        ibuf_RVCExpander_n138), .Y(ibuf_RVCExpander_n125) );
  AND2X1_LVT ibuf_RVCExpander_U270 ( .A1(ibuf_RVCExpander_n111), .A2(
        ibuf_RVCExpander_n65), .Y(ibuf_RVCExpander_n138) );
  INVX1_LVT ibuf_RVCExpander_U269 ( .A(ibuf_RVCExpander_n108), .Y(
        ibuf_RVCExpander_n178) );
  NAND3X0_LVT ibuf_RVCExpander_U268 ( .A1(ibuf_RVCExpander_n104), .A2(
        ibuf_RVCExpander_n103), .A3(ibuf_RVCExpander_n170), .Y(
        ibuf_RVCExpander_n105) );
  AND2X1_LVT ibuf_RVCExpander_U267 ( .A1(ibuf_RVCExpander_n288), .A2(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n286) );
  NAND3X0_LVT ibuf_RVCExpander_U266 ( .A1(ibuf_RVCExpander_n103), .A2(
        ibuf_RVCExpander_n61), .A3(ibuf_RVCExpander_n102), .Y(
        ibuf_RVCExpander_n104) );
  AND2X1_LVT ibuf_RVCExpander_U265 ( .A1(ibuf_RVCExpander_n37), .A2(
        ibuf_RVCExpander_n302), .Y(ibuf_RVCExpander_n103) );
  NAND2X0_LVT ibuf_RVCExpander_U264 ( .A1(ibuf_RVCExpander_n302), .A2(
        ibuf_RVCExpander_n228), .Y(ibuf_RVCExpander_n97) );
  NAND2X0_LVT ibuf_RVCExpander_U263 ( .A1(ibuf_RVCExpander_n62), .A2(
        ibuf_RVCExpander_n100), .Y(ibuf_RVCExpander_n99) );
  NAND2X0_LVT ibuf_RVCExpander_U262 ( .A1(ibuf_RVCExpander_n95), .A2(
        ibuf_RVCExpander_n108), .Y(ibuf_RVCExpander_n100) );
  AND2X1_LVT ibuf_RVCExpander_U261 ( .A1(ibuf_RVCExpander_n169), .A2(
        ibuf_RVCExpander_n94), .Y(ibuf_RVCExpander_n108) );
  NAND2X0_LVT ibuf_RVCExpander_U260 ( .A1(ibuf_RVCExpander_n93), .A2(
        ibuf_RVCExpander_n320), .Y(ibuf_RVCExpander_n288) );
  AND2X1_LVT ibuf_RVCExpander_U259 ( .A1(ibuf_RVCExpander_n92), .A2(
        ibuf_RVCExpander_n320), .Y(ibuf_RVCExpander_n291) );
  AND2X1_LVT ibuf_RVCExpander_U258 ( .A1(ibuf_RVCExpander_n91), .A2(
        ibuf_RVCExpander_n170), .Y(ibuf_RVCExpander_n169) );
  AND2X1_LVT ibuf_RVCExpander_U257 ( .A1(ibuf_n130), .A2(ibuf_RVCExpander_n89), 
        .Y(ibuf_RVCExpander_n112) );
  INVX1_LVT ibuf_RVCExpander_U256 ( .A(ibuf_RVCExpander_n213), .Y(
        ibuf_RVCExpander_n95) );
  NAND2X0_LVT ibuf_RVCExpander_U255 ( .A1(ibuf_RVCExpander_n88), .A2(
        ibuf_RVCExpander_n190), .Y(ibuf_RVCExpander_n229) );
  OR2X1_LVT ibuf_RVCExpander_U254 ( .A1(ibuf_RVCExpander_n120), .A2(
        ibuf_RVCExpander_n210), .Y(ibuf_RVCExpander_n87) );
  INVX1_LVT ibuf_RVCExpander_U253 ( .A(ibuf_io_inst_0_bits_raw[19]), .Y(
        ibuf_RVCExpander_n86) );
  AND3X1_LVT ibuf_RVCExpander_U252 ( .A1(ibuf_RVCExpander_n349), .A2(
        ibuf_RVCExpander_n84), .A3(ibuf_RVCExpander_n224), .Y(
        ibuf_RVCExpander_n85) );
  NAND2X0_LVT ibuf_RVCExpander_U251 ( .A1(ibuf_n122), .A2(
        ibuf_io_inst_0_bits_raw[18]), .Y(ibuf_RVCExpander_n224) );
  NAND2X0_LVT ibuf_RVCExpander_U250 ( .A1(ibuf_n127), .A2(ibuf_RVCExpander_n48), .Y(ibuf_RVCExpander_n84) );
  AND2X1_LVT ibuf_RVCExpander_U249 ( .A1(ibuf_RVCExpander_n201), .A2(
        ibuf_RVCExpander_n68), .Y(ibuf_RVCExpander_n225) );
  NAND4X0_LVT ibuf_RVCExpander_U248 ( .A1(ibuf_RVCExpander_n79), .A2(
        ibuf_RVCExpander_n78), .A3(ibuf_RVCExpander_n228), .A4(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n80) );
  INVX1_LVT ibuf_RVCExpander_U247 ( .A(ibuf_RVCExpander_n126), .Y(
        ibuf_RVCExpander_n228) );
  INVX1_LVT ibuf_RVCExpander_U246 ( .A(ibuf_RVCExpander_n212), .Y(
        ibuf_RVCExpander_n79) );
  OR2X1_LVT ibuf_RVCExpander_U245 ( .A1(ibuf_RVCExpander_n300), .A2(
        ibuf_RVCExpander_n205), .Y(ibuf_RVCExpander_n81) );
  NAND2X0_LVT ibuf_RVCExpander_U244 ( .A1(ibuf_n122), .A2(
        ibuf_io_inst_0_bits_raw[16]), .Y(ibuf_RVCExpander_n207) );
  AO21X1_LVT ibuf_RVCExpander_U243 ( .A1(ibuf_RVCExpander_n244), .A2(
        ibuf_RVCExpander_n211), .A3(ibuf_RVCExpander_n300), .Y(
        ibuf_RVCExpander_n82) );
  NOR3X0_LVT ibuf_RVCExpander_U242 ( .A1(ibuf_RVCExpander_n48), .A2(
        ibuf_RVCExpander_n270), .A3(ibuf_RVCExpander_n296), .Y(
        ibuf_RVCExpander_n244) );
  NAND2X0_LVT ibuf_RVCExpander_U241 ( .A1(ibuf_RVCExpander_n57), .A2(ibuf_n125), .Y(ibuf_RVCExpander_n117) );
  NAND2X0_LVT ibuf_RVCExpander_U240 ( .A1(ibuf_RVCExpander_n67), .A2(
        ibuf_RVCExpander_n242), .Y(ibuf_RVCExpander_n280) );
  NAND2X0_LVT ibuf_RVCExpander_U239 ( .A1(ibuf_RVCExpander_n241), .A2(
        ibuf_RVCExpander_n90), .Y(ibuf_RVCExpander_n256) );
  AND3X1_LVT ibuf_RVCExpander_U238 ( .A1(ibuf_RVCExpander_n50), .A2(
        ibuf_RVCExpander_n76), .A3(ibuf_RVCExpander_n77), .Y(
        ibuf_RVCExpander_n203) );
  NAND2X0_LVT ibuf_RVCExpander_U237 ( .A1(ibuf_n126), .A2(
        ibuf_RVCExpander_n172), .Y(ibuf_RVCExpander_n77) );
  AND2X1_LVT ibuf_RVCExpander_U236 ( .A1(ibuf_RVCExpander_n180), .A2(
        ibuf_RVCExpander_n211), .Y(ibuf_RVCExpander_n76) );
  NAND2X0_LVT ibuf_RVCExpander_U235 ( .A1(ibuf_RVCExpander_n126), .A2(
        ibuf_RVCExpander_n89), .Y(ibuf_RVCExpander_n180) );
  AND2X1_LVT ibuf_RVCExpander_U234 ( .A1(ibuf_RVCExpander_n320), .A2(
        ibuf_RVCExpander_n190), .Y(ibuf_RVCExpander_n126) );
  AO22X1_LVT ibuf_RVCExpander_U233 ( .A1(ibuf_RVCExpander_n320), .A2(
        ibuf_RVCExpander_n38), .A3(ibuf_n122), .A4(ibuf_io_inst_0_bits_raw[23]), .Y(ibuf_RVCExpander_n261) );
  NAND2X0_LVT ibuf_RVCExpander_U232 ( .A1(ibuf_n122), .A2(
        ibuf_io_inst_0_bits_raw[22]), .Y(ibuf_RVCExpander_n246) );
  NAND2X0_LVT ibuf_RVCExpander_U231 ( .A1(ibuf_n122), .A2(ibuf_n_T_55_84_), 
        .Y(ibuf_RVCExpander_n234) );
  AND2X1_LVT ibuf_RVCExpander_U230 ( .A1(ibuf_RVCExpander_n153), .A2(
        ibuf_RVCExpander_n154), .Y(ibuf_RVCExpander_n133) );
  OA21X1_LVT ibuf_RVCExpander_U229 ( .A1(ibuf_RVCExpander_n350), .A2(
        ibuf_RVCExpander_n71), .A3(ibuf_RVCExpander_n59), .Y(
        ibuf_RVCExpander_n181) );
  AND2X1_LVT ibuf_RVCExpander_U228 ( .A1(ibuf_RVCExpander_n96), .A2(
        ibuf_RVCExpander_n288), .Y(ibuf_RVCExpander_n94) );
  AND4X1_LVT ibuf_RVCExpander_U227 ( .A1(ibuf_RVCExpander_n317), .A2(
        ibuf_RVCExpander_n63), .A3(ibuf_RVCExpander_n242), .A4(
        ibuf_RVCExpander_n297), .Y(ibuf_RVCExpander_n243) );
  NAND3X0_LVT ibuf_RVCExpander_U226 ( .A1(ibuf_RVCExpander_n203), .A2(
        ibuf_RVCExpander_n68), .A3(ibuf_RVCExpander_n244), .Y(
        ibuf_RVCExpander_n83) );
  AND2X2_LVT ibuf_RVCExpander_U225 ( .A1(ibuf_RVCExpander_n113), .A2(ibuf_n130), .Y(ibuf_RVCExpander_n320) );
  OR2X2_LVT ibuf_RVCExpander_U224 ( .A1(ibuf_RVCExpander_n57), .A2(
        ibuf_RVCExpander_n333), .Y(ibuf_RVCExpander_n211) );
  OR2X2_LVT ibuf_RVCExpander_U223 ( .A1(ibuf_RVCExpander_n89), .A2(
        ibuf_RVCExpander_n182), .Y(ibuf_RVCExpander_n242) );
  AND2X1_LVT ibuf_RVCExpander_U222 ( .A1(ibuf_RVCExpander_n57), .A2(ibuf_n123), 
        .Y(ibuf_RVCExpander_n93) );
  OR2X2_LVT ibuf_RVCExpander_U221 ( .A1(ibuf_RVCExpander_n210), .A2(
        ibuf_RVCExpander_n209), .Y(ibuf_RVCExpander_n277) );
  OA21X2_LVT ibuf_RVCExpander_U220 ( .A1(ibuf_RVCExpander_n47), .A2(
        ibuf_RVCExpander_n178), .A3(ibuf_RVCExpander_n39), .Y(
        ibuf_io_inst_0_bits_inst_rd[4]) );
  INVX1_LVT ibuf_RVCExpander_U219 ( .A(ibuf_RVCExpander_n242), .Y(
        ibuf_RVCExpander_n174) );
  INVX1_LVT ibuf_RVCExpander_U218 ( .A(ibuf_RVCExpander_n283), .Y(
        ibuf_RVCExpander_n328) );
  NAND3X2_LVT ibuf_RVCExpander_U217 ( .A1(ibuf_RVCExpander_n226), .A2(
        ibuf_RVCExpander_n225), .A3(ibuf_RVCExpander_n85), .Y(
        ibuf_io_inst_0_bits_inst_rs1[3]) );
  INVX1_LVT ibuf_RVCExpander_U216 ( .A(ibuf_RVCExpander_n350), .Y(
        ibuf_RVCExpander_n70) );
  OR2X1_LVT ibuf_RVCExpander_U215 ( .A1(ibuf_RVCExpander_n195), .A2(
        ibuf_RVCExpander_n173), .Y(ibuf_RVCExpander_n248) );
  AND3X2_LVT ibuf_RVCExpander_U214 ( .A1(ibuf_RVCExpander_n130), .A2(
        ibuf_RVCExpander_n129), .A3(ibuf_RVCExpander_n128), .Y(n9529) );
  INVX1_LVT ibuf_RVCExpander_U213 ( .A(ibuf_RVCExpander_n296), .Y(
        ibuf_RVCExpander_n266) );
  INVX1_LVT ibuf_RVCExpander_U212 ( .A(ibuf_RVCExpander_n55), .Y(
        ibuf_RVCExpander_n301) );
  AND2X1_LVT ibuf_RVCExpander_U211 ( .A1(ibuf_RVCExpander_n315), .A2(
        ibuf_RVCExpander_n314), .Y(n9521) );
  OR2X1_LVT ibuf_RVCExpander_U210 ( .A1(ibuf_RVCExpander_n350), .A2(
        ibuf_RVCExpander_n49), .Y(ibuf_RVCExpander_n232) );
  NOR2X0_LVT ibuf_RVCExpander_U209 ( .A1(ibuf_n130), .A2(ibuf_RVCExpander_n283), .Y(ibuf_RVCExpander_n336) );
  NAND3X0_LVT ibuf_RVCExpander_U208 ( .A1(ibuf_RVCExpander_n348), .A2(
        ibuf_RVCExpander_n339), .A3(ibuf_RVCExpander_n338), .Y(n9519) );
  NAND3X0_LVT ibuf_RVCExpander_U207 ( .A1(ibuf_RVCExpander_n328), .A2(
        ibuf_RVCExpander_n228), .A3(ibuf_RVCExpander_n40), .Y(
        ibuf_RVCExpander_n206) );
  AND3X1_LVT ibuf_RVCExpander_U206 ( .A1(ibuf_RVCExpander_n286), .A2(
        ibuf_RVCExpander_n333), .A3(ibuf_RVCExpander_n59), .Y(
        ibuf_RVCExpander_n106) );
  AO22X1_LVT ibuf_RVCExpander_U205 ( .A1(ibuf_RVCExpander_n241), .A2(
        ibuf_RVCExpander_n55), .A3(ibuf_RVCExpander_n100), .A4(
        ibuf_io_inst_0_bits_raw[8]), .Y(ibuf_io_inst_0_bits_inst_rd[1]) );
  AOI22X1_LVT ibuf_RVCExpander_U204 ( .A1(ibuf_n122), .A2(
        ibuf_io_inst_0_bits_raw[30]), .A3(ibuf_RVCExpander_n340), .A4(
        ibuf_io_inst_0_bits_raw[8]), .Y(ibuf_RVCExpander_n347) );
  OR2X2_LVT ibuf_RVCExpander_U203 ( .A1(ibuf_RVCExpander_n283), .A2(
        ibuf_RVCExpander_n340), .Y(ibuf_RVCExpander_n296) );
  IBUFFX2_LVT ibuf_RVCExpander_U202 ( .A(ibuf_n125), .Y(ibuf_RVCExpander_n216)
         );
  NAND3X1_LVT ibuf_RVCExpander_U201 ( .A1(ibuf_RVCExpander_n321), .A2(
        ibuf_n125), .A3(ibuf_RVCExpander_n320), .Y(ibuf_RVCExpander_n323) );
  INVX1_LVT ibuf_RVCExpander_U200 ( .A(ibuf_io_inst_0_bits_raw[4]), .Y(
        ibuf_RVCExpander_n245) );
  NAND4X0_LVT ibuf_RVCExpander_U199 ( .A1(ibuf_RVCExpander_n348), .A2(
        ibuf_RVCExpander_n347), .A3(ibuf_RVCExpander_n346), .A4(
        ibuf_RVCExpander_n345), .Y(n9518) );
  AND2X1_LVT ibuf_RVCExpander_U198 ( .A1(ibuf_RVCExpander_n101), .A2(ibuf_n123), .Y(ibuf_RVCExpander_n88) );
  NAND4X1_LVT ibuf_RVCExpander_U197 ( .A1(ibuf_RVCExpander_n329), .A2(
        ibuf_RVCExpander_n55), .A3(ibuf_RVCExpander_n264), .A4(
        ibuf_RVCExpander_n65), .Y(ibuf_RVCExpander_n165) );
  AND2X1_LVT ibuf_RVCExpander_U196 ( .A1(ibuf_RVCExpander_n256), .A2(
        ibuf_RVCExpander_n242), .Y(ibuf_RVCExpander_n68) );
  NAND2X0_LVT ibuf_RVCExpander_U195 ( .A1(ibuf_RVCExpander_n241), .A2(
        ibuf_RVCExpander_n90), .Y(ibuf_RVCExpander_n67) );
  NAND3X0_LVT ibuf_RVCExpander_U194 ( .A1(ibuf_RVCExpander_n67), .A2(
        ibuf_RVCExpander_n38), .A3(ibuf_RVCExpander_n333), .Y(
        ibuf_RVCExpander_n255) );
  AND2X1_LVT ibuf_RVCExpander_U193 ( .A1(ibuf_RVCExpander_n75), .A2(
        ibuf_RVCExpander_n60), .Y(ibuf_RVCExpander_n101) );
  OA21X1_LVT ibuf_RVCExpander_U192 ( .A1(ibuf_RVCExpander_n216), .A2(
        ibuf_RVCExpander_n184), .A3(ibuf_RVCExpander_n183), .Y(
        ibuf_RVCExpander_n185) );
  INVX1_LVT ibuf_RVCExpander_U191 ( .A(ibuf_RVCExpander_n270), .Y(
        ibuf_RVCExpander_n201) );
  IBUFFX2_LVT ibuf_RVCExpander_U190 ( .A(ibuf_RVCExpander_n60), .Y(
        ibuf_RVCExpander_n113) );
  NAND3X0_LVT ibuf_RVCExpander_U189 ( .A1(ibuf_RVCExpander_n154), .A2(
        ibuf_RVCExpander_n153), .A3(ibuf_RVCExpander_n152), .Y(
        ibuf_RVCExpander_n158) );
  NAND2X0_LVT ibuf_RVCExpander_U188 ( .A1(ibuf_RVCExpander_n288), .A2(
        ibuf_RVCExpander_n96), .Y(ibuf_RVCExpander_n171) );
  OR2X1_LVT ibuf_RVCExpander_U187 ( .A1(ibuf_RVCExpander_n340), .A2(
        ibuf_RVCExpander_n215), .Y(ibuf_RVCExpander_n218) );
  OA21X1_LVT ibuf_RVCExpander_U186 ( .A1(ibuf_RVCExpander_n172), .A2(
        ibuf_RVCExpander_n340), .A3(ibuf_RVCExpander_n170), .Y(
        ibuf_RVCExpander_n176) );
  NAND2X0_LVT ibuf_RVCExpander_U185 ( .A1(ibuf_RVCExpander_n92), .A2(
        ibuf_RVCExpander_n101), .Y(ibuf_RVCExpander_n65) );
  NAND4X0_LVT ibuf_RVCExpander_U184 ( .A1(ibuf_RVCExpander_n200), .A2(
        ibuf_RVCExpander_n199), .A3(ibuf_RVCExpander_n198), .A4(
        ibuf_RVCExpander_n197), .Y(n9523) );
  AND3X1_LVT ibuf_RVCExpander_U183 ( .A1(ibuf_RVCExpander_n209), .A2(
        ibuf_RVCExpander_n47), .A3(ibuf_RVCExpander_n118), .Y(
        ibuf_RVCExpander_n64) );
  OA21X2_LVT ibuf_RVCExpander_U182 ( .A1(ibuf_n130), .A2(ibuf_RVCExpander_n93), 
        .A3(ibuf_RVCExpander_n60), .Y(ibuf_RVCExpander_n73) );
  NBUFFX2_LVT ibuf_RVCExpander_U181 ( .A(ibuf_n131), .Y(ibuf_RVCExpander_n60)
         );
  NAND2X0_LVT ibuf_RVCExpander_U180 ( .A1(ibuf_RVCExpander_n320), .A2(
        ibuf_RVCExpander_n89), .Y(ibuf_RVCExpander_n58) );
  OR2X1_LVT ibuf_RVCExpander_U179 ( .A1(ibuf_RVCExpander_n58), .A2(
        ibuf_RVCExpander_n90), .Y(ibuf_RVCExpander_n59) );
  NBUFFX2_LVT ibuf_RVCExpander_U178 ( .A(ibuf_n124), .Y(ibuf_RVCExpander_n57)
         );
  AND3X1_LVT ibuf_RVCExpander_U177 ( .A1(ibuf_RVCExpander_n342), .A2(
        ibuf_RVCExpander_n74), .A3(ibuf_RVCExpander_n290), .Y(
        ibuf_RVCExpander_n56) );
  NBUFFX2_LVT ibuf_RVCExpander_U176 ( .A(ibuf_n129), .Y(ibuf_RVCExpander_n55)
         );
  NAND3X0_LVT ibuf_RVCExpander_U175 ( .A1(ibuf_RVCExpander_n160), .A2(
        ibuf_RVCExpander_n349), .A3(ibuf_RVCExpander_n159), .Y(n9525) );
  NOR2X2_LVT ibuf_RVCExpander_U174 ( .A1(ibuf_RVCExpander_n283), .A2(
        ibuf_RVCExpander_n340), .Y(ibuf_RVCExpander_n349) );
  NAND3X0_LVT ibuf_RVCExpander_U173 ( .A1(ibuf_RVCExpander_n209), .A2(
        ibuf_RVCExpander_n47), .A3(ibuf_RVCExpander_n118), .Y(
        ibuf_RVCExpander_n316) );
  OR3X2_LVT ibuf_RVCExpander_U172 ( .A1(ibuf_RVCExpander_n5), .A2(
        ibuf_io_inst_0_bits_raw[11]), .A3(ibuf_RVCExpander_n116), .Y(
        ibuf_RVCExpander_n209) );
  NAND3X0_LVT ibuf_RVCExpander_U171 ( .A1(ibuf_RVCExpander_n209), .A2(
        ibuf_RVCExpander_n47), .A3(ibuf_RVCExpander_n118), .Y(
        ibuf_RVCExpander_n54) );
  NAND3X0_LVT ibuf_RVCExpander_U170 ( .A1(ibuf_RVCExpander_n209), .A2(
        ibuf_RVCExpander_n47), .A3(ibuf_RVCExpander_n118), .Y(
        ibuf_RVCExpander_n53) );
  INVX1_LVT ibuf_RVCExpander_U169 ( .A(ibuf_RVCExpander_n168), .Y(
        ibuf_RVCExpander_n66) );
  OA22X1_LVT ibuf_RVCExpander_U168 ( .A1(ibuf_RVCExpander_n290), .A2(
        ibuf_RVCExpander_n302), .A3(ibuf_RVCExpander_n289), .A4(
        ibuf_RVCExpander_n288), .Y(ibuf_RVCExpander_n294) );
  NAND2X0_LVT ibuf_RVCExpander_U167 ( .A1(ibuf_RVCExpander_n288), .A2(
        ibuf_RVCExpander_n96), .Y(ibuf_RVCExpander_n51) );
  IBUFFX2_LVT ibuf_RVCExpander_U166 ( .A(ibuf_io_inst_0_bits_raw[2]), .Y(
        ibuf_RVCExpander_n290) );
  NAND4X0_LVT ibuf_RVCExpander_U165 ( .A1(ibuf_RVCExpander_n82), .A2(
        ibuf_RVCExpander_n207), .A3(ibuf_RVCExpander_n81), .A4(
        ibuf_RVCExpander_n80), .Y(ibuf_io_inst_0_bits_inst_rs1[1]) );
  NAND2X0_LVT ibuf_RVCExpander_U164 ( .A1(ibuf_RVCExpander_n110), .A2(
        ibuf_RVCExpander_n172), .Y(ibuf_RVCExpander_n50) );
  NAND2X0_LVT ibuf_RVCExpander_U163 ( .A1(ibuf_RVCExpander_n110), .A2(
        ibuf_RVCExpander_n172), .Y(ibuf_RVCExpander_n49) );
  NOR3X0_LVT ibuf_RVCExpander_U162 ( .A1(ibuf_RVCExpander_n89), .A2(
        ibuf_RVCExpander_n216), .A3(ibuf_RVCExpander_n57), .Y(
        ibuf_RVCExpander_n92) );
  AND2X1_LVT ibuf_RVCExpander_U161 ( .A1(ibuf_RVCExpander_n92), .A2(
        ibuf_RVCExpander_n101), .Y(ibuf_RVCExpander_n340) );
  OR2X1_LVT ibuf_RVCExpander_U160 ( .A1(ibuf_n125), .A2(ibuf_RVCExpander_n333), 
        .Y(ibuf_RVCExpander_n177) );
  NAND2X0_LVT ibuf_RVCExpander_U159 ( .A1(ibuf_RVCExpander_n56), .A2(
        ibuf_RVCExpander_n172), .Y(ibuf_RVCExpander_n46) );
  AND2X4_LVT ibuf_RVCExpander_U158 ( .A1(ibuf_RVCExpander_n60), .A2(ibuf_n130), 
        .Y(ibuf_n122) );
  NAND3X0_LVT ibuf_RVCExpander_U157 ( .A1(ibuf_RVCExpander_n121), .A2(
        ibuf_RVCExpander_n216), .A3(ibuf_RVCExpander_n242), .Y(
        ibuf_RVCExpander_n122) );
  INVX1_LVT ibuf_RVCExpander_U156 ( .A(ibuf_n_T_55_85_), .Y(
        ibuf_RVCExpander_n72) );
  INVX0_LVT ibuf_RVCExpander_U155 ( .A(ibuf_n_T_55_91_), .Y(
        ibuf_RVCExpander_n303) );
  NOR2X1_LVT ibuf_RVCExpander_U154 ( .A1(ibuf_io_inst_0_bits_raw[4]), .A2(
        ibuf_RVCExpander_n55), .Y(ibuf_RVCExpander_n74) );
  INVX0_LVT ibuf_RVCExpander_U153 ( .A(ibuf_RVCExpander_n63), .Y(
        ibuf_RVCExpander_n298) );
  INVX0_LVT ibuf_RVCExpander_U152 ( .A(ibuf_RVCExpander_n342), .Y(
        ibuf_RVCExpander_n196) );
  NAND3X0_LVT ibuf_RVCExpander_U151 ( .A1(ibuf_io_inst_0_bits_raw[8]), .A2(
        ibuf_RVCExpander_n216), .A3(ibuf_n123), .Y(ibuf_RVCExpander_n217) );
  INVX1_LVT ibuf_RVCExpander_U150 ( .A(ibuf_RVCExpander_n241), .Y(
        ibuf_RVCExpander_n182) );
  OAI21X1_LVT ibuf_RVCExpander_U149 ( .A1(ibuf_RVCExpander_n245), .A2(
        ibuf_RVCExpander_n73), .A3(ibuf_RVCExpander_n246), .Y(
        ibuf_io_inst_0_bits_inst_rs2[2]) );
  OR2X1_LVT ibuf_RVCExpander_U148 ( .A1(ibuf_RVCExpander_n72), .A2(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n237) );
  OR2X1_LVT ibuf_RVCExpander_U147 ( .A1(ibuf_RVCExpander_n1), .A2(
        ibuf_RVCExpander_n40), .Y(ibuf_RVCExpander_n129) );
  NOR2X1_LVT ibuf_RVCExpander_U146 ( .A1(ibuf_RVCExpander_n89), .A2(
        ibuf_RVCExpander_n71), .Y(ibuf_RVCExpander_n204) );
  NOR2X1_LVT ibuf_RVCExpander_U145 ( .A1(ibuf_RVCExpander_n5), .A2(
        ibuf_RVCExpander_n39), .Y(ibuf_RVCExpander_n109) );
  OAI21X1_LVT ibuf_RVCExpander_U144 ( .A1(ibuf_RVCExpander_n301), .A2(
        ibuf_RVCExpander_n73), .A3(ibuf_RVCExpander_n237), .Y(
        ibuf_io_inst_0_bits_inst_rs2[1]) );
  OR2X1_LVT ibuf_RVCExpander_U143 ( .A1(ibuf_RVCExpander_n350), .A2(
        ibuf_RVCExpander_n53), .Y(ibuf_RVCExpander_n275) );
  AND2X1_LVT ibuf_RVCExpander_U142 ( .A1(ibuf_RVCExpander_n211), .A2(
        ibuf_RVCExpander_n177), .Y(ibuf_RVCExpander_n317) );
  OR2X1_LVT ibuf_RVCExpander_U141 ( .A1(ibuf_RVCExpander_n61), .A2(
        ibuf_RVCExpander_n110), .Y(ibuf_RVCExpander_n170) );
  AND2X1_LVT ibuf_RVCExpander_U140 ( .A1(ibuf_RVCExpander_n190), .A2(
        ibuf_RVCExpander_n34), .Y(ibuf_RVCExpander_n270) );
  NOR2X1_LVT ibuf_RVCExpander_U139 ( .A1(ibuf_n122), .A2(ibuf_RVCExpander_n291), .Y(ibuf_RVCExpander_n96) );
  INVX1_LVT ibuf_RVCExpander_U138 ( .A(ibuf_RVCExpander_n277), .Y(
        ibuf_RVCExpander_n325) );
  INVX0_LVT ibuf_RVCExpander_U137 ( .A(ibuf_RVCExpander_n317), .Y(
        ibuf_RVCExpander_n257) );
  OR2X1_LVT ibuf_RVCExpander_U136 ( .A1(ibuf_RVCExpander_n261), .A2(
        ibuf_RVCExpander_n336), .Y(ibuf_io_inst_0_bits_inst_rs2[3]) );
  NOR2X1_LVT ibuf_RVCExpander_U135 ( .A1(ibuf_RVCExpander_n174), .A2(
        ibuf_RVCExpander_n279), .Y(ibuf_RVCExpander_n264) );
  INVX0_LVT ibuf_RVCExpander_U134 ( .A(ibuf_RVCExpander_n279), .Y(
        ibuf_RVCExpander_n161) );
  NOR2X1_LVT ibuf_RVCExpander_U133 ( .A1(ibuf_RVCExpander_n280), .A2(
        ibuf_RVCExpander_n279), .Y(ibuf_RVCExpander_n337) );
  INVX0_LVT ibuf_RVCExpander_U132 ( .A(ibuf_RVCExpander_n104), .Y(
        ibuf_RVCExpander_n107) );
  NAND3X1_LVT ibuf_RVCExpander_U131 ( .A1(ibuf_RVCExpander_n194), .A2(
        ibuf_RVCExpander_n193), .A3(ibuf_RVCExpander_n192), .Y(n9524) );
  AO22X1_LVT ibuf_RVCExpander_U130 ( .A1(ibuf_RVCExpander_n107), .A2(
        ibuf_RVCExpander_n106), .A3(ibuf_n127), .A4(ibuf_RVCExpander_n105), 
        .Y(ibuf_io_inst_0_bits_inst_rd[3]) );
  NAND3X0_LVT ibuf_RVCExpander_U129 ( .A1(ibuf_RVCExpander_n99), .A2(
        ibuf_RVCExpander_n232), .A3(ibuf_RVCExpander_n98), .Y(
        ibuf_io_inst_0_bits_inst_rd[0]) );
  INVX1_LVT ibuf_RVCExpander_U128 ( .A(ibuf_n126), .Y(ibuf_RVCExpander_n350)
         );
  INVX0_LVT ibuf_RVCExpander_U127 ( .A(ibuf_n127), .Y(ibuf_RVCExpander_n344)
         );
  IBUFFX2_LVT ibuf_RVCExpander_U126 ( .A(ibuf_n122), .Y(ibuf_RVCExpander_n40)
         );
  INVX0_LVT ibuf_RVCExpander_U125 ( .A(ibuf_n130), .Y(ibuf_RVCExpander_n75) );
  NOR2X1_LVT ibuf_RVCExpander_U124 ( .A1(ibuf_RVCExpander_n117), .A2(
        ibuf_RVCExpander_n333), .Y(ibuf_RVCExpander_n48) );
  OR2X1_LVT ibuf_RVCExpander_U123 ( .A1(ibuf_RVCExpander_n117), .A2(
        ibuf_RVCExpander_n333), .Y(ibuf_RVCExpander_n210) );
  INVX1_LVT ibuf_RVCExpander_U122 ( .A(ibuf_RVCExpander_n211), .Y(
        ibuf_RVCExpander_n115) );
  NAND2X1_LVT ibuf_RVCExpander_U121 ( .A1(ibuf_RVCExpander_n227), .A2(
        ibuf_RVCExpander_n87), .Y(ibuf_io_inst_0_bits_inst_rs1[4]) );
  OR2X2_LVT ibuf_RVCExpander_U120 ( .A1(ibuf_RVCExpander_n97), .A2(
        ibuf_RVCExpander_n51), .Y(ibuf_RVCExpander_n162) );
  AND3X2_LVT ibuf_RVCExpander_U119 ( .A1(ibuf_RVCExpander_n75), .A2(
        ibuf_RVCExpander_n60), .A3(ibuf_RVCExpander_n89), .Y(
        ibuf_RVCExpander_n47) );
  NAND3X2_LVT ibuf_RVCExpander_U118 ( .A1(ibuf_RVCExpander_n75), .A2(
        ibuf_RVCExpander_n60), .A3(ibuf_RVCExpander_n89), .Y(
        ibuf_RVCExpander_n333) );
  NOR2X4_LVT ibuf_RVCExpander_U117 ( .A1(ibuf_n130), .A2(ibuf_RVCExpander_n60), 
        .Y(ibuf_RVCExpander_n241) );
  NAND3X2_LVT ibuf_RVCExpander_U116 ( .A1(ibuf_RVCExpander_n112), .A2(
        ibuf_RVCExpander_n113), .A3(ibuf_RVCExpander_n90), .Y(
        ibuf_RVCExpander_n302) );
  AND3X4_LVT ibuf_RVCExpander_U115 ( .A1(ibuf_RVCExpander_n320), .A2(ibuf_n123), .A3(ibuf_RVCExpander_n190), .Y(ibuf_RVCExpander_n172) );
  NAND3X1_LVT ibuf_RVCExpander_U114 ( .A1(ibuf_RVCExpander_n320), .A2(
        ibuf_n123), .A3(ibuf_RVCExpander_n190), .Y(ibuf_RVCExpander_n61) );
  NAND3X2_LVT ibuf_RVCExpander_U113 ( .A1(ibuf_RVCExpander_n270), .A2(
        ibuf_RVCExpander_n9), .A3(ibuf_RVCExpander_n38), .Y(
        ibuf_RVCExpander_n183) );
  IBUFFX2_LVT ibuf_RVCExpander_U112 ( .A(ibuf_RVCExpander_n2), .Y(
        ibuf_RVCExpander_n151) );
  IBUFFX2_LVT ibuf_RVCExpander_U111 ( .A(ibuf_RVCExpander_n163), .Y(
        ibuf_RVCExpander_n233) );
  NAND3X2_LVT ibuf_RVCExpander_U110 ( .A1(ibuf_RVCExpander_n90), .A2(
        ibuf_RVCExpander_n320), .A3(ibuf_RVCExpander_n70), .Y(
        ibuf_RVCExpander_n268) );
  IBUFFX2_LVT ibuf_RVCExpander_U109 ( .A(ibuf_io_inst_0_bits_raw[11]), .Y(
        ibuf_RVCExpander_n120) );
  NAND2X0_LVT ibuf_RVCExpander_U108 ( .A1(ibuf_RVCExpander_n92), .A2(
        ibuf_RVCExpander_n320), .Y(ibuf_RVCExpander_n37) );
  NAND2X0_LVT ibuf_RVCExpander_U107 ( .A1(ibuf_RVCExpander_n332), .A2(
        ibuf_RVCExpander_n331), .Y(n9520) );
  OR2X2_LVT ibuf_RVCExpander_U106 ( .A1(ibuf_RVCExpander_n188), .A2(
        ibuf_RVCExpander_n229), .Y(ibuf_RVCExpander_n334) );
  AND3X4_LVT ibuf_RVCExpander_U105 ( .A1(ibuf_RVCExpander_n229), .A2(
        ibuf_RVCExpander_n228), .A3(ibuf_RVCExpander_n242), .Y(
        ibuf_RVCExpander_n250) );
  OR3X2_LVT ibuf_RVCExpander_U104 ( .A1(ibuf_RVCExpander_n101), .A2(
        ibuf_RVCExpander_n290), .A3(ibuf_RVCExpander_n162), .Y(
        ibuf_RVCExpander_n98) );
  NAND3X2_LVT ibuf_RVCExpander_U103 ( .A1(ibuf_RVCExpander_n101), .A2(
        ibuf_n123), .A3(ibuf_n125), .Y(ibuf_RVCExpander_n102) );
  AO22X2_LVT ibuf_RVCExpander_U102 ( .A1(ibuf_RVCExpander_n241), .A2(
        ibuf_RVCExpander_n52), .A3(ibuf_RVCExpander_n100), .A4(
        ibuf_RVCExpander_n66), .Y(ibuf_io_inst_0_bits_inst_rd[2]) );
  AND2X4_LVT ibuf_RVCExpander_U101 ( .A1(ibuf_RVCExpander_n168), .A2(
        ibuf_RVCExpander_n120), .Y(ibuf_RVCExpander_n153) );
  AND4X2_LVT ibuf_RVCExpander_U100 ( .A1(ibuf_RVCExpander_n115), .A2(
        ibuf_RVCExpander_n114), .A3(ibuf_RVCExpander_n300), .A4(
        ibuf_RVCExpander_n289), .Y(ibuf_RVCExpander_n36) );
  AOI21X1_LVT ibuf_RVCExpander_U99 ( .A1(ibuf_RVCExpander_n35), .A2(
        ibuf_RVCExpander_n163), .A3(ibuf_RVCExpander_n36), .Y(
        ibuf_RVCExpander_n119) );
  OR2X2_LVT ibuf_RVCExpander_U98 ( .A1(ibuf_RVCExpander_n172), .A2(
        ibuf_RVCExpander_n171), .Y(ibuf_RVCExpander_n309) );
  IBUFFX2_LVT ibuf_RVCExpander_U97 ( .A(ibuf_RVCExpander_n120), .Y(
        ibuf_RVCExpander_n39) );
  AND4X2_LVT ibuf_RVCExpander_U96 ( .A1(ibuf_n125), .A2(ibuf_RVCExpander_n120), 
        .A3(ibuf_RVCExpander_n168), .A4(ibuf_RVCExpander_n344), .Y(
        ibuf_RVCExpander_n114) );
  OA21X2_LVT ibuf_RVCExpander_U95 ( .A1(ibuf_RVCExpander_n53), .A2(
        ibuf_RVCExpander_n301), .A3(ibuf_RVCExpander_n334), .Y(
        ibuf_RVCExpander_n194) );
  AND2X4_LVT ibuf_RVCExpander_U94 ( .A1(ibuf_RVCExpander_n334), .A2(
        ibuf_RVCExpander_n317), .Y(ibuf_RVCExpander_n276) );
  NAND3X2_LVT ibuf_RVCExpander_U93 ( .A1(ibuf_RVCExpander_n318), .A2(
        ibuf_RVCExpander_n317), .A3(ibuf_RVCExpander_n334), .Y(
        ibuf_RVCExpander_n319) );
  AND2X1_LVT ibuf_RVCExpander_U92 ( .A1(ibuf_RVCExpander_n101), .A2(ibuf_n123), 
        .Y(ibuf_RVCExpander_n34) );
  NAND3X1_LVT ibuf_RVCExpander_U91 ( .A1(ibuf_RVCExpander_n277), .A2(
        ibuf_RVCExpander_n317), .A3(ibuf_RVCExpander_n343), .Y(
        ibuf_RVCExpander_n265) );
  OR2X4_LVT ibuf_RVCExpander_U90 ( .A1(ibuf_RVCExpander_n343), .A2(
        ibuf_RVCExpander_n344), .Y(ibuf_RVCExpander_n345) );
  NAND2X2_LVT ibuf_RVCExpander_U89 ( .A1(ibuf_RVCExpander_n274), .A2(
        ibuf_RVCExpander_n273), .Y(n9522) );
  OR3X2_LVT ibuf_RVCExpander_U88 ( .A1(ibuf_RVCExpander_n146), .A2(
        ibuf_RVCExpander_n171), .A3(ibuf_RVCExpander_n145), .Y(
        ibuf_RVCExpander_n150) );
  INVX1_LVT ibuf_RVCExpander_U87 ( .A(ibuf_RVCExpander_n151), .Y(
        ibuf_RVCExpander_n38) );
  INVX0_LVT ibuf_RVCExpander_U85 ( .A(ibuf_RVCExpander_n235), .Y(
        ibuf_RVCExpander_n32) );
  OA221X1_LVT ibuf_RVCExpander_U83 ( .A1(ibuf_RVCExpander_n263), .A2(
        ibuf_RVCExpander_n264), .A3(ibuf_RVCExpander_n263), .A4(
        ibuf_RVCExpander_n39), .A5(ibuf_RVCExpander_n336), .Y(
        ibuf_RVCExpander_n30) );
  AND2X4_LVT ibuf_RVCExpander_U82 ( .A1(ibuf_RVCExpander_n300), .A2(
        ibuf_RVCExpander_n29), .Y(ibuf_RVCExpander_n212) );
  NAND2X0_LVT ibuf_RVCExpander_U81 ( .A1(ibuf_RVCExpander_n67), .A2(
        ibuf_RVCExpander_n242), .Y(ibuf_RVCExpander_n29) );
  NAND2X0_LVT ibuf_RVCExpander_U80 ( .A1(ibuf_RVCExpander_n226), .A2(
        ibuf_RVCExpander_n28), .Y(io_fpu_inst[18]) );
  AND4X1_LVT ibuf_RVCExpander_U79 ( .A1(ibuf_RVCExpander_n224), .A2(
        ibuf_RVCExpander_n328), .A3(ibuf_RVCExpander_n225), .A4(
        ibuf_RVCExpander_n235), .Y(ibuf_RVCExpander_n28) );
  NAND3X0_LVT ibuf_RVCExpander_U78 ( .A1(ibuf_RVCExpander_n222), .A2(
        ibuf_RVCExpander_n26), .A3(ibuf_RVCExpander_n27), .Y(io_fpu_inst[15])
         );
  INVX0_LVT ibuf_RVCExpander_U77 ( .A(ibuf_RVCExpander_n204), .Y(
        ibuf_RVCExpander_n27) );
  AOI22X1_LVT ibuf_RVCExpander_U76 ( .A1(ibuf_RVCExpander_n62), .A2(
        ibuf_RVCExpander_n221), .A3(ibuf_RVCExpander_n64), .A4(
        ibuf_RVCExpander_n38), .Y(ibuf_RVCExpander_n26) );
  OA21X1_LVT ibuf_RVCExpander_U75 ( .A1(ibuf_RVCExpander_n178), .A2(
        ibuf_RVCExpander_n25), .A3(ibuf_RVCExpander_n39), .Y(io_fpu_inst[11])
         );
  NAND4X0_LVT ibuf_RVCExpander_U74 ( .A1(ibuf_RVCExpander_n242), .A2(
        ibuf_RVCExpander_n210), .A3(ibuf_RVCExpander_n317), .A4(
        ibuf_RVCExpander_n328), .Y(ibuf_RVCExpander_n25) );
  NAND3X0_LVT ibuf_RVCExpander_U73 ( .A1(ibuf_RVCExpander_n24), .A2(
        ibuf_RVCExpander_n23), .A3(ibuf_RVCExpander_n22), .Y(io_fpu_inst[9])
         );
  OR2X1_LVT ibuf_RVCExpander_U72 ( .A1(ibuf_RVCExpander_n168), .A2(
        ibuf_RVCExpander_n17), .Y(ibuf_RVCExpander_n24) );
  NAND2X0_LVT ibuf_RVCExpander_U71 ( .A1(ibuf_RVCExpander_n283), .A2(
        ibuf_RVCExpander_n52), .Y(ibuf_RVCExpander_n23) );
  NAND2X0_LVT ibuf_RVCExpander_U70 ( .A1(ibuf_RVCExpander_n10), .A2(
        ibuf_RVCExpander_n21), .Y(ibuf_RVCExpander_n22) );
  NAND3X0_LVT ibuf_RVCExpander_U69 ( .A1(ibuf_RVCExpander_n20), .A2(
        ibuf_RVCExpander_n19), .A3(ibuf_RVCExpander_n18), .Y(
        ibuf_RVCExpander_n21) );
  NAND2X0_LVT ibuf_RVCExpander_U68 ( .A1(ibuf_RVCExpander_n66), .A2(
        ibuf_RVCExpander_n279), .Y(ibuf_RVCExpander_n20) );
  NAND3X0_LVT ibuf_RVCExpander_U67 ( .A1(ibuf_RVCExpander_n174), .A2(
        ibuf_RVCExpander_n216), .A3(ibuf_RVCExpander_n63), .Y(
        ibuf_RVCExpander_n19) );
  NAND3X0_LVT ibuf_RVCExpander_U66 ( .A1(ibuf_RVCExpander_n349), .A2(
        ibuf_RVCExpander_n52), .A3(ibuf_RVCExpander_n264), .Y(
        ibuf_RVCExpander_n18) );
  OAI222X1_LVT ibuf_RVCExpander_U64 ( .A1(ibuf_RVCExpander_n11), .A2(
        ibuf_RVCExpander_n12), .A3(ibuf_RVCExpander_n163), .A4(
        ibuf_RVCExpander_n232), .A5(ibuf_RVCExpander_n162), .A6(
        ibuf_RVCExpander_n15), .Y(io_fpu_inst[7]) );
  NAND3X0_LVT ibuf_RVCExpander_U62 ( .A1(ibuf_RVCExpander_n266), .A2(
        ibuf_RVCExpander_n1), .A3(ibuf_RVCExpander_n264), .Y(
        ibuf_RVCExpander_n13) );
  INVX0_LVT ibuf_RVCExpander_U61 ( .A(ibuf_RVCExpander_n164), .Y(
        ibuf_RVCExpander_n12) );
  INVX0_LVT ibuf_RVCExpander_U60 ( .A(ibuf_RVCExpander_n62), .Y(
        ibuf_RVCExpander_n11) );
  INVX1_LVT ibuf_RVCExpander_U59 ( .A(ibuf_n123), .Y(ibuf_RVCExpander_n89) );
  IBUFFX2_LVT ibuf_RVCExpander_U58 ( .A(ibuf_io_inst_0_bits_raw[8]), .Y(
        ibuf_RVCExpander_n300) );
  INVX1_LVT ibuf_RVCExpander_U57 ( .A(ibuf_RVCExpander_n289), .Y(
        ibuf_RVCExpander_n62) );
  NAND3X0_LVT ibuf_RVCExpander_U56 ( .A1(ibuf_RVCExpander_n185), .A2(
        ibuf_RVCExpander_n186), .A3(ibuf_RVCExpander_n200), .Y(io_fpu_inst[12]) );
  INVX1_LVT ibuf_RVCExpander_U55 ( .A(ibuf_RVCExpander_n162), .Y(
        ibuf_RVCExpander_n329) );
  OA21X1_LVT ibuf_RVCExpander_U54 ( .A1(ibuf_RVCExpander_n270), .A2(
        ibuf_RVCExpander_n325), .A3(ibuf_RVCExpander_n343), .Y(
        ibuf_RVCExpander_n271) );
  INVX1_LVT ibuf_RVCExpander_U53 ( .A(ibuf_RVCExpander_n248), .Y(
        ibuf_RVCExpander_n35) );
  NAND4X0_LVT ibuf_RVCExpander_U52 ( .A1(ibuf_RVCExpander_n155), .A2(
        ibuf_RVCExpander_n157), .A3(ibuf_RVCExpander_n156), .A4(
        ibuf_RVCExpander_n260), .Y(n9526) );
  INVX1_LVT ibuf_RVCExpander_U51 ( .A(ibuf_RVCExpander_n245), .Y(
        ibuf_RVCExpander_n52) );
  INVX1_LVT ibuf_RVCExpander_U50 ( .A(ibuf_n122), .Y(ibuf_RVCExpander_n71) );
  AO21X1_LVT ibuf_RVCExpander_U49 ( .A1(ibuf_RVCExpander_n70), .A2(
        ibuf_RVCExpander_n163), .A3(ibuf_RVCExpander_n49), .Y(
        ibuf_RVCExpander_n127) );
  IBUFFX2_LVT ibuf_RVCExpander_U48 ( .A(ibuf_RVCExpander_n101), .Y(
        ibuf_RVCExpander_n78) );
  OR2X2_LVT ibuf_RVCExpander_U47 ( .A1(ibuf_n125), .A2(ibuf_RVCExpander_n57), 
        .Y(ibuf_RVCExpander_n90) );
  NOR2X2_LVT ibuf_RVCExpander_U46 ( .A1(ibuf_n125), .A2(ibuf_RVCExpander_n57), 
        .Y(ibuf_RVCExpander_n190) );
  NAND3X2_LVT ibuf_RVCExpander_U45 ( .A1(ibuf_RVCExpander_n330), .A2(
        ibuf_RVCExpander_n329), .A3(ibuf_RVCExpander_n328), .Y(
        ibuf_RVCExpander_n331) );
  NAND3X0_LVT ibuf_RVCExpander_U44 ( .A1(ibuf_RVCExpander_n144), .A2(
        ibuf_RVCExpander_n143), .A3(ibuf_RVCExpander_n142), .Y(n9528) );
  NAND3X2_LVT ibuf_RVCExpander_U43 ( .A1(ibuf_RVCExpander_n10), .A2(
        ibuf_RVCExpander_n244), .A3(ibuf_RVCExpander_n243), .Y(
        ibuf_RVCExpander_n254) );
  NAND3X0_LVT ibuf_RVCExpander_U42 ( .A1(ibuf_RVCExpander_n140), .A2(
        ibuf_RVCExpander_n329), .A3(ibuf_RVCExpander_n328), .Y(
        ibuf_RVCExpander_n144) );
  AND2X4_LVT ibuf_RVCExpander_U41 ( .A1(ibuf_RVCExpander_n101), .A2(
        ibuf_RVCExpander_n93), .Y(ibuf_RVCExpander_n283) );
  NAND2X0_LVT ibuf_RVCExpander_U40 ( .A1(ibuf_RVCExpander_n353), .A2(
        ibuf_RVCExpander_n352), .Y(n9517) );
  AO21X2_LVT ibuf_RVCExpander_U39 ( .A1(ibuf_RVCExpander_n283), .A2(
        ibuf_RVCExpander_n216), .A3(ibuf_RVCExpander_n279), .Y(
        ibuf_RVCExpander_n213) );
  IBUFFX2_LVT ibuf_RVCExpander_U38 ( .A(ibuf_RVCExpander_n320), .Y(
        ibuf_RVCExpander_n285) );
  DELLN2X2_LVT ibuf_RVCExpander_U37 ( .A(ibuf_n128), .Y(ibuf_RVCExpander_n63)
         );
  IBUFFX2_LVT ibuf_RVCExpander_U36 ( .A(ibuf_RVCExpander_n162), .Y(
        ibuf_RVCExpander_n10) );
  AND2X4_LVT ibuf_RVCExpander_U35 ( .A1(ibuf_RVCExpander_n180), .A2(
        ibuf_RVCExpander_n302), .Y(ibuf_RVCExpander_n91) );
  OA22X2_LVT ibuf_RVCExpander_U34 ( .A1(ibuf_RVCExpander_n71), .A2(
        ibuf_RVCExpander_n86), .A3(ibuf_RVCExpander_n120), .A4(
        ibuf_RVCExpander_n203), .Y(ibuf_RVCExpander_n227) );
  NAND3X2_LVT ibuf_RVCExpander_U33 ( .A1(ibuf_RVCExpander_n203), .A2(
        ibuf_RVCExpander_n68), .A3(ibuf_RVCExpander_n202), .Y(
        ibuf_RVCExpander_n221) );
  AND3X2_LVT ibuf_RVCExpander_U32 ( .A1(ibuf_RVCExpander_n342), .A2(
        ibuf_RVCExpander_n300), .A3(ibuf_RVCExpander_n350), .Y(
        ibuf_RVCExpander_n132) );
  NAND3X2_LVT ibuf_RVCExpander_U31 ( .A1(ibuf_RVCExpander_n56), .A2(
        ibuf_RVCExpander_n48), .A3(ibuf_RVCExpander_n350), .Y(
        ibuf_RVCExpander_n111) );
  NBUFFX2_LVT ibuf_RVCExpander_U30 ( .A(ibuf_n128), .Y(ibuf_RVCExpander_n9) );
  AND2X4_LVT ibuf_RVCExpander_U29 ( .A1(ibuf_n122), .A2(
        ibuf_io_inst_0_bits_raw[17]), .Y(ibuf_RVCExpander_n223) );
  NAND3X2_LVT ibuf_RVCExpander_U28 ( .A1(ibuf_RVCExpander_n154), .A2(
        ibuf_RVCExpander_n153), .A3(ibuf_RVCExpander_n152), .Y(
        ibuf_RVCExpander_n8) );
  OR2X4_LVT ibuf_RVCExpander_U27 ( .A1(ibuf_RVCExpander_n179), .A2(
        ibuf_RVCExpander_n6), .Y(ibuf_RVCExpander_n343) );
  NAND2X0_LVT ibuf_RVCExpander_U26 ( .A1(ibuf_RVCExpander_n7), .A2(
        ibuf_RVCExpander_n333), .Y(ibuf_RVCExpander_n279) );
  NAND2X0_LVT ibuf_RVCExpander_U25 ( .A1(ibuf_RVCExpander_n88), .A2(
        ibuf_RVCExpander_n190), .Y(ibuf_RVCExpander_n7) );
  NAND2X0_LVT ibuf_RVCExpander_U24 ( .A1(ibuf_RVCExpander_n88), .A2(
        ibuf_RVCExpander_n190), .Y(ibuf_RVCExpander_n6) );
  AO21X2_LVT ibuf_RVCExpander_U23 ( .A1(ibuf_RVCExpander_n83), .A2(
        ibuf_RVCExpander_n62), .A3(ibuf_RVCExpander_n204), .Y(
        ibuf_io_inst_0_bits_inst_rs1[0]) );
  OR2X4_LVT ibuf_RVCExpander_U22 ( .A1(ibuf_n127), .A2(
        ibuf_io_inst_0_bits_raw[7]), .Y(ibuf_RVCExpander_n116) );
  NBUFFX2_LVT ibuf_RVCExpander_U21 ( .A(ibuf_io_inst_0_bits_raw[9]), .Y(
        ibuf_RVCExpander_n5) );
  AO22X1_LVT ibuf_RVCExpander_U20 ( .A1(ibuf_RVCExpander_n320), .A2(
        ibuf_RVCExpander_n9), .A3(ibuf_n122), .A4(ibuf_io_inst_0_bits_raw[24]), 
        .Y(ibuf_RVCExpander_n354) );
  AO22X2_LVT ibuf_RVCExpander_U19 ( .A1(ibuf_RVCExpander_n320), .A2(
        ibuf_RVCExpander_n9), .A3(ibuf_n122), .A4(ibuf_io_inst_0_bits_raw[24]), 
        .Y(ibuf_io_inst_0_bits_inst_rs2[4]) );
  AND3X2_LVT ibuf_RVCExpander_U18 ( .A1(ibuf_RVCExpander_n154), .A2(
        ibuf_RVCExpander_n109), .A3(ibuf_RVCExpander_n300), .Y(
        ibuf_RVCExpander_n163) );
  AND2X1_LVT ibuf_RVCExpander_U17 ( .A1(ibuf_RVCExpander_n56), .A2(
        ibuf_RVCExpander_n172), .Y(ibuf_RVCExpander_n3) );
  NBUFFX2_LVT ibuf_RVCExpander_U16 ( .A(ibuf_io_inst_0_bits_raw[5]), .Y(
        ibuf_RVCExpander_n2) );
  NBUFFX2_LVT ibuf_RVCExpander_U15 ( .A(ibuf_io_inst_0_bits_raw[2]), .Y(
        ibuf_RVCExpander_n1) );
  NAND3X0_LVT ibuf_RVCExpander_U14 ( .A1(ibuf_RVCExpander_n133), .A2(
        ibuf_RVCExpander_n342), .A3(ibuf_RVCExpander_n152), .Y(
        ibuf_RVCExpander_n121) );
  OAI21X2_LVT ibuf_RVCExpander_U13 ( .A1(ibuf_RVCExpander_n290), .A2(
        ibuf_RVCExpander_n73), .A3(ibuf_RVCExpander_n234), .Y(
        ibuf_io_inst_0_bits_inst_rs2[0]) );
  AND3X1_LVT ibuf_RVCExpander_U12 ( .A1(ibuf_RVCExpander_n46), .A2(
        ibuf_RVCExpander_n77), .A3(ibuf_RVCExpander_n180), .Y(
        ibuf_RVCExpander_n205) );
  OA21X1_LVT ibuf_RVCExpander_U11 ( .A1(ibuf_RVCExpander_n70), .A2(
        ibuf_RVCExpander_n46), .A3(ibuf_RVCExpander_n248), .Y(
        ibuf_RVCExpander_n141) );
  AO21X1_LVT ibuf_RVCExpander_U10 ( .A1(ibuf_RVCExpander_n66), .A2(
        ibuf_RVCExpander_n83), .A3(ibuf_RVCExpander_n223), .Y(
        ibuf_io_inst_0_bits_inst_rs1[2]) );
  AND3X1_LVT ibuf_RVCExpander_U9 ( .A1(ibuf_RVCExpander_n342), .A2(
        ibuf_RVCExpander_n74), .A3(ibuf_RVCExpander_n290), .Y(
        ibuf_RVCExpander_n110) );
  OR2X1_LVT ibuf_RVCExpander_U8 ( .A1(ibuf_RVCExpander_n344), .A2(
        ibuf_RVCExpander_n203), .Y(ibuf_RVCExpander_n226) );
  NOR2X2_LVT ibuf_RVCExpander_U7 ( .A1(ibuf_n128), .A2(ibuf_RVCExpander_n2), 
        .Y(ibuf_RVCExpander_n342) );
  OA221X1_LVT ibuf_RVCExpander_U6 ( .A1(1'b0), .A2(ibuf_RVCExpander_n335), 
        .A3(ibuf_RVCExpander_n289), .A4(ibuf_RVCExpander_n161), .A5(
        ibuf_RVCExpander_n13), .Y(ibuf_RVCExpander_n15) );
  OA221X1_LVT ibuf_RVCExpander_U5 ( .A1(1'b0), .A2(ibuf_RVCExpander_n40), .A3(
        ibuf_n125), .A4(ibuf_RVCExpander_n288), .A5(ibuf_RVCExpander_n169), 
        .Y(ibuf_RVCExpander_n17) );
  AO221X1_LVT ibuf_RVCExpander_U4 ( .A1(1'b1), .A2(ibuf_RVCExpander_n30), .A3(
        ibuf_RVCExpander_n63), .A4(ibuf_RVCExpander_n265), .A5(
        ibuf_RVCExpander_n354), .Y(io_fpu_inst[24]) );
  AO221X1_LVT ibuf_RVCExpander_U3 ( .A1(1'b1), .A2(ibuf_RVCExpander_n223), 
        .A3(ibuf_RVCExpander_n66), .A4(ibuf_RVCExpander_n221), .A5(
        ibuf_RVCExpander_n32), .Y(io_fpu_inst[17]) );
  NAND2X0_LVT csr_U2908 ( .A1(csr_n589), .A2(csr_n1907), .Y(csr_n1908) );
  NAND2X0_LVT csr_U2907 ( .A1(csr_n1474), .A2(csr_n1905), .Y(csr_n1906) );
  NAND2X0_LVT csr_U2906 ( .A1(csr_n589), .A2(csr_n1904), .Y(csr_n1905) );
  AND2X1_LVT csr_U2905 ( .A1(io_imem_sfence_bits_addr[1]), .A2(csr_n516), .Y(
        csr_n1900) );
  OA21X1_LVT csr_U2904 ( .A1(csr_n1474), .A2(csr_n1475), .A3(
        csr_read_mideleg_1), .Y(csr_n1901) );
  AO221X1_LVT csr_U2903 ( .A1(csr_n1899), .A2(csr_n407), .A3(csr_n1899), .A4(
        csr_n1898), .A5(csr_n1476), .Y(csr_n1902) );
  AND3X1_LVT csr_U2902 ( .A1(csr_io_rw_addr[1]), .A2(csr_n504), .A3(csr_n1486), 
        .Y(csr_n2166) );
  AND2X1_LVT csr_U2901 ( .A1(csr_n1487), .A2(csr_n504), .Y(csr_n2167) );
  AND2X1_LVT csr_U2900 ( .A1(csr_n504), .A2(csr_n1465), .Y(csr_n2168) );
  AND2X1_LVT csr_U2899 ( .A1(csr_n504), .A2(csr_n1484), .Y(csr_n2169) );
  AO22X1_LVT csr_U2898 ( .A1(csr_n515), .A2(csr_wdata_1_), .A3(csr_n450), .A4(
        csr_io_pc[1]), .Y(csr_net35301) );
  AO22X1_LVT csr_U2897 ( .A1(csr_n514), .A2(csr_wdata_1_), .A3(csr_n449), .A4(
        csr_io_pc[1]), .Y(csr_net35079) );
  AO22X1_LVT csr_U2896 ( .A1(csr_n513), .A2(csr_wdata_1_), .A3(csr_n448), .A4(
        csr_io_pc[1]), .Y(csr_net34877) );
  AND2X1_LVT csr_U2895 ( .A1(csr_n1897), .A2(io_ptw_pmp_7_addr[6]), .Y(
        io_ptw_pmp_7_mask[9]) );
  AND2X1_LVT csr_U2894 ( .A1(csr_n1896), .A2(io_ptw_pmp_7_addr[5]), .Y(
        io_ptw_pmp_7_mask[8]) );
  AND2X1_LVT csr_U2893 ( .A1(csr_n1895), .A2(io_ptw_pmp_7_addr[4]), .Y(
        io_ptw_pmp_7_mask[7]) );
  AND2X1_LVT csr_U2892 ( .A1(csr_n1894), .A2(io_ptw_pmp_7_addr[2]), .Y(
        io_ptw_pmp_7_mask[5]) );
  AND2X1_LVT csr_U2891 ( .A1(csr_n1893), .A2(io_ptw_pmp_7_addr[1]), .Y(
        io_ptw_pmp_7_mask[4]) );
  AND2X1_LVT csr_U2890 ( .A1(csr_n1892), .A2(io_ptw_pmp_7_addr[0]), .Y(
        io_ptw_pmp_7_mask[3]) );
  AND2X1_LVT csr_U2889 ( .A1(csr_n1891), .A2(io_ptw_pmp_7_addr[28]), .Y(
        io_ptw_pmp_7_mask[31]) );
  AND2X1_LVT csr_U2888 ( .A1(csr_n1890), .A2(io_ptw_pmp_7_addr[27]), .Y(
        io_ptw_pmp_7_mask[30]) );
  AND2X1_LVT csr_U2887 ( .A1(csr_n1889), .A2(io_ptw_pmp_7_addr[26]), .Y(
        io_ptw_pmp_7_mask[29]) );
  AND2X1_LVT csr_U2886 ( .A1(csr_n1888), .A2(io_ptw_pmp_7_addr[25]), .Y(
        io_ptw_pmp_7_mask[28]) );
  AND2X1_LVT csr_U2885 ( .A1(csr_n1887), .A2(io_ptw_pmp_7_addr[24]), .Y(
        io_ptw_pmp_7_mask[27]) );
  AND2X1_LVT csr_U2884 ( .A1(csr_n1886), .A2(io_ptw_pmp_7_addr[23]), .Y(
        io_ptw_pmp_7_mask[26]) );
  AND2X1_LVT csr_U2883 ( .A1(csr_n1885), .A2(io_ptw_pmp_7_addr[22]), .Y(
        io_ptw_pmp_7_mask[25]) );
  AND2X1_LVT csr_U2882 ( .A1(csr_n1884), .A2(io_ptw_pmp_7_addr[21]), .Y(
        io_ptw_pmp_7_mask[24]) );
  AND2X1_LVT csr_U2881 ( .A1(csr_n1883), .A2(io_ptw_pmp_7_addr[20]), .Y(
        io_ptw_pmp_7_mask[23]) );
  AND2X1_LVT csr_U2880 ( .A1(csr_n1882), .A2(io_ptw_pmp_7_addr[19]), .Y(
        io_ptw_pmp_7_mask[22]) );
  AND2X1_LVT csr_U2879 ( .A1(csr_n1881), .A2(io_ptw_pmp_7_addr[18]), .Y(
        io_ptw_pmp_7_mask[21]) );
  AND2X1_LVT csr_U2878 ( .A1(csr_n1880), .A2(io_ptw_pmp_7_addr[17]), .Y(
        io_ptw_pmp_7_mask[20]) );
  AND2X1_LVT csr_U2877 ( .A1(csr_n1879), .A2(io_ptw_pmp_7_addr[16]), .Y(
        io_ptw_pmp_7_mask[19]) );
  AND2X1_LVT csr_U2876 ( .A1(csr_n1878), .A2(io_ptw_pmp_7_addr[15]), .Y(
        io_ptw_pmp_7_mask[18]) );
  AND2X1_LVT csr_U2875 ( .A1(csr_n1877), .A2(io_ptw_pmp_7_addr[14]), .Y(
        io_ptw_pmp_7_mask[17]) );
  AND2X1_LVT csr_U2874 ( .A1(csr_n1876), .A2(io_ptw_pmp_7_addr[13]), .Y(
        io_ptw_pmp_7_mask[16]) );
  AND2X1_LVT csr_U2873 ( .A1(csr_n1875), .A2(io_ptw_pmp_7_addr[12]), .Y(
        io_ptw_pmp_7_mask[15]) );
  AND2X1_LVT csr_U2872 ( .A1(csr_n1874), .A2(io_ptw_pmp_7_addr[10]), .Y(
        io_ptw_pmp_7_mask[13]) );
  AND2X1_LVT csr_U2871 ( .A1(csr_n1873), .A2(io_ptw_pmp_7_addr[8]), .Y(
        io_ptw_pmp_7_mask[11]) );
  AND2X1_LVT csr_U2870 ( .A1(csr_n1872), .A2(io_ptw_pmp_6_addr[6]), .Y(
        io_ptw_pmp_6_mask[9]) );
  AND2X1_LVT csr_U2869 ( .A1(csr_n1871), .A2(io_ptw_pmp_6_addr[5]), .Y(
        io_ptw_pmp_6_mask[8]) );
  AND2X1_LVT csr_U2868 ( .A1(csr_n1870), .A2(io_ptw_pmp_6_addr[4]), .Y(
        io_ptw_pmp_6_mask[7]) );
  AND2X1_LVT csr_U2867 ( .A1(csr_n1869), .A2(io_ptw_pmp_6_addr[2]), .Y(
        io_ptw_pmp_6_mask[5]) );
  AND2X1_LVT csr_U2866 ( .A1(csr_n1868), .A2(io_ptw_pmp_6_addr[1]), .Y(
        io_ptw_pmp_6_mask[4]) );
  AND2X1_LVT csr_U2865 ( .A1(csr_n1867), .A2(io_ptw_pmp_6_addr[0]), .Y(
        io_ptw_pmp_6_mask[3]) );
  AND2X1_LVT csr_U2864 ( .A1(csr_n1866), .A2(io_ptw_pmp_6_addr[28]), .Y(
        io_ptw_pmp_6_mask[31]) );
  AND2X1_LVT csr_U2863 ( .A1(csr_n1865), .A2(io_ptw_pmp_6_addr[27]), .Y(
        io_ptw_pmp_6_mask[30]) );
  AND2X1_LVT csr_U2862 ( .A1(csr_n1864), .A2(io_ptw_pmp_6_addr[26]), .Y(
        io_ptw_pmp_6_mask[29]) );
  AND2X1_LVT csr_U2861 ( .A1(csr_n1863), .A2(io_ptw_pmp_6_addr[25]), .Y(
        io_ptw_pmp_6_mask[28]) );
  AND2X1_LVT csr_U2860 ( .A1(csr_n1862), .A2(io_ptw_pmp_6_addr[24]), .Y(
        io_ptw_pmp_6_mask[27]) );
  AND2X1_LVT csr_U2859 ( .A1(csr_n1861), .A2(io_ptw_pmp_6_addr[23]), .Y(
        io_ptw_pmp_6_mask[26]) );
  AND2X1_LVT csr_U2858 ( .A1(csr_n1860), .A2(io_ptw_pmp_6_addr[22]), .Y(
        io_ptw_pmp_6_mask[25]) );
  AND2X1_LVT csr_U2857 ( .A1(csr_n1859), .A2(io_ptw_pmp_6_addr[21]), .Y(
        io_ptw_pmp_6_mask[24]) );
  AND2X1_LVT csr_U2856 ( .A1(csr_n1858), .A2(io_ptw_pmp_6_addr[20]), .Y(
        io_ptw_pmp_6_mask[23]) );
  AND2X1_LVT csr_U2855 ( .A1(csr_n1857), .A2(io_ptw_pmp_6_addr[19]), .Y(
        io_ptw_pmp_6_mask[22]) );
  AND2X1_LVT csr_U2854 ( .A1(csr_n1856), .A2(io_ptw_pmp_6_addr[18]), .Y(
        io_ptw_pmp_6_mask[21]) );
  AND2X1_LVT csr_U2853 ( .A1(csr_n1855), .A2(io_ptw_pmp_6_addr[17]), .Y(
        io_ptw_pmp_6_mask[20]) );
  AND2X1_LVT csr_U2852 ( .A1(csr_n1854), .A2(io_ptw_pmp_6_addr[16]), .Y(
        io_ptw_pmp_6_mask[19]) );
  AND2X1_LVT csr_U2851 ( .A1(csr_n1853), .A2(io_ptw_pmp_6_addr[15]), .Y(
        io_ptw_pmp_6_mask[18]) );
  AND2X1_LVT csr_U2850 ( .A1(csr_n1852), .A2(io_ptw_pmp_6_addr[14]), .Y(
        io_ptw_pmp_6_mask[17]) );
  AND2X1_LVT csr_U2849 ( .A1(csr_n1851), .A2(io_ptw_pmp_6_addr[13]), .Y(
        io_ptw_pmp_6_mask[16]) );
  AND2X1_LVT csr_U2848 ( .A1(csr_n1850), .A2(io_ptw_pmp_6_addr[12]), .Y(
        io_ptw_pmp_6_mask[15]) );
  AND2X1_LVT csr_U2847 ( .A1(csr_n1849), .A2(io_ptw_pmp_6_addr[10]), .Y(
        io_ptw_pmp_6_mask[13]) );
  AND2X1_LVT csr_U2846 ( .A1(csr_n1848), .A2(io_ptw_pmp_6_addr[8]), .Y(
        io_ptw_pmp_6_mask[11]) );
  AND2X1_LVT csr_U2845 ( .A1(csr_n1847), .A2(io_ptw_pmp_5_addr[6]), .Y(
        io_ptw_pmp_5_mask[9]) );
  AND2X1_LVT csr_U2844 ( .A1(csr_n1846), .A2(io_ptw_pmp_5_addr[5]), .Y(
        io_ptw_pmp_5_mask[8]) );
  AND2X1_LVT csr_U2843 ( .A1(csr_n1845), .A2(io_ptw_pmp_5_addr[4]), .Y(
        io_ptw_pmp_5_mask[7]) );
  AND2X1_LVT csr_U2842 ( .A1(csr_n1844), .A2(io_ptw_pmp_5_addr[2]), .Y(
        io_ptw_pmp_5_mask[5]) );
  AND2X1_LVT csr_U2841 ( .A1(csr_n1843), .A2(io_ptw_pmp_5_addr[1]), .Y(
        io_ptw_pmp_5_mask[4]) );
  AND2X1_LVT csr_U2840 ( .A1(csr_n1842), .A2(io_ptw_pmp_5_addr[0]), .Y(
        io_ptw_pmp_5_mask[3]) );
  AND2X1_LVT csr_U2839 ( .A1(csr_n1841), .A2(io_ptw_pmp_5_addr[28]), .Y(
        io_ptw_pmp_5_mask[31]) );
  AND2X1_LVT csr_U2838 ( .A1(csr_n1840), .A2(io_ptw_pmp_5_addr[27]), .Y(
        io_ptw_pmp_5_mask[30]) );
  AND2X1_LVT csr_U2837 ( .A1(csr_n1839), .A2(io_ptw_pmp_5_addr[26]), .Y(
        io_ptw_pmp_5_mask[29]) );
  AND2X1_LVT csr_U2836 ( .A1(csr_n1838), .A2(io_ptw_pmp_5_addr[25]), .Y(
        io_ptw_pmp_5_mask[28]) );
  AND2X1_LVT csr_U2835 ( .A1(csr_n1837), .A2(io_ptw_pmp_5_addr[24]), .Y(
        io_ptw_pmp_5_mask[27]) );
  AND2X1_LVT csr_U2834 ( .A1(csr_n1836), .A2(io_ptw_pmp_5_addr[23]), .Y(
        io_ptw_pmp_5_mask[26]) );
  AND2X1_LVT csr_U2833 ( .A1(csr_n1835), .A2(io_ptw_pmp_5_addr[22]), .Y(
        io_ptw_pmp_5_mask[25]) );
  AND2X1_LVT csr_U2832 ( .A1(csr_n1834), .A2(io_ptw_pmp_5_addr[21]), .Y(
        io_ptw_pmp_5_mask[24]) );
  AND2X1_LVT csr_U2831 ( .A1(csr_n1833), .A2(io_ptw_pmp_5_addr[20]), .Y(
        io_ptw_pmp_5_mask[23]) );
  AND2X1_LVT csr_U2830 ( .A1(csr_n1832), .A2(io_ptw_pmp_5_addr[19]), .Y(
        io_ptw_pmp_5_mask[22]) );
  AND2X1_LVT csr_U2829 ( .A1(csr_n1831), .A2(io_ptw_pmp_5_addr[18]), .Y(
        io_ptw_pmp_5_mask[21]) );
  AND2X1_LVT csr_U2828 ( .A1(csr_n1830), .A2(io_ptw_pmp_5_addr[17]), .Y(
        io_ptw_pmp_5_mask[20]) );
  AND2X1_LVT csr_U2827 ( .A1(csr_n1829), .A2(io_ptw_pmp_5_addr[16]), .Y(
        io_ptw_pmp_5_mask[19]) );
  AND2X1_LVT csr_U2826 ( .A1(csr_n1828), .A2(io_ptw_pmp_5_addr[15]), .Y(
        io_ptw_pmp_5_mask[18]) );
  AND2X1_LVT csr_U2825 ( .A1(csr_n1827), .A2(io_ptw_pmp_5_addr[14]), .Y(
        io_ptw_pmp_5_mask[17]) );
  AND2X1_LVT csr_U2824 ( .A1(csr_n1826), .A2(io_ptw_pmp_5_addr[13]), .Y(
        io_ptw_pmp_5_mask[16]) );
  AND2X1_LVT csr_U2823 ( .A1(csr_n1825), .A2(io_ptw_pmp_5_addr[12]), .Y(
        io_ptw_pmp_5_mask[15]) );
  AND2X1_LVT csr_U2822 ( .A1(csr_n1824), .A2(io_ptw_pmp_5_addr[10]), .Y(
        io_ptw_pmp_5_mask[13]) );
  AND2X1_LVT csr_U2821 ( .A1(csr_n1823), .A2(io_ptw_pmp_5_addr[8]), .Y(
        io_ptw_pmp_5_mask[11]) );
  AND2X1_LVT csr_U2820 ( .A1(csr_n1822), .A2(io_ptw_pmp_4_addr[6]), .Y(
        io_ptw_pmp_4_mask[9]) );
  AND2X1_LVT csr_U2819 ( .A1(csr_n1821), .A2(io_ptw_pmp_4_addr[5]), .Y(
        io_ptw_pmp_4_mask[8]) );
  AND2X1_LVT csr_U2818 ( .A1(csr_n1820), .A2(io_ptw_pmp_4_addr[4]), .Y(
        io_ptw_pmp_4_mask[7]) );
  AND2X1_LVT csr_U2817 ( .A1(csr_n1819), .A2(io_ptw_pmp_4_addr[2]), .Y(
        io_ptw_pmp_4_mask[5]) );
  AND2X1_LVT csr_U2816 ( .A1(csr_n1818), .A2(io_ptw_pmp_4_addr[1]), .Y(
        io_ptw_pmp_4_mask[4]) );
  AND2X1_LVT csr_U2815 ( .A1(csr_n1817), .A2(io_ptw_pmp_4_addr[0]), .Y(
        io_ptw_pmp_4_mask[3]) );
  AND2X1_LVT csr_U2814 ( .A1(csr_n1816), .A2(io_ptw_pmp_4_addr[28]), .Y(
        io_ptw_pmp_4_mask[31]) );
  AND2X1_LVT csr_U2813 ( .A1(csr_n1815), .A2(io_ptw_pmp_4_addr[27]), .Y(
        io_ptw_pmp_4_mask[30]) );
  AND2X1_LVT csr_U2812 ( .A1(csr_n1814), .A2(io_ptw_pmp_4_addr[26]), .Y(
        io_ptw_pmp_4_mask[29]) );
  AND2X1_LVT csr_U2811 ( .A1(csr_n1813), .A2(io_ptw_pmp_4_addr[25]), .Y(
        io_ptw_pmp_4_mask[28]) );
  AND2X1_LVT csr_U2810 ( .A1(csr_n1812), .A2(io_ptw_pmp_4_addr[24]), .Y(
        io_ptw_pmp_4_mask[27]) );
  AND2X1_LVT csr_U2809 ( .A1(csr_n1811), .A2(io_ptw_pmp_4_addr[23]), .Y(
        io_ptw_pmp_4_mask[26]) );
  AND2X1_LVT csr_U2808 ( .A1(csr_n1810), .A2(io_ptw_pmp_4_addr[22]), .Y(
        io_ptw_pmp_4_mask[25]) );
  AND2X1_LVT csr_U2807 ( .A1(csr_n1809), .A2(io_ptw_pmp_4_addr[21]), .Y(
        io_ptw_pmp_4_mask[24]) );
  AND2X1_LVT csr_U2806 ( .A1(csr_n1808), .A2(io_ptw_pmp_4_addr[20]), .Y(
        io_ptw_pmp_4_mask[23]) );
  AND2X1_LVT csr_U2805 ( .A1(csr_n1807), .A2(io_ptw_pmp_4_addr[19]), .Y(
        io_ptw_pmp_4_mask[22]) );
  AND2X1_LVT csr_U2804 ( .A1(csr_n1806), .A2(io_ptw_pmp_4_addr[18]), .Y(
        io_ptw_pmp_4_mask[21]) );
  AND2X1_LVT csr_U2803 ( .A1(csr_n1805), .A2(io_ptw_pmp_4_addr[17]), .Y(
        io_ptw_pmp_4_mask[20]) );
  AND2X1_LVT csr_U2802 ( .A1(csr_n1804), .A2(io_ptw_pmp_4_addr[16]), .Y(
        io_ptw_pmp_4_mask[19]) );
  AND2X1_LVT csr_U2801 ( .A1(csr_n1803), .A2(io_ptw_pmp_4_addr[15]), .Y(
        io_ptw_pmp_4_mask[18]) );
  AND2X1_LVT csr_U2800 ( .A1(csr_n1802), .A2(io_ptw_pmp_4_addr[14]), .Y(
        io_ptw_pmp_4_mask[17]) );
  AND2X1_LVT csr_U2799 ( .A1(csr_n1801), .A2(io_ptw_pmp_4_addr[13]), .Y(
        io_ptw_pmp_4_mask[16]) );
  AND2X1_LVT csr_U2798 ( .A1(csr_n1800), .A2(io_ptw_pmp_4_addr[12]), .Y(
        io_ptw_pmp_4_mask[15]) );
  AND2X1_LVT csr_U2797 ( .A1(csr_n1799), .A2(io_ptw_pmp_4_addr[10]), .Y(
        io_ptw_pmp_4_mask[13]) );
  AND2X1_LVT csr_U2796 ( .A1(csr_n1798), .A2(io_ptw_pmp_4_addr[8]), .Y(
        io_ptw_pmp_4_mask[11]) );
  AND2X1_LVT csr_U2795 ( .A1(csr_n1797), .A2(io_ptw_pmp_3_addr[6]), .Y(
        io_ptw_pmp_3_mask[9]) );
  AND2X1_LVT csr_U2794 ( .A1(csr_n1796), .A2(io_ptw_pmp_3_addr[5]), .Y(
        io_ptw_pmp_3_mask[8]) );
  AND2X1_LVT csr_U2793 ( .A1(csr_n1795), .A2(io_ptw_pmp_3_addr[4]), .Y(
        io_ptw_pmp_3_mask[7]) );
  AND2X1_LVT csr_U2792 ( .A1(csr_n1794), .A2(io_ptw_pmp_3_addr[2]), .Y(
        io_ptw_pmp_3_mask[5]) );
  AND2X1_LVT csr_U2791 ( .A1(csr_n1793), .A2(io_ptw_pmp_3_addr[1]), .Y(
        io_ptw_pmp_3_mask[4]) );
  AND2X1_LVT csr_U2790 ( .A1(csr_n1792), .A2(io_ptw_pmp_3_addr[0]), .Y(
        io_ptw_pmp_3_mask[3]) );
  AND2X1_LVT csr_U2789 ( .A1(csr_n1791), .A2(io_ptw_pmp_3_addr[28]), .Y(
        io_ptw_pmp_3_mask[31]) );
  AND2X1_LVT csr_U2788 ( .A1(csr_n1790), .A2(io_ptw_pmp_3_addr[27]), .Y(
        io_ptw_pmp_3_mask[30]) );
  AND2X1_LVT csr_U2787 ( .A1(csr_n1789), .A2(io_ptw_pmp_3_addr[26]), .Y(
        io_ptw_pmp_3_mask[29]) );
  AND2X1_LVT csr_U2786 ( .A1(csr_n1788), .A2(io_ptw_pmp_3_addr[25]), .Y(
        io_ptw_pmp_3_mask[28]) );
  AND2X1_LVT csr_U2785 ( .A1(csr_n1787), .A2(io_ptw_pmp_3_addr[24]), .Y(
        io_ptw_pmp_3_mask[27]) );
  AND2X1_LVT csr_U2784 ( .A1(csr_n1786), .A2(io_ptw_pmp_3_addr[23]), .Y(
        io_ptw_pmp_3_mask[26]) );
  AND2X1_LVT csr_U2783 ( .A1(csr_n1785), .A2(io_ptw_pmp_3_addr[22]), .Y(
        io_ptw_pmp_3_mask[25]) );
  AND2X1_LVT csr_U2782 ( .A1(csr_n1784), .A2(io_ptw_pmp_3_addr[21]), .Y(
        io_ptw_pmp_3_mask[24]) );
  AND2X1_LVT csr_U2781 ( .A1(csr_n1783), .A2(io_ptw_pmp_3_addr[20]), .Y(
        io_ptw_pmp_3_mask[23]) );
  AND2X1_LVT csr_U2780 ( .A1(csr_n1782), .A2(io_ptw_pmp_3_addr[19]), .Y(
        io_ptw_pmp_3_mask[22]) );
  AND2X1_LVT csr_U2779 ( .A1(csr_n1781), .A2(io_ptw_pmp_3_addr[18]), .Y(
        io_ptw_pmp_3_mask[21]) );
  AND2X1_LVT csr_U2778 ( .A1(csr_n1780), .A2(io_ptw_pmp_3_addr[17]), .Y(
        io_ptw_pmp_3_mask[20]) );
  AND2X1_LVT csr_U2777 ( .A1(csr_n1779), .A2(io_ptw_pmp_3_addr[16]), .Y(
        io_ptw_pmp_3_mask[19]) );
  AND2X1_LVT csr_U2776 ( .A1(csr_n1778), .A2(io_ptw_pmp_3_addr[15]), .Y(
        io_ptw_pmp_3_mask[18]) );
  AND2X1_LVT csr_U2775 ( .A1(csr_n1777), .A2(io_ptw_pmp_3_addr[14]), .Y(
        io_ptw_pmp_3_mask[17]) );
  AND2X1_LVT csr_U2774 ( .A1(csr_n1776), .A2(io_ptw_pmp_3_addr[13]), .Y(
        io_ptw_pmp_3_mask[16]) );
  AND2X1_LVT csr_U2773 ( .A1(csr_n1775), .A2(io_ptw_pmp_3_addr[12]), .Y(
        io_ptw_pmp_3_mask[15]) );
  AND2X1_LVT csr_U2772 ( .A1(csr_n1774), .A2(io_ptw_pmp_3_addr[10]), .Y(
        io_ptw_pmp_3_mask[13]) );
  AND2X1_LVT csr_U2771 ( .A1(csr_n1773), .A2(io_ptw_pmp_3_addr[8]), .Y(
        io_ptw_pmp_3_mask[11]) );
  AND2X1_LVT csr_U2770 ( .A1(csr_n1772), .A2(io_ptw_pmp_2_addr[6]), .Y(
        io_ptw_pmp_2_mask[9]) );
  AND2X1_LVT csr_U2769 ( .A1(csr_n1771), .A2(io_ptw_pmp_2_addr[5]), .Y(
        io_ptw_pmp_2_mask[8]) );
  AND2X1_LVT csr_U2768 ( .A1(csr_n1770), .A2(io_ptw_pmp_2_addr[4]), .Y(
        io_ptw_pmp_2_mask[7]) );
  AND2X1_LVT csr_U2767 ( .A1(csr_n1769), .A2(io_ptw_pmp_2_addr[2]), .Y(
        io_ptw_pmp_2_mask[5]) );
  AND2X1_LVT csr_U2766 ( .A1(csr_n1768), .A2(io_ptw_pmp_2_addr[1]), .Y(
        io_ptw_pmp_2_mask[4]) );
  AND2X1_LVT csr_U2765 ( .A1(csr_n1767), .A2(io_ptw_pmp_2_addr[0]), .Y(
        io_ptw_pmp_2_mask[3]) );
  AND2X1_LVT csr_U2764 ( .A1(csr_n1766), .A2(io_ptw_pmp_2_addr[28]), .Y(
        io_ptw_pmp_2_mask[31]) );
  AND2X1_LVT csr_U2763 ( .A1(csr_n1765), .A2(io_ptw_pmp_2_addr[27]), .Y(
        io_ptw_pmp_2_mask[30]) );
  AND2X1_LVT csr_U2762 ( .A1(csr_n1764), .A2(io_ptw_pmp_2_addr[26]), .Y(
        io_ptw_pmp_2_mask[29]) );
  AND2X1_LVT csr_U2761 ( .A1(csr_n1763), .A2(io_ptw_pmp_2_addr[25]), .Y(
        io_ptw_pmp_2_mask[28]) );
  AND2X1_LVT csr_U2760 ( .A1(csr_n1762), .A2(io_ptw_pmp_2_addr[24]), .Y(
        io_ptw_pmp_2_mask[27]) );
  AND2X1_LVT csr_U2759 ( .A1(csr_n1761), .A2(io_ptw_pmp_2_addr[23]), .Y(
        io_ptw_pmp_2_mask[26]) );
  AND2X1_LVT csr_U2758 ( .A1(csr_n1760), .A2(io_ptw_pmp_2_addr[22]), .Y(
        io_ptw_pmp_2_mask[25]) );
  AND2X1_LVT csr_U2757 ( .A1(csr_n1759), .A2(io_ptw_pmp_2_addr[21]), .Y(
        io_ptw_pmp_2_mask[24]) );
  AND2X1_LVT csr_U2756 ( .A1(csr_n1758), .A2(io_ptw_pmp_2_addr[20]), .Y(
        io_ptw_pmp_2_mask[23]) );
  AND2X1_LVT csr_U2755 ( .A1(csr_n1757), .A2(io_ptw_pmp_2_addr[19]), .Y(
        io_ptw_pmp_2_mask[22]) );
  AND2X1_LVT csr_U2754 ( .A1(csr_n1756), .A2(io_ptw_pmp_2_addr[18]), .Y(
        io_ptw_pmp_2_mask[21]) );
  AND2X1_LVT csr_U2753 ( .A1(csr_n1755), .A2(io_ptw_pmp_2_addr[17]), .Y(
        io_ptw_pmp_2_mask[20]) );
  AND2X1_LVT csr_U2752 ( .A1(csr_n1754), .A2(io_ptw_pmp_2_addr[16]), .Y(
        io_ptw_pmp_2_mask[19]) );
  AND2X1_LVT csr_U2751 ( .A1(csr_n1753), .A2(io_ptw_pmp_2_addr[15]), .Y(
        io_ptw_pmp_2_mask[18]) );
  AND2X1_LVT csr_U2750 ( .A1(csr_n1752), .A2(io_ptw_pmp_2_addr[14]), .Y(
        io_ptw_pmp_2_mask[17]) );
  AND2X1_LVT csr_U2749 ( .A1(csr_n1751), .A2(io_ptw_pmp_2_addr[13]), .Y(
        io_ptw_pmp_2_mask[16]) );
  AND2X1_LVT csr_U2748 ( .A1(csr_n1750), .A2(io_ptw_pmp_2_addr[12]), .Y(
        io_ptw_pmp_2_mask[15]) );
  AND2X1_LVT csr_U2747 ( .A1(csr_n1749), .A2(io_ptw_pmp_2_addr[10]), .Y(
        io_ptw_pmp_2_mask[13]) );
  AND2X1_LVT csr_U2746 ( .A1(csr_n1748), .A2(io_ptw_pmp_2_addr[8]), .Y(
        io_ptw_pmp_2_mask[11]) );
  AND2X1_LVT csr_U2745 ( .A1(csr_n1747), .A2(io_ptw_pmp_1_addr[6]), .Y(
        io_ptw_pmp_1_mask[9]) );
  AND2X1_LVT csr_U2744 ( .A1(csr_n1746), .A2(io_ptw_pmp_1_addr[5]), .Y(
        io_ptw_pmp_1_mask[8]) );
  AND2X1_LVT csr_U2743 ( .A1(csr_n1745), .A2(io_ptw_pmp_1_addr[4]), .Y(
        io_ptw_pmp_1_mask[7]) );
  AND2X1_LVT csr_U2742 ( .A1(csr_n1744), .A2(io_ptw_pmp_1_addr[2]), .Y(
        io_ptw_pmp_1_mask[5]) );
  AND2X1_LVT csr_U2741 ( .A1(csr_n1743), .A2(io_ptw_pmp_1_addr[1]), .Y(
        io_ptw_pmp_1_mask[4]) );
  AND2X1_LVT csr_U2740 ( .A1(csr_n1742), .A2(io_ptw_pmp_1_addr[0]), .Y(
        io_ptw_pmp_1_mask[3]) );
  AND2X1_LVT csr_U2739 ( .A1(csr_n1741), .A2(io_ptw_pmp_1_addr[28]), .Y(
        io_ptw_pmp_1_mask[31]) );
  AND2X1_LVT csr_U2738 ( .A1(csr_n1740), .A2(io_ptw_pmp_1_addr[27]), .Y(
        io_ptw_pmp_1_mask[30]) );
  AND2X1_LVT csr_U2737 ( .A1(csr_n1739), .A2(io_ptw_pmp_1_addr[26]), .Y(
        io_ptw_pmp_1_mask[29]) );
  AND2X1_LVT csr_U2736 ( .A1(csr_n1738), .A2(io_ptw_pmp_1_addr[25]), .Y(
        io_ptw_pmp_1_mask[28]) );
  AND2X1_LVT csr_U2735 ( .A1(csr_n1737), .A2(io_ptw_pmp_1_addr[24]), .Y(
        io_ptw_pmp_1_mask[27]) );
  AND2X1_LVT csr_U2734 ( .A1(csr_n1736), .A2(io_ptw_pmp_1_addr[23]), .Y(
        io_ptw_pmp_1_mask[26]) );
  AND2X1_LVT csr_U2733 ( .A1(csr_n1735), .A2(io_ptw_pmp_1_addr[22]), .Y(
        io_ptw_pmp_1_mask[25]) );
  AND2X1_LVT csr_U2732 ( .A1(csr_n1734), .A2(io_ptw_pmp_1_addr[21]), .Y(
        io_ptw_pmp_1_mask[24]) );
  AND2X1_LVT csr_U2731 ( .A1(csr_n1733), .A2(io_ptw_pmp_1_addr[20]), .Y(
        io_ptw_pmp_1_mask[23]) );
  AND2X1_LVT csr_U2730 ( .A1(csr_n1732), .A2(io_ptw_pmp_1_addr[19]), .Y(
        io_ptw_pmp_1_mask[22]) );
  AND2X1_LVT csr_U2729 ( .A1(csr_n1731), .A2(io_ptw_pmp_1_addr[18]), .Y(
        io_ptw_pmp_1_mask[21]) );
  AND2X1_LVT csr_U2728 ( .A1(csr_n1730), .A2(io_ptw_pmp_1_addr[17]), .Y(
        io_ptw_pmp_1_mask[20]) );
  AND2X1_LVT csr_U2727 ( .A1(csr_n1729), .A2(io_ptw_pmp_1_addr[16]), .Y(
        io_ptw_pmp_1_mask[19]) );
  AND2X1_LVT csr_U2726 ( .A1(csr_n1728), .A2(io_ptw_pmp_1_addr[15]), .Y(
        io_ptw_pmp_1_mask[18]) );
  AND2X1_LVT csr_U2725 ( .A1(csr_n1727), .A2(io_ptw_pmp_1_addr[14]), .Y(
        io_ptw_pmp_1_mask[17]) );
  AND2X1_LVT csr_U2724 ( .A1(csr_n1726), .A2(io_ptw_pmp_1_addr[13]), .Y(
        io_ptw_pmp_1_mask[16]) );
  AND2X1_LVT csr_U2723 ( .A1(csr_n1725), .A2(io_ptw_pmp_1_addr[12]), .Y(
        io_ptw_pmp_1_mask[15]) );
  AND2X1_LVT csr_U2722 ( .A1(csr_n1724), .A2(io_ptw_pmp_1_addr[10]), .Y(
        io_ptw_pmp_1_mask[13]) );
  AND2X1_LVT csr_U2721 ( .A1(csr_n1723), .A2(io_ptw_pmp_1_addr[8]), .Y(
        io_ptw_pmp_1_mask[11]) );
  AND2X1_LVT csr_U2720 ( .A1(csr_n1722), .A2(io_ptw_pmp_0_addr[6]), .Y(
        io_ptw_pmp_0_mask[9]) );
  AND2X1_LVT csr_U2719 ( .A1(csr_n1721), .A2(io_ptw_pmp_0_addr[5]), .Y(
        io_ptw_pmp_0_mask[8]) );
  AND2X1_LVT csr_U2718 ( .A1(csr_n1720), .A2(io_ptw_pmp_0_addr[4]), .Y(
        io_ptw_pmp_0_mask[7]) );
  AND2X1_LVT csr_U2717 ( .A1(csr_n1719), .A2(io_ptw_pmp_0_addr[2]), .Y(
        io_ptw_pmp_0_mask[5]) );
  AND2X1_LVT csr_U2716 ( .A1(csr_n1718), .A2(io_ptw_pmp_0_addr[1]), .Y(
        io_ptw_pmp_0_mask[4]) );
  AND2X1_LVT csr_U2715 ( .A1(csr_n1717), .A2(io_ptw_pmp_0_addr[0]), .Y(
        io_ptw_pmp_0_mask[3]) );
  AND2X1_LVT csr_U2714 ( .A1(csr_n1716), .A2(io_ptw_pmp_0_addr[28]), .Y(
        io_ptw_pmp_0_mask[31]) );
  AND2X1_LVT csr_U2713 ( .A1(csr_n1715), .A2(io_ptw_pmp_0_addr[27]), .Y(
        io_ptw_pmp_0_mask[30]) );
  AND2X1_LVT csr_U2712 ( .A1(csr_n1714), .A2(io_ptw_pmp_0_addr[26]), .Y(
        io_ptw_pmp_0_mask[29]) );
  AND2X1_LVT csr_U2711 ( .A1(csr_n1713), .A2(io_ptw_pmp_0_addr[25]), .Y(
        io_ptw_pmp_0_mask[28]) );
  AND2X1_LVT csr_U2710 ( .A1(csr_n1712), .A2(io_ptw_pmp_0_addr[24]), .Y(
        io_ptw_pmp_0_mask[27]) );
  AND2X1_LVT csr_U2709 ( .A1(csr_n1711), .A2(io_ptw_pmp_0_addr[23]), .Y(
        io_ptw_pmp_0_mask[26]) );
  AND2X1_LVT csr_U2708 ( .A1(csr_n1710), .A2(io_ptw_pmp_0_addr[22]), .Y(
        io_ptw_pmp_0_mask[25]) );
  AND2X1_LVT csr_U2707 ( .A1(csr_n1709), .A2(io_ptw_pmp_0_addr[21]), .Y(
        io_ptw_pmp_0_mask[24]) );
  AND2X1_LVT csr_U2706 ( .A1(csr_n1708), .A2(io_ptw_pmp_0_addr[20]), .Y(
        io_ptw_pmp_0_mask[23]) );
  AND2X1_LVT csr_U2705 ( .A1(csr_n1707), .A2(io_ptw_pmp_0_addr[19]), .Y(
        io_ptw_pmp_0_mask[22]) );
  AND2X1_LVT csr_U2704 ( .A1(csr_n1706), .A2(io_ptw_pmp_0_addr[18]), .Y(
        io_ptw_pmp_0_mask[21]) );
  AND2X1_LVT csr_U2703 ( .A1(csr_n1705), .A2(io_ptw_pmp_0_addr[17]), .Y(
        io_ptw_pmp_0_mask[20]) );
  AND2X1_LVT csr_U2702 ( .A1(csr_n1704), .A2(io_ptw_pmp_0_addr[16]), .Y(
        io_ptw_pmp_0_mask[19]) );
  AND2X1_LVT csr_U2701 ( .A1(csr_n1703), .A2(io_ptw_pmp_0_addr[15]), .Y(
        io_ptw_pmp_0_mask[18]) );
  AND2X1_LVT csr_U2700 ( .A1(csr_n1702), .A2(io_ptw_pmp_0_addr[14]), .Y(
        io_ptw_pmp_0_mask[17]) );
  AND2X1_LVT csr_U2699 ( .A1(csr_n1701), .A2(io_ptw_pmp_0_addr[13]), .Y(
        io_ptw_pmp_0_mask[16]) );
  AND2X1_LVT csr_U2698 ( .A1(csr_n1700), .A2(io_ptw_pmp_0_addr[12]), .Y(
        io_ptw_pmp_0_mask[15]) );
  AND2X1_LVT csr_U2697 ( .A1(csr_n1699), .A2(io_ptw_pmp_0_addr[10]), .Y(
        io_ptw_pmp_0_mask[13]) );
  AND2X1_LVT csr_U2696 ( .A1(csr_n1698), .A2(io_ptw_pmp_0_addr[8]), .Y(
        io_ptw_pmp_0_mask[11]) );
  AO22X1_LVT csr_U2695 ( .A1(csr_n512), .A2(csr_wdata_8_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[8]), .Y(csr_n_GEN_307[8]) );
  AO22X1_LVT csr_U2694 ( .A1(csr_n512), .A2(csr_wdata_6_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[6]), .Y(csr_n_GEN_307[6]) );
  AO22X1_LVT csr_U2693 ( .A1(csr_n512), .A2(csr_wdata_5_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[5]), .Y(csr_n_GEN_307[5]) );
  AO22X1_LVT csr_U2692 ( .A1(csr_n512), .A2(csr_wdata_4_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[4]), .Y(csr_n_GEN_307[4]) );
  AO22X1_LVT csr_U2691 ( .A1(csr_n512), .A2(csr_wdata_2_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[2]), .Y(csr_n_GEN_307[2]) );
  AO22X1_LVT csr_U2690 ( .A1(csr_n512), .A2(csr_wdata_29_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[29]), .Y(csr_n_GEN_307[29]) );
  AO22X1_LVT csr_U2689 ( .A1(csr_n512), .A2(csr_wdata_28_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[28]), .Y(csr_n_GEN_307[28]) );
  AO22X1_LVT csr_U2688 ( .A1(csr_n512), .A2(csr_wdata_27_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[27]), .Y(csr_n_GEN_307[27]) );
  AO22X1_LVT csr_U2687 ( .A1(csr_n512), .A2(csr_wdata_26_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[26]), .Y(csr_n_GEN_307[26]) );
  AO22X1_LVT csr_U2686 ( .A1(csr_n512), .A2(csr_wdata_25_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[25]), .Y(csr_n_GEN_307[25]) );
  AO22X1_LVT csr_U2685 ( .A1(csr_n512), .A2(csr_wdata_24_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[24]), .Y(csr_n_GEN_307[24]) );
  AO22X1_LVT csr_U2684 ( .A1(csr_n512), .A2(csr_wdata_23_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[23]), .Y(csr_n_GEN_307[23]) );
  AO22X1_LVT csr_U2683 ( .A1(csr_n512), .A2(csr_wdata_22_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[22]), .Y(csr_n_GEN_307[22]) );
  AO22X1_LVT csr_U2682 ( .A1(csr_n512), .A2(csr_wdata_21_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[21]), .Y(csr_n_GEN_307[21]) );
  AO22X1_LVT csr_U2681 ( .A1(csr_n512), .A2(csr_wdata_20_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[20]), .Y(csr_n_GEN_307[20]) );
  AO22X1_LVT csr_U2680 ( .A1(csr_n512), .A2(csr_wdata_1_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[1]), .Y(csr_n_GEN_307[1]) );
  AO22X1_LVT csr_U2679 ( .A1(csr_n512), .A2(csr_wdata_19_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[19]), .Y(csr_n_GEN_307[19]) );
  AO22X1_LVT csr_U2678 ( .A1(csr_n512), .A2(csr_wdata_18_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[18]), .Y(csr_n_GEN_307[18]) );
  AO22X1_LVT csr_U2677 ( .A1(csr_n512), .A2(csr_wdata_17_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[17]), .Y(csr_n_GEN_307[17]) );
  AO22X1_LVT csr_U2676 ( .A1(csr_n512), .A2(csr_wdata_16_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[16]), .Y(csr_n_GEN_307[16]) );
  AO22X1_LVT csr_U2675 ( .A1(csr_n512), .A2(csr_wdata_15_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[15]), .Y(csr_n_GEN_307[15]) );
  AO22X1_LVT csr_U2674 ( .A1(csr_n512), .A2(csr_wdata_14_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[14]), .Y(csr_n_GEN_307[14]) );
  AO22X1_LVT csr_U2673 ( .A1(csr_n512), .A2(csr_wdata_13_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[13]), .Y(csr_n_GEN_307[13]) );
  AO22X1_LVT csr_U2672 ( .A1(csr_n512), .A2(csr_wdata_12_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[12]), .Y(csr_n_GEN_307[12]) );
  AO22X1_LVT csr_U2671 ( .A1(csr_n512), .A2(csr_wdata_10_), .A3(csr_n386), 
        .A4(io_ptw_pmp_7_addr[10]), .Y(csr_n_GEN_307[10]) );
  AO22X1_LVT csr_U2670 ( .A1(csr_n512), .A2(csr_wdata_0_), .A3(csr_n386), .A4(
        io_ptw_pmp_7_addr[0]), .Y(csr_n_GEN_307[0]) );
  AO22X1_LVT csr_U2669 ( .A1(csr_n511), .A2(csr_wdata_8_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[8]), .Y(csr_n_GEN_300[8]) );
  AO22X1_LVT csr_U2668 ( .A1(csr_n511), .A2(csr_wdata_6_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[6]), .Y(csr_n_GEN_300[6]) );
  AO22X1_LVT csr_U2667 ( .A1(csr_n511), .A2(csr_wdata_5_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[5]), .Y(csr_n_GEN_300[5]) );
  AO22X1_LVT csr_U2666 ( .A1(csr_n511), .A2(csr_wdata_4_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[4]), .Y(csr_n_GEN_300[4]) );
  AO22X1_LVT csr_U2665 ( .A1(csr_n511), .A2(csr_wdata_2_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[2]), .Y(csr_n_GEN_300[2]) );
  AO22X1_LVT csr_U2664 ( .A1(csr_n511), .A2(csr_wdata_29_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[29]), .Y(csr_n_GEN_300[29]) );
  AO22X1_LVT csr_U2663 ( .A1(csr_n511), .A2(csr_wdata_28_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[28]), .Y(csr_n_GEN_300[28]) );
  AO22X1_LVT csr_U2662 ( .A1(csr_n511), .A2(csr_wdata_27_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[27]), .Y(csr_n_GEN_300[27]) );
  AO22X1_LVT csr_U2661 ( .A1(csr_n511), .A2(csr_wdata_26_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[26]), .Y(csr_n_GEN_300[26]) );
  AO22X1_LVT csr_U2660 ( .A1(csr_n511), .A2(csr_wdata_25_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[25]), .Y(csr_n_GEN_300[25]) );
  AO22X1_LVT csr_U2659 ( .A1(csr_n511), .A2(csr_wdata_24_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[24]), .Y(csr_n_GEN_300[24]) );
  AO22X1_LVT csr_U2658 ( .A1(csr_n511), .A2(csr_wdata_23_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[23]), .Y(csr_n_GEN_300[23]) );
  AO22X1_LVT csr_U2657 ( .A1(csr_n511), .A2(csr_wdata_22_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[22]), .Y(csr_n_GEN_300[22]) );
  AO22X1_LVT csr_U2656 ( .A1(csr_n511), .A2(csr_wdata_21_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[21]), .Y(csr_n_GEN_300[21]) );
  AO22X1_LVT csr_U2655 ( .A1(csr_n511), .A2(csr_wdata_20_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[20]), .Y(csr_n_GEN_300[20]) );
  AO22X1_LVT csr_U2654 ( .A1(csr_n511), .A2(csr_wdata_1_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[1]), .Y(csr_n_GEN_300[1]) );
  AO22X1_LVT csr_U2653 ( .A1(csr_n511), .A2(csr_wdata_19_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[19]), .Y(csr_n_GEN_300[19]) );
  AO22X1_LVT csr_U2652 ( .A1(csr_n511), .A2(csr_wdata_18_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[18]), .Y(csr_n_GEN_300[18]) );
  AO22X1_LVT csr_U2651 ( .A1(csr_n511), .A2(csr_wdata_17_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[17]), .Y(csr_n_GEN_300[17]) );
  AO22X1_LVT csr_U2650 ( .A1(csr_n511), .A2(csr_wdata_16_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[16]), .Y(csr_n_GEN_300[16]) );
  AO22X1_LVT csr_U2649 ( .A1(csr_n511), .A2(csr_wdata_15_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[15]), .Y(csr_n_GEN_300[15]) );
  AO22X1_LVT csr_U2648 ( .A1(csr_n511), .A2(csr_wdata_14_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[14]), .Y(csr_n_GEN_300[14]) );
  AO22X1_LVT csr_U2647 ( .A1(csr_n511), .A2(csr_wdata_13_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[13]), .Y(csr_n_GEN_300[13]) );
  AO22X1_LVT csr_U2646 ( .A1(csr_n511), .A2(csr_wdata_12_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[12]), .Y(csr_n_GEN_300[12]) );
  AO22X1_LVT csr_U2645 ( .A1(csr_n511), .A2(csr_wdata_10_), .A3(csr_n435), 
        .A4(io_ptw_pmp_6_addr[10]), .Y(csr_n_GEN_300[10]) );
  AO22X1_LVT csr_U2644 ( .A1(csr_n511), .A2(csr_wdata_0_), .A3(csr_n435), .A4(
        io_ptw_pmp_6_addr[0]), .Y(csr_n_GEN_300[0]) );
  AO22X1_LVT csr_U2643 ( .A1(csr_n510), .A2(csr_wdata_8_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[8]), .Y(csr_n_GEN_293[8]) );
  AO22X1_LVT csr_U2642 ( .A1(csr_n510), .A2(csr_wdata_6_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[6]), .Y(csr_n_GEN_293[6]) );
  AO22X1_LVT csr_U2641 ( .A1(csr_n510), .A2(csr_wdata_5_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[5]), .Y(csr_n_GEN_293[5]) );
  AO22X1_LVT csr_U2640 ( .A1(csr_n510), .A2(csr_wdata_4_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[4]), .Y(csr_n_GEN_293[4]) );
  AO22X1_LVT csr_U2639 ( .A1(csr_n510), .A2(csr_wdata_2_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[2]), .Y(csr_n_GEN_293[2]) );
  AO22X1_LVT csr_U2638 ( .A1(csr_n510), .A2(csr_wdata_29_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[29]), .Y(csr_n_GEN_293[29]) );
  AO22X1_LVT csr_U2637 ( .A1(csr_n510), .A2(csr_wdata_28_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[28]), .Y(csr_n_GEN_293[28]) );
  AO22X1_LVT csr_U2636 ( .A1(csr_n510), .A2(csr_wdata_27_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[27]), .Y(csr_n_GEN_293[27]) );
  AO22X1_LVT csr_U2635 ( .A1(csr_n510), .A2(csr_wdata_26_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[26]), .Y(csr_n_GEN_293[26]) );
  AO22X1_LVT csr_U2634 ( .A1(csr_n510), .A2(csr_wdata_25_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[25]), .Y(csr_n_GEN_293[25]) );
  AO22X1_LVT csr_U2633 ( .A1(csr_n510), .A2(csr_wdata_24_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[24]), .Y(csr_n_GEN_293[24]) );
  AO22X1_LVT csr_U2632 ( .A1(csr_n510), .A2(csr_wdata_23_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[23]), .Y(csr_n_GEN_293[23]) );
  AO22X1_LVT csr_U2631 ( .A1(csr_n510), .A2(csr_wdata_22_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[22]), .Y(csr_n_GEN_293[22]) );
  AO22X1_LVT csr_U2630 ( .A1(csr_n510), .A2(csr_wdata_21_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[21]), .Y(csr_n_GEN_293[21]) );
  AO22X1_LVT csr_U2629 ( .A1(csr_n510), .A2(csr_wdata_20_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[20]), .Y(csr_n_GEN_293[20]) );
  AO22X1_LVT csr_U2628 ( .A1(csr_n510), .A2(csr_wdata_1_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[1]), .Y(csr_n_GEN_293[1]) );
  AO22X1_LVT csr_U2627 ( .A1(csr_n510), .A2(csr_wdata_19_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[19]), .Y(csr_n_GEN_293[19]) );
  AO22X1_LVT csr_U2626 ( .A1(csr_n510), .A2(csr_wdata_18_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[18]), .Y(csr_n_GEN_293[18]) );
  AO22X1_LVT csr_U2625 ( .A1(csr_n510), .A2(csr_wdata_17_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[17]), .Y(csr_n_GEN_293[17]) );
  AO22X1_LVT csr_U2624 ( .A1(csr_n510), .A2(csr_wdata_16_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[16]), .Y(csr_n_GEN_293[16]) );
  AO22X1_LVT csr_U2623 ( .A1(csr_n510), .A2(csr_wdata_15_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[15]), .Y(csr_n_GEN_293[15]) );
  AO22X1_LVT csr_U2622 ( .A1(csr_n510), .A2(csr_wdata_14_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[14]), .Y(csr_n_GEN_293[14]) );
  AO22X1_LVT csr_U2621 ( .A1(csr_n510), .A2(csr_wdata_13_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[13]), .Y(csr_n_GEN_293[13]) );
  AO22X1_LVT csr_U2620 ( .A1(csr_n510), .A2(csr_wdata_12_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[12]), .Y(csr_n_GEN_293[12]) );
  AO22X1_LVT csr_U2619 ( .A1(csr_n510), .A2(csr_wdata_10_), .A3(csr_n434), 
        .A4(io_ptw_pmp_5_addr[10]), .Y(csr_n_GEN_293[10]) );
  AO22X1_LVT csr_U2618 ( .A1(csr_n510), .A2(csr_wdata_0_), .A3(csr_n434), .A4(
        io_ptw_pmp_5_addr[0]), .Y(csr_n_GEN_293[0]) );
  AO22X1_LVT csr_U2617 ( .A1(csr_n509), .A2(csr_wdata_8_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[8]), .Y(csr_n_GEN_286[8]) );
  AO22X1_LVT csr_U2616 ( .A1(csr_n509), .A2(csr_wdata_6_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[6]), .Y(csr_n_GEN_286[6]) );
  AO22X1_LVT csr_U2615 ( .A1(csr_n509), .A2(csr_wdata_5_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[5]), .Y(csr_n_GEN_286[5]) );
  AO22X1_LVT csr_U2614 ( .A1(csr_n509), .A2(csr_wdata_4_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[4]), .Y(csr_n_GEN_286[4]) );
  AO22X1_LVT csr_U2613 ( .A1(csr_n509), .A2(csr_wdata_2_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[2]), .Y(csr_n_GEN_286[2]) );
  AO22X1_LVT csr_U2612 ( .A1(csr_n509), .A2(csr_wdata_29_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[29]), .Y(csr_n_GEN_286[29]) );
  AO22X1_LVT csr_U2611 ( .A1(csr_n509), .A2(csr_wdata_28_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[28]), .Y(csr_n_GEN_286[28]) );
  AO22X1_LVT csr_U2610 ( .A1(csr_n509), .A2(csr_wdata_27_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[27]), .Y(csr_n_GEN_286[27]) );
  AO22X1_LVT csr_U2609 ( .A1(csr_n509), .A2(csr_wdata_26_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[26]), .Y(csr_n_GEN_286[26]) );
  AO22X1_LVT csr_U2608 ( .A1(csr_n509), .A2(csr_wdata_25_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[25]), .Y(csr_n_GEN_286[25]) );
  AO22X1_LVT csr_U2607 ( .A1(csr_n509), .A2(csr_wdata_24_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[24]), .Y(csr_n_GEN_286[24]) );
  AO22X1_LVT csr_U2606 ( .A1(csr_n509), .A2(csr_wdata_23_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[23]), .Y(csr_n_GEN_286[23]) );
  AO22X1_LVT csr_U2605 ( .A1(csr_n509), .A2(csr_wdata_22_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[22]), .Y(csr_n_GEN_286[22]) );
  AO22X1_LVT csr_U2604 ( .A1(csr_n509), .A2(csr_wdata_21_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[21]), .Y(csr_n_GEN_286[21]) );
  AO22X1_LVT csr_U2603 ( .A1(csr_n509), .A2(csr_wdata_20_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[20]), .Y(csr_n_GEN_286[20]) );
  AO22X1_LVT csr_U2602 ( .A1(csr_n509), .A2(csr_wdata_1_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[1]), .Y(csr_n_GEN_286[1]) );
  AO22X1_LVT csr_U2601 ( .A1(csr_n509), .A2(csr_wdata_19_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[19]), .Y(csr_n_GEN_286[19]) );
  AO22X1_LVT csr_U2600 ( .A1(csr_n509), .A2(csr_wdata_18_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[18]), .Y(csr_n_GEN_286[18]) );
  AO22X1_LVT csr_U2599 ( .A1(csr_n509), .A2(csr_wdata_17_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[17]), .Y(csr_n_GEN_286[17]) );
  AO22X1_LVT csr_U2598 ( .A1(csr_n509), .A2(csr_wdata_16_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[16]), .Y(csr_n_GEN_286[16]) );
  AO22X1_LVT csr_U2597 ( .A1(csr_n509), .A2(csr_wdata_15_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[15]), .Y(csr_n_GEN_286[15]) );
  AO22X1_LVT csr_U2596 ( .A1(csr_n509), .A2(csr_wdata_14_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[14]), .Y(csr_n_GEN_286[14]) );
  AO22X1_LVT csr_U2595 ( .A1(csr_n509), .A2(csr_wdata_13_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[13]), .Y(csr_n_GEN_286[13]) );
  AO22X1_LVT csr_U2594 ( .A1(csr_n509), .A2(csr_wdata_12_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[12]), .Y(csr_n_GEN_286[12]) );
  AO22X1_LVT csr_U2593 ( .A1(csr_n509), .A2(csr_wdata_10_), .A3(csr_n433), 
        .A4(io_ptw_pmp_4_addr[10]), .Y(csr_n_GEN_286[10]) );
  AO22X1_LVT csr_U2592 ( .A1(csr_n509), .A2(csr_wdata_0_), .A3(csr_n433), .A4(
        io_ptw_pmp_4_addr[0]), .Y(csr_n_GEN_286[0]) );
  AO22X1_LVT csr_U2591 ( .A1(csr_n508), .A2(csr_wdata_8_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[8]), .Y(csr_n_GEN_279[8]) );
  AO22X1_LVT csr_U2590 ( .A1(csr_n508), .A2(csr_wdata_6_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[6]), .Y(csr_n_GEN_279[6]) );
  AO22X1_LVT csr_U2589 ( .A1(csr_n508), .A2(csr_wdata_5_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[5]), .Y(csr_n_GEN_279[5]) );
  AO22X1_LVT csr_U2588 ( .A1(csr_n508), .A2(csr_wdata_4_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[4]), .Y(csr_n_GEN_279[4]) );
  AO22X1_LVT csr_U2587 ( .A1(csr_n508), .A2(csr_wdata_2_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[2]), .Y(csr_n_GEN_279[2]) );
  AO22X1_LVT csr_U2586 ( .A1(csr_n508), .A2(csr_wdata_29_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[29]), .Y(csr_n_GEN_279[29]) );
  AO22X1_LVT csr_U2585 ( .A1(csr_n508), .A2(csr_wdata_28_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[28]), .Y(csr_n_GEN_279[28]) );
  AO22X1_LVT csr_U2584 ( .A1(csr_n508), .A2(csr_wdata_27_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[27]), .Y(csr_n_GEN_279[27]) );
  AO22X1_LVT csr_U2583 ( .A1(csr_n508), .A2(csr_wdata_26_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[26]), .Y(csr_n_GEN_279[26]) );
  AO22X1_LVT csr_U2582 ( .A1(csr_n508), .A2(csr_wdata_25_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[25]), .Y(csr_n_GEN_279[25]) );
  AO22X1_LVT csr_U2581 ( .A1(csr_n508), .A2(csr_wdata_24_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[24]), .Y(csr_n_GEN_279[24]) );
  AO22X1_LVT csr_U2580 ( .A1(csr_n508), .A2(csr_wdata_23_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[23]), .Y(csr_n_GEN_279[23]) );
  AO22X1_LVT csr_U2579 ( .A1(csr_n508), .A2(csr_wdata_22_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[22]), .Y(csr_n_GEN_279[22]) );
  AO22X1_LVT csr_U2578 ( .A1(csr_n508), .A2(csr_wdata_21_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[21]), .Y(csr_n_GEN_279[21]) );
  AO22X1_LVT csr_U2577 ( .A1(csr_n508), .A2(csr_wdata_20_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[20]), .Y(csr_n_GEN_279[20]) );
  AO22X1_LVT csr_U2576 ( .A1(csr_n508), .A2(csr_wdata_1_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[1]), .Y(csr_n_GEN_279[1]) );
  AO22X1_LVT csr_U2575 ( .A1(csr_n508), .A2(csr_wdata_19_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[19]), .Y(csr_n_GEN_279[19]) );
  AO22X1_LVT csr_U2574 ( .A1(csr_n508), .A2(csr_wdata_18_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[18]), .Y(csr_n_GEN_279[18]) );
  AO22X1_LVT csr_U2573 ( .A1(csr_n508), .A2(csr_wdata_17_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[17]), .Y(csr_n_GEN_279[17]) );
  AO22X1_LVT csr_U2572 ( .A1(csr_n508), .A2(csr_wdata_16_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[16]), .Y(csr_n_GEN_279[16]) );
  AO22X1_LVT csr_U2571 ( .A1(csr_n508), .A2(csr_wdata_15_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[15]), .Y(csr_n_GEN_279[15]) );
  AO22X1_LVT csr_U2570 ( .A1(csr_n508), .A2(csr_wdata_14_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[14]), .Y(csr_n_GEN_279[14]) );
  AO22X1_LVT csr_U2569 ( .A1(csr_n508), .A2(csr_wdata_13_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[13]), .Y(csr_n_GEN_279[13]) );
  AO22X1_LVT csr_U2568 ( .A1(csr_n508), .A2(csr_wdata_12_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[12]), .Y(csr_n_GEN_279[12]) );
  AO22X1_LVT csr_U2567 ( .A1(csr_n508), .A2(csr_wdata_10_), .A3(csr_n436), 
        .A4(io_ptw_pmp_3_addr[10]), .Y(csr_n_GEN_279[10]) );
  AO22X1_LVT csr_U2566 ( .A1(csr_n508), .A2(csr_wdata_0_), .A3(csr_n436), .A4(
        io_ptw_pmp_3_addr[0]), .Y(csr_n_GEN_279[0]) );
  AO22X1_LVT csr_U2565 ( .A1(csr_n507), .A2(csr_wdata_8_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[8]), .Y(csr_n_GEN_272[8]) );
  AO22X1_LVT csr_U2564 ( .A1(csr_n507), .A2(csr_wdata_6_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[6]), .Y(csr_n_GEN_272[6]) );
  AO22X1_LVT csr_U2563 ( .A1(csr_n507), .A2(csr_wdata_5_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[5]), .Y(csr_n_GEN_272[5]) );
  AO22X1_LVT csr_U2562 ( .A1(csr_n507), .A2(csr_wdata_4_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[4]), .Y(csr_n_GEN_272[4]) );
  AO22X1_LVT csr_U2561 ( .A1(csr_n507), .A2(csr_wdata_2_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[2]), .Y(csr_n_GEN_272[2]) );
  AO22X1_LVT csr_U2560 ( .A1(csr_n507), .A2(csr_wdata_29_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[29]), .Y(csr_n_GEN_272[29]) );
  AO22X1_LVT csr_U2559 ( .A1(csr_n507), .A2(csr_wdata_28_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[28]), .Y(csr_n_GEN_272[28]) );
  AO22X1_LVT csr_U2558 ( .A1(csr_n507), .A2(csr_wdata_27_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[27]), .Y(csr_n_GEN_272[27]) );
  AO22X1_LVT csr_U2557 ( .A1(csr_n507), .A2(csr_wdata_26_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[26]), .Y(csr_n_GEN_272[26]) );
  AO22X1_LVT csr_U2556 ( .A1(csr_n507), .A2(csr_wdata_25_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[25]), .Y(csr_n_GEN_272[25]) );
  AO22X1_LVT csr_U2555 ( .A1(csr_n507), .A2(csr_wdata_24_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[24]), .Y(csr_n_GEN_272[24]) );
  AO22X1_LVT csr_U2554 ( .A1(csr_n507), .A2(csr_wdata_23_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[23]), .Y(csr_n_GEN_272[23]) );
  AO22X1_LVT csr_U2553 ( .A1(csr_n507), .A2(csr_wdata_22_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[22]), .Y(csr_n_GEN_272[22]) );
  AO22X1_LVT csr_U2552 ( .A1(csr_n507), .A2(csr_wdata_21_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[21]), .Y(csr_n_GEN_272[21]) );
  AO22X1_LVT csr_U2551 ( .A1(csr_n507), .A2(csr_wdata_20_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[20]), .Y(csr_n_GEN_272[20]) );
  AO22X1_LVT csr_U2550 ( .A1(csr_n507), .A2(csr_wdata_1_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[1]), .Y(csr_n_GEN_272[1]) );
  AO22X1_LVT csr_U2549 ( .A1(csr_n507), .A2(csr_wdata_19_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[19]), .Y(csr_n_GEN_272[19]) );
  AO22X1_LVT csr_U2548 ( .A1(csr_n507), .A2(csr_wdata_18_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[18]), .Y(csr_n_GEN_272[18]) );
  AO22X1_LVT csr_U2547 ( .A1(csr_n507), .A2(csr_wdata_17_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[17]), .Y(csr_n_GEN_272[17]) );
  AO22X1_LVT csr_U2546 ( .A1(csr_n507), .A2(csr_wdata_16_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[16]), .Y(csr_n_GEN_272[16]) );
  AO22X1_LVT csr_U2545 ( .A1(csr_n507), .A2(csr_wdata_15_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[15]), .Y(csr_n_GEN_272[15]) );
  AO22X1_LVT csr_U2544 ( .A1(csr_n507), .A2(csr_wdata_14_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[14]), .Y(csr_n_GEN_272[14]) );
  AO22X1_LVT csr_U2543 ( .A1(csr_n507), .A2(csr_wdata_13_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[13]), .Y(csr_n_GEN_272[13]) );
  AO22X1_LVT csr_U2542 ( .A1(csr_n507), .A2(csr_wdata_12_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[12]), .Y(csr_n_GEN_272[12]) );
  AO22X1_LVT csr_U2541 ( .A1(csr_n507), .A2(csr_wdata_10_), .A3(csr_n432), 
        .A4(io_ptw_pmp_2_addr[10]), .Y(csr_n_GEN_272[10]) );
  AO22X1_LVT csr_U2540 ( .A1(csr_n507), .A2(csr_wdata_0_), .A3(csr_n432), .A4(
        io_ptw_pmp_2_addr[0]), .Y(csr_n_GEN_272[0]) );
  AO22X1_LVT csr_U2539 ( .A1(csr_n506), .A2(csr_wdata_8_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[8]), .Y(csr_n_GEN_265[8]) );
  AO22X1_LVT csr_U2538 ( .A1(csr_n506), .A2(csr_wdata_6_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[6]), .Y(csr_n_GEN_265[6]) );
  AO22X1_LVT csr_U2537 ( .A1(csr_n506), .A2(csr_wdata_5_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[5]), .Y(csr_n_GEN_265[5]) );
  AO22X1_LVT csr_U2536 ( .A1(csr_n506), .A2(csr_wdata_4_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[4]), .Y(csr_n_GEN_265[4]) );
  AO22X1_LVT csr_U2535 ( .A1(csr_n506), .A2(csr_wdata_2_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[2]), .Y(csr_n_GEN_265[2]) );
  AO22X1_LVT csr_U2534 ( .A1(csr_n506), .A2(csr_wdata_29_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[29]), .Y(csr_n_GEN_265[29]) );
  AO22X1_LVT csr_U2533 ( .A1(csr_n506), .A2(csr_wdata_28_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[28]), .Y(csr_n_GEN_265[28]) );
  AO22X1_LVT csr_U2532 ( .A1(csr_n506), .A2(csr_wdata_27_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[27]), .Y(csr_n_GEN_265[27]) );
  AO22X1_LVT csr_U2531 ( .A1(csr_n506), .A2(csr_wdata_26_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[26]), .Y(csr_n_GEN_265[26]) );
  AO22X1_LVT csr_U2530 ( .A1(csr_n506), .A2(csr_wdata_25_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[25]), .Y(csr_n_GEN_265[25]) );
  AO22X1_LVT csr_U2529 ( .A1(csr_n506), .A2(csr_wdata_24_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[24]), .Y(csr_n_GEN_265[24]) );
  AO22X1_LVT csr_U2528 ( .A1(csr_n506), .A2(csr_wdata_23_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[23]), .Y(csr_n_GEN_265[23]) );
  AO22X1_LVT csr_U2527 ( .A1(csr_n506), .A2(csr_wdata_22_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[22]), .Y(csr_n_GEN_265[22]) );
  AO22X1_LVT csr_U2526 ( .A1(csr_n506), .A2(csr_wdata_21_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[21]), .Y(csr_n_GEN_265[21]) );
  AO22X1_LVT csr_U2525 ( .A1(csr_n506), .A2(csr_wdata_20_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[20]), .Y(csr_n_GEN_265[20]) );
  AO22X1_LVT csr_U2524 ( .A1(csr_n506), .A2(csr_wdata_1_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[1]), .Y(csr_n_GEN_265[1]) );
  AO22X1_LVT csr_U2523 ( .A1(csr_n506), .A2(csr_wdata_19_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[19]), .Y(csr_n_GEN_265[19]) );
  AO22X1_LVT csr_U2522 ( .A1(csr_n506), .A2(csr_wdata_18_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[18]), .Y(csr_n_GEN_265[18]) );
  AO22X1_LVT csr_U2521 ( .A1(csr_n506), .A2(csr_wdata_17_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[17]), .Y(csr_n_GEN_265[17]) );
  AO22X1_LVT csr_U2520 ( .A1(csr_n506), .A2(csr_wdata_16_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[16]), .Y(csr_n_GEN_265[16]) );
  AO22X1_LVT csr_U2519 ( .A1(csr_n506), .A2(csr_wdata_15_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[15]), .Y(csr_n_GEN_265[15]) );
  AO22X1_LVT csr_U2518 ( .A1(csr_n506), .A2(csr_wdata_14_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[14]), .Y(csr_n_GEN_265[14]) );
  AO22X1_LVT csr_U2517 ( .A1(csr_n506), .A2(csr_wdata_13_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[13]), .Y(csr_n_GEN_265[13]) );
  AO22X1_LVT csr_U2516 ( .A1(csr_n506), .A2(csr_wdata_12_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[12]), .Y(csr_n_GEN_265[12]) );
  AO22X1_LVT csr_U2515 ( .A1(csr_n506), .A2(csr_wdata_10_), .A3(csr_n431), 
        .A4(io_ptw_pmp_1_addr[10]), .Y(csr_n_GEN_265[10]) );
  AO22X1_LVT csr_U2514 ( .A1(csr_n506), .A2(csr_wdata_0_), .A3(csr_n431), .A4(
        io_ptw_pmp_1_addr[0]), .Y(csr_n_GEN_265[0]) );
  AO22X1_LVT csr_U2513 ( .A1(csr_n505), .A2(csr_wdata_8_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[8]), .Y(csr_n_GEN_258[8]) );
  AO22X1_LVT csr_U2512 ( .A1(csr_n505), .A2(csr_wdata_6_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[6]), .Y(csr_n_GEN_258[6]) );
  AO22X1_LVT csr_U2511 ( .A1(csr_n505), .A2(csr_wdata_5_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[5]), .Y(csr_n_GEN_258[5]) );
  AO22X1_LVT csr_U2510 ( .A1(csr_n505), .A2(csr_wdata_4_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[4]), .Y(csr_n_GEN_258[4]) );
  AO22X1_LVT csr_U2509 ( .A1(csr_n505), .A2(csr_wdata_2_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[2]), .Y(csr_n_GEN_258[2]) );
  AO22X1_LVT csr_U2508 ( .A1(csr_n505), .A2(csr_wdata_29_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[29]), .Y(csr_n_GEN_258[29]) );
  AO22X1_LVT csr_U2507 ( .A1(csr_n505), .A2(csr_wdata_28_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[28]), .Y(csr_n_GEN_258[28]) );
  AO22X1_LVT csr_U2506 ( .A1(csr_n505), .A2(csr_wdata_27_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[27]), .Y(csr_n_GEN_258[27]) );
  AO22X1_LVT csr_U2505 ( .A1(csr_n505), .A2(csr_wdata_26_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[26]), .Y(csr_n_GEN_258[26]) );
  AO22X1_LVT csr_U2504 ( .A1(csr_n505), .A2(csr_wdata_25_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[25]), .Y(csr_n_GEN_258[25]) );
  AO22X1_LVT csr_U2503 ( .A1(csr_n505), .A2(csr_wdata_24_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[24]), .Y(csr_n_GEN_258[24]) );
  AO22X1_LVT csr_U2502 ( .A1(csr_n505), .A2(csr_wdata_23_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[23]), .Y(csr_n_GEN_258[23]) );
  AO22X1_LVT csr_U2501 ( .A1(csr_n505), .A2(csr_wdata_22_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[22]), .Y(csr_n_GEN_258[22]) );
  AO22X1_LVT csr_U2500 ( .A1(csr_n505), .A2(csr_wdata_21_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[21]), .Y(csr_n_GEN_258[21]) );
  AO22X1_LVT csr_U2499 ( .A1(csr_n505), .A2(csr_wdata_20_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[20]), .Y(csr_n_GEN_258[20]) );
  AO22X1_LVT csr_U2498 ( .A1(csr_n505), .A2(csr_wdata_1_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[1]), .Y(csr_n_GEN_258[1]) );
  AO22X1_LVT csr_U2497 ( .A1(csr_n505), .A2(csr_wdata_19_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[19]), .Y(csr_n_GEN_258[19]) );
  AO22X1_LVT csr_U2496 ( .A1(csr_n505), .A2(csr_wdata_18_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[18]), .Y(csr_n_GEN_258[18]) );
  AO22X1_LVT csr_U2495 ( .A1(csr_n505), .A2(csr_wdata_17_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[17]), .Y(csr_n_GEN_258[17]) );
  AO22X1_LVT csr_U2494 ( .A1(csr_n505), .A2(csr_wdata_16_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[16]), .Y(csr_n_GEN_258[16]) );
  AO22X1_LVT csr_U2493 ( .A1(csr_n505), .A2(csr_wdata_15_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[15]), .Y(csr_n_GEN_258[15]) );
  AO22X1_LVT csr_U2492 ( .A1(csr_n505), .A2(csr_wdata_14_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[14]), .Y(csr_n_GEN_258[14]) );
  AO22X1_LVT csr_U2491 ( .A1(csr_n505), .A2(csr_wdata_13_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[13]), .Y(csr_n_GEN_258[13]) );
  AO22X1_LVT csr_U2490 ( .A1(csr_n505), .A2(csr_wdata_12_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[12]), .Y(csr_n_GEN_258[12]) );
  AO22X1_LVT csr_U2489 ( .A1(csr_n505), .A2(csr_wdata_10_), .A3(csr_n430), 
        .A4(io_ptw_pmp_0_addr[10]), .Y(csr_n_GEN_258[10]) );
  AO22X1_LVT csr_U2488 ( .A1(csr_n505), .A2(csr_wdata_0_), .A3(csr_n430), .A4(
        io_ptw_pmp_0_addr[0]), .Y(csr_n_GEN_258[0]) );
  AO22X1_LVT csr_U2487 ( .A1(csr_n1477), .A2(csr_wdata_6_), .A3(csr_n1696), 
        .A4(csr_wdata_1_), .Y(csr_n_GEN_155[1]) );
  AO22X1_LVT csr_U2486 ( .A1(csr_n1477), .A2(csr_wdata_5_), .A3(csr_n1696), 
        .A4(csr_wdata_0_), .Y(csr_n_GEN_155[0]) );
  AND2X1_LVT csr_U2485 ( .A1(csr_n1504), .A2(csr_n504), .Y(csr_N670) );
  OA21X1_LVT csr_U2484 ( .A1(csr_io_rw_addr[9]), .A2(csr_read_mideleg_5), .A3(
        csr_wdata_5_), .Y(csr_n1695) );
  OA21X1_LVT csr_U2483 ( .A1(csr_io_rw_addr[9]), .A2(csr_read_mideleg_1), .A3(
        csr_wdata_1_), .Y(csr_n1693) );
  AND2X1_LVT csr_U2482 ( .A1(csr_n1510), .A2(csr_n504), .Y(csr_N475) );
  AND2X1_LVT csr_U2481 ( .A1(csr_n504), .A2(csr_n1469), .Y(csr_N460) );
  AND2X1_LVT csr_U2480 ( .A1(csr_n504), .A2(csr_n1691), .Y(csr_N459) );
  AOI22X1_LVT csr_U2479 ( .A1(csr_n1485), .A2(csr_reg_mscratch[58]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[58]), .Y(csr_n1688) );
  AOI22X1_LVT csr_U2478 ( .A1(csr_n1485), .A2(csr_reg_mscratch[57]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[57]), .Y(csr_n1687) );
  AOI22X1_LVT csr_U2477 ( .A1(csr_n1507), .A2(io_ptw_pmp_7_cfg_r), .A3(
        csr_n1508), .A4(csr_reg_sscratch[56]), .Y(csr_n1686) );
  AOI22X1_LVT csr_U2476 ( .A1(csr_n1510), .A2(csr_reg_dscratch[52]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[52]), .Y(csr_n1685) );
  AOI22X1_LVT csr_U2475 ( .A1(csr_n1510), .A2(csr_reg_dscratch[51]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[51]), .Y(csr_n1684) );
  AOI22X1_LVT csr_U2474 ( .A1(csr_n1485), .A2(csr_reg_mscratch[50]), .A3(
        csr_n1507), .A4(io_ptw_pmp_6_cfg_x), .Y(csr_n1683) );
  AOI22X1_LVT csr_U2473 ( .A1(csr_n1510), .A2(csr_reg_dscratch[49]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[49]), .Y(csr_n1682) );
  AOI22X1_LVT csr_U2472 ( .A1(csr_n1510), .A2(csr_reg_dscratch[48]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[48]), .Y(csr_n1681) );
  AOI22X1_LVT csr_U2471 ( .A1(csr_n1510), .A2(csr_reg_dscratch[47]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[47]), .Y(csr_n1680) );
  AOI22X1_LVT csr_U2470 ( .A1(csr_n1510), .A2(csr_reg_dscratch[43]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[43]), .Y(csr_n1678) );
  AOI22X1_LVT csr_U2469 ( .A1(csr_n1510), .A2(csr_reg_dscratch[42]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[42]), .Y(csr_n1677) );
  AOI22X1_LVT csr_U2468 ( .A1(csr_n1510), .A2(csr_reg_dscratch[41]), .A3(
        csr_n1507), .A4(io_ptw_pmp_5_cfg_w), .Y(csr_n1676) );
  AOI22X1_LVT csr_U2467 ( .A1(csr_n1507), .A2(io_ptw_pmp_5_cfg_r), .A3(
        csr_n1508), .A4(csr_reg_sscratch[40]), .Y(csr_n1675) );
  NAND2X0_LVT csr_U2466 ( .A1(csr_n488), .A2(csr_n504), .Y(csr_n1673) );
  AND2X1_LVT csr_U2465 ( .A1(csr_n1508), .A2(csr_n504), .Y(csr_N1422) );
  AO22X1_LVT csr_U2464 ( .A1(csr_n1485), .A2(csr_reg_mscratch[63]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[63]), .Y(csr_n1672) );
  OR3X1_LVT csr_U2463 ( .A1(csr_n1666), .A2(csr_n1665), .A3(csr_n1664), .Y(
        csr_n1667) );
  OR3X1_LVT csr_U2462 ( .A1(csr_n1663), .A2(csr_n1662), .A3(csr_n1661), .Y(
        csr_n1664) );
  AO22X1_LVT csr_U2461 ( .A1(csr_n1507), .A2(io_ptw_pmp_0_cfg_x), .A3(
        csr_read_medeleg_2_), .A4(csr_n1469), .Y(csr_n1661) );
  AO22X1_LVT csr_U2460 ( .A1(csr_n488), .A2(io_ptw_ptbr_ppn[2]), .A3(csr_n1472), .A4(io_ptw_pmp_5_addr[2]), .Y(csr_n1662) );
  AO22X1_LVT csr_U2459 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[2]), .A3(
        csr_n1489), .A4(csr_reg_mepc_2_), .Y(csr_n1665) );
  AO22X1_LVT csr_U2458 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[2]), .A3(
        csr_reg_mtvec_2_), .A4(csr_n1470), .Y(csr_n1668) );
  AO22X1_LVT csr_U2457 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[2]), .A3(
        csr_n1506), .A4(csr_reg_sepc_2_), .Y(csr_n1660) );
  AO22X1_LVT csr_U2456 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[2]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[2]), .Y(csr_n1658) );
  AO22X1_LVT csr_U2455 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[2]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[2]), .Y(csr_n1659) );
  AO22X1_LVT csr_U2454 ( .A1(csr_n1487), .A2(csr_n428), .A3(csr_n1492), .A4(
        io_ptw_pmp_2_addr[0]), .Y(csr_n1655) );
  AO22X1_LVT csr_U2453 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[0]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[0]), .Y(csr_n1657) );
  AO22X1_LVT csr_U2452 ( .A1(csr_n1485), .A2(csr_reg_mscratch[0]), .A3(
        csr_read_medeleg_0), .A4(csr_n1469), .Y(csr_n1654) );
  AO22X1_LVT csr_U2451 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[0]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[0]), .Y(csr_n1651) );
  AO22X1_LVT csr_U2450 ( .A1(csr_n1508), .A2(csr_reg_sscratch[0]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[0]), .Y(csr_n1652) );
  AO22X1_LVT csr_U2449 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[0]), .A3(
        csr_n1484), .A4(csr_read_mcounteren_0_), .Y(csr_n1653) );
  AND2X1_LVT csr_U2448 ( .A1(csr_n1485), .A2(csr_n504), .Y(csr_N1033) );
  AO22X1_LVT csr_U2447 ( .A1(csr_n1489), .A2(csr_reg_mepc_39_), .A3(csr_n1506), 
        .A4(csr_reg_sepc_39_), .Y(csr_n1649) );
  AO22X1_LVT csr_U2446 ( .A1(csr_n1487), .A2(csr_reg_stvec_38_), .A3(csr_n1490), .A4(csr_io_bp_0_address[38]), .Y(csr_n1650) );
  OR4X1_LVT csr_U2445 ( .A1(csr_n1647), .A2(csr_n1646), .A3(csr_n1645), .A4(
        csr_n1644), .Y(csr_n1648) );
  AO22X1_LVT csr_U2444 ( .A1(csr_n1493), .A2(csr_reg_dpc_37_), .A3(csr_n1506), 
        .A4(csr_reg_sepc_37_), .Y(csr_n1646) );
  AO22X1_LVT csr_U2443 ( .A1(csr_n1510), .A2(csr_reg_dscratch[37]), .A3(
        csr_n1489), .A4(csr_reg_mepc_37_), .Y(csr_n1647) );
  OR4X1_LVT csr_U2442 ( .A1(csr_n1642), .A2(csr_n1641), .A3(csr_n1640), .A4(
        csr_n1639), .Y(csr_n1643) );
  AO22X1_LVT csr_U2441 ( .A1(csr_n1493), .A2(csr_reg_dpc_36_), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[36]), .Y(csr_n1639) );
  AO22X1_LVT csr_U2440 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[36]), .A3(
        csr_n1510), .A4(csr_reg_dscratch[36]), .Y(csr_n1641) );
  AO22X1_LVT csr_U2439 ( .A1(csr_n1489), .A2(csr_reg_mepc_36_), .A3(csr_n1485), 
        .A4(csr_reg_mscratch[36]), .Y(csr_n1642) );
  OR4X1_LVT csr_U2438 ( .A1(csr_n1637), .A2(csr_n1636), .A3(csr_n1635), .A4(
        csr_n1634), .Y(csr_n1638) );
  AO22X1_LVT csr_U2437 ( .A1(csr_n1485), .A2(csr_reg_mscratch[34]), .A3(
        csr_n1507), .A4(io_ptw_pmp_4_cfg_x), .Y(csr_n1637) );
  OR4X1_LVT csr_U2436 ( .A1(csr_n1632), .A2(csr_n1631), .A3(csr_n1630), .A4(
        csr_n1629), .Y(csr_n1633) );
  AO22X1_LVT csr_U2435 ( .A1(csr_n1507), .A2(io_ptw_pmp_4_cfg_r), .A3(
        csr_n1508), .A4(csr_reg_sscratch[32]), .Y(csr_n1632) );
  AO22X1_LVT csr_U2434 ( .A1(csr_n1508), .A2(csr_reg_sscratch[30]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_30_), .Y(csr_n1628) );
  AO22X1_LVT csr_U2433 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[29]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[29]), .Y(csr_n1625) );
  AO21X1_LVT csr_U2432 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[29]), .A3(
        csr_n1670), .Y(csr_n1626) );
  AO22X1_LVT csr_U2431 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[29]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_29_), .Y(csr_n1623) );
  AO22X1_LVT csr_U2430 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[29]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[29]), .Y(csr_n1624) );
  AO22X1_LVT csr_U2429 ( .A1(csr_n1485), .A2(csr_reg_mscratch[29]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[29]), .Y(csr_n1620) );
  AO22X1_LVT csr_U2428 ( .A1(csr_n1510), .A2(csr_reg_dscratch[29]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[29]), .Y(csr_n1621) );
  AO22X1_LVT csr_U2427 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[29]), .A3(
        csr_n1506), .A4(csr_reg_sepc_29_), .Y(csr_n1622) );
  AO22X1_LVT csr_U2426 ( .A1(csr_n1487), .A2(csr_reg_stvec_27_), .A3(csr_n1497), .A4(csr_reg_mtvec_27_), .Y(csr_n1617) );
  AO22X1_LVT csr_U2425 ( .A1(csr_n1510), .A2(csr_reg_dscratch[27]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[27]), .Y(csr_n1618) );
  AO22X1_LVT csr_U2424 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[27]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[27]), .Y(csr_n1619) );
  AO22X1_LVT csr_U2423 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[27]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[27]), .Y(csr_n1615) );
  AO22X1_LVT csr_U2422 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[27]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[27]), .Y(csr_n1616) );
  AO22X1_LVT csr_U2421 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[27]), .A3(
        csr_n1489), .A4(csr_reg_mepc_27_), .Y(csr_n1614) );
  AO22X1_LVT csr_U2420 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[24]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[24]), .Y(csr_n1612) );
  AO22X1_LVT csr_U2419 ( .A1(csr_n1489), .A2(csr_reg_mepc_24_), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[24]), .Y(csr_n1608) );
  AO22X1_LVT csr_U2418 ( .A1(csr_n1510), .A2(csr_reg_dscratch[24]), .A3(
        csr_n1506), .A4(csr_reg_sepc_24_), .Y(csr_n1609) );
  AO22X1_LVT csr_U2417 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[24]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[24]), .Y(csr_n1610) );
  AO22X1_LVT csr_U2416 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[24]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[24]), .Y(csr_n1611) );
  AO22X1_LVT csr_U2415 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[24]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[24]), .Y(csr_n1606) );
  AO22X1_LVT csr_U2414 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[24]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[24]), .Y(csr_n1607) );
  AO21X1_LVT csr_U2413 ( .A1(csr_n1487), .A2(csr_reg_stvec_23_), .A3(csr_n1603), .Y(csr_n1604) );
  AO22X1_LVT csr_U2412 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[23]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[23]), .Y(csr_n1602) );
  AO22X1_LVT csr_U2411 ( .A1(csr_n1485), .A2(csr_reg_mscratch[23]), .A3(
        csr_n1493), .A4(csr_reg_dpc_23_), .Y(csr_n1598) );
  AO22X1_LVT csr_U2410 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[23]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[23]), .Y(csr_n1599) );
  AO22X1_LVT csr_U2409 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[23]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[23]), .Y(csr_n1600) );
  AO22X1_LVT csr_U2408 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[23]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_23_), .Y(csr_n1601) );
  AO21X1_LVT csr_U2407 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[20]), .A3(
        csr_n1596), .Y(csr_n1597) );
  AO22X1_LVT csr_U2406 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[20]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[20]), .Y(csr_n1595) );
  AO22X1_LVT csr_U2405 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[20]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[20]), .Y(csr_n1592) );
  AO22X1_LVT csr_U2404 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[20]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_20_), .Y(csr_n1593) );
  AO22X1_LVT csr_U2403 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[20]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[20]), .Y(csr_n1594) );
  AO22X1_LVT csr_U2402 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[19]), .A3(
        csr_n1506), .A4(csr_reg_sepc_19_), .Y(csr_n1588) );
  AO22X1_LVT csr_U2401 ( .A1(csr_n1489), .A2(csr_reg_mepc_19_), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[19]), .Y(csr_n1589) );
  AO22X1_LVT csr_U2400 ( .A1(csr_n1510), .A2(csr_reg_dscratch[19]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[19]), .Y(csr_n1590) );
  AO22X1_LVT csr_U2399 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[19]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[19]), .Y(csr_n1587) );
  AO22X1_LVT csr_U2398 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[18]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[18]), .Y(csr_n1585) );
  AO22X1_LVT csr_U2397 ( .A1(csr_n1485), .A2(csr_reg_mscratch[18]), .A3(
        csr_n1493), .A4(csr_reg_dpc_18_), .Y(csr_n1586) );
  AO22X1_LVT csr_U2396 ( .A1(csr_n1489), .A2(csr_reg_mepc_18_), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[18]), .Y(csr_n1583) );
  AO22X1_LVT csr_U2395 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[18]), .A3(
        csr_n1506), .A4(csr_reg_sepc_18_), .Y(csr_n1584) );
  AO22X1_LVT csr_U2394 ( .A1(csr_n1488), .A2(io_ptw_ptbr_ppn[18]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[18]), .Y(csr_n1582) );
  NAND2X0_LVT csr_U2393 ( .A1(csr_n1487), .A2(csr_reg_stvec_17_), .Y(csr_n1579) );
  AO22X1_LVT csr_U2392 ( .A1(csr_n1510), .A2(csr_reg_dscratch[17]), .A3(
        csr_n1506), .A4(csr_reg_sepc_17_), .Y(csr_n1575) );
  AO22X1_LVT csr_U2391 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[17]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[17]), .Y(csr_n1576) );
  AO22X1_LVT csr_U2390 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[17]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[17]), .Y(csr_n1571) );
  AO22X1_LVT csr_U2389 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[17]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_17_), .Y(csr_n1572) );
  AO22X1_LVT csr_U2388 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[17]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[17]), .Y(csr_n1574) );
  AO21X1_LVT csr_U2387 ( .A1(csr_n1487), .A2(csr_reg_stvec_16_), .A3(csr_n1568), .Y(csr_n1569) );
  AO22X1_LVT csr_U2386 ( .A1(csr_n488), .A2(io_ptw_ptbr_ppn[16]), .A3(
        csr_n1506), .A4(csr_reg_sepc_16_), .Y(csr_n1568) );
  AO22X1_LVT csr_U2385 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[16]), .A3(
        csr_n1489), .A4(csr_reg_mepc_16_), .Y(csr_n1564) );
  AO22X1_LVT csr_U2384 ( .A1(csr_n1485), .A2(csr_reg_mscratch[16]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[16]), .Y(csr_n1565) );
  AO22X1_LVT csr_U2383 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[16]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[16]), .Y(csr_n1566) );
  AO22X1_LVT csr_U2382 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[16]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[16]), .Y(csr_n1567) );
  AO22X1_LVT csr_U2381 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[16]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_16_), .Y(csr_n1561) );
  AO22X1_LVT csr_U2380 ( .A1(csr_n1507), .A2(io_ptw_pmp_2_cfg_r), .A3(
        csr_n1508), .A4(csr_reg_sscratch[16]), .Y(csr_n1562) );
  AO22X1_LVT csr_U2379 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[16]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[16]), .Y(csr_n1563) );
  AO22X1_LVT csr_U2378 ( .A1(csr_n1506), .A2(csr_reg_sepc_15_), .A3(
        csr_read_medeleg_15), .A4(csr_n1469), .Y(csr_n1560) );
  AO22X1_LVT csr_U2377 ( .A1(csr_n1493), .A2(csr_reg_dpc_13_), .A3(csr_n1506), 
        .A4(csr_reg_sepc_13_), .Y(csr_n1559) );
  AND2X1_LVT csr_U2376 ( .A1(csr_io_rw_addr[0]), .A2(csr_n1656), .Y(csr_n1670)
         );
  AND4X1_LVT csr_U2375 ( .A1(csr_io_rw_addr[1]), .A2(csr_n1558), .A3(csr_n1557), .A4(csr_n1556), .Y(csr_n1656) );
  AND2X1_LVT csr_U2374 ( .A1(csr_io_rw_addr[10]), .A2(csr_io_rw_addr[11]), .Y(
        csr_n1556) );
  AO22X1_LVT csr_U2372 ( .A1(csr_n1502), .A2(csr_reg_mie_1_), .A3(csr_n1465), 
        .A4(csr_read_scounteren_1_), .Y(csr_n1554) );
  NAND3X0_LVT csr_U2371 ( .A1(csr_n1505), .A2(csr_n1509), .A3(csr_n_T_61_1), 
        .Y(csr_n1552) );
  NAND3X0_LVT csr_U2370 ( .A1(csr_n1504), .A2(csr_reg_mie_1_), .A3(csr_n1515), 
        .Y(csr_n1692) );
  AO22X1_LVT csr_U2369 ( .A1(csr_n1510), .A2(csr_reg_dscratch[1]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[1]), .Y(csr_n1548) );
  AO22X1_LVT csr_U2368 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[1]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[1]), .Y(csr_n1549) );
  AO22X1_LVT csr_U2367 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[1]), .A3(
        csr_n1466), .A4(io_fpu_fcsr_rm[1]), .Y(csr_n1550) );
  AND2X1_LVT csr_U2366 ( .A1(csr_n1474), .A2(csr_n_T_61_1), .Y(csr_n1551) );
  AO22X1_LVT csr_U2365 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[1]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[1]), .Y(csr_n1547) );
  AO22X1_LVT csr_U2364 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[1]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[1]), .Y(csr_n1545) );
  AO22X1_LVT csr_U2363 ( .A1(csr_n1488), .A2(io_ptw_ptbr_ppn[1]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[1]), .Y(csr_n1546) );
  OR3X1_LVT csr_U2362 ( .A1(csr_n1542), .A2(csr_n1541), .A3(csr_n1540), .Y(
        csr_n1543) );
  AO22X1_LVT csr_U2361 ( .A1(csr_n1474), .A2(csr_n_T_61_5_), .A3(csr_n1493), 
        .A4(csr_reg_dpc_5_), .Y(csr_n1542) );
  NAND3X0_LVT csr_U2360 ( .A1(csr_n1553), .A2(csr_n1694), .A3(csr_n1538), .Y(
        csr_n1539) );
  NAND3X0_LVT csr_U2359 ( .A1(csr_n1505), .A2(csr_n1509), .A3(csr_n_T_61_5_), 
        .Y(csr_n1538) );
  NAND2X0_LVT csr_U2358 ( .A1(csr_n1503), .A2(csr_reg_mie_5_), .Y(csr_n1694)
         );
  AO22X1_LVT csr_U2357 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[5]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[5]), .Y(csr_n1534) );
  AO22X1_LVT csr_U2356 ( .A1(csr_n488), .A2(io_ptw_ptbr_ppn[5]), .A3(csr_n1473), .A4(io_ptw_pmp_3_addr[5]), .Y(csr_n1535) );
  AO22X1_LVT csr_U2355 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[5]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[5]), .Y(csr_n1536) );
  AO22X1_LVT csr_U2354 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[5]), .A3(
        csr_n1506), .A4(csr_reg_sepc_5_), .Y(csr_n1537) );
  AO22X1_LVT csr_U2353 ( .A1(csr_n1493), .A2(csr_reg_dpc_8_), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_8_), .Y(csr_n1533) );
  NAND2X0_LVT csr_U2352 ( .A1(csr_n1674), .A2(csr_n1530), .Y(csr_n1531) );
  NAND3X0_LVT csr_U2351 ( .A1(csr_io_rw_addr[10]), .A2(csr_io_rw_addr[11]), 
        .A3(csr_n1511), .Y(csr_n1530) );
  AND3X1_LVT csr_U2350 ( .A1(csr_n1517), .A2(csr_n1528), .A3(csr_n1518), .Y(
        csr_n1557) );
  NAND3X0_LVT csr_U2348 ( .A1(csr_io_rw_addr[7]), .A2(csr_io_rw_addr[5]), .A3(
        csr_n1513), .Y(csr_n1524) );
  AND4X1_LVT csr_U2347 ( .A1(csr_io_rw_addr[7]), .A2(csr_io_rw_addr[5]), .A3(
        csr_n1558), .A4(csr_n1513), .Y(csr_n1523) );
  NOR3X0_LVT csr_U2346 ( .A1(csr_n1521), .A2(csr_n1525), .A3(csr_io_rw_addr[3]), .Y(csr_n1558) );
  NAND3X0_LVT csr_U2345 ( .A1(csr_io_rw_addr[9]), .A2(csr_io_rw_addr[8]), .A3(
        csr_n1516), .Y(csr_n1525) );
  AND3X1_LVT csr_U2344 ( .A1(csr_io_rw_addr[8]), .A2(csr_n1529), .A3(csr_n1517), .Y(csr_n1522) );
  AND2X1_LVT csr_U2343 ( .A1(csr_n1490), .A2(csr_n1464), .Y(csr_n2163) );
  OR2X1_LVT csr_U2342 ( .A1(csr_n376), .A2(csr_N604), .Y(csr_N595) );
  AND2X1_LVT csr_U2341 ( .A1(csr_n1463), .A2(csr_n442), .Y(csr_N604) );
  OR2X1_LVT csr_U2340 ( .A1(csr_n376), .A2(csr_N542), .Y(csr_N539) );
  AND2X1_LVT csr_U2339 ( .A1(csr_n1463), .A2(csr_n441), .Y(csr_N542) );
  NAND2X0_LVT csr_U2338 ( .A1(csr_n448), .A2(csr_n1462), .Y(csr_net34759) );
  NAND3X0_LVT csr_U2337 ( .A1(csr_n1461), .A2(csr_n590), .A3(csr_n1460), .Y(
        csr_N880) );
  AO21X1_LVT csr_U2336 ( .A1(csr_n1459), .A2(csr_n_T_45_5_), .A3(csr_n1458), 
        .Y(csr_N1496) );
  NAND2X0_LVT csr_U2335 ( .A1(csr_n1457), .A2(csr_n1461), .Y(csr_N992) );
  OR2X1_LVT csr_U2334 ( .A1(csr_n376), .A2(csr_N518), .Y(csr_N515) );
  AND2X1_LVT csr_U2333 ( .A1(csr_n1463), .A2(csr_n453), .Y(csr_N518) );
  OR2X1_LVT csr_U2332 ( .A1(csr_n376), .A2(csr_N568), .Y(csr_N559) );
  NAND2X0_LVT csr_U2331 ( .A1(csr_n1456), .A2(csr_n1462), .Y(csr_N1381) );
  NAND2X0_LVT csr_U2330 ( .A1(csr_n1455), .A2(csr_n1462), .Y(csr_N1269) );
  AO21X1_LVT csr_U2329 ( .A1(csr_n1497), .A2(csr_n504), .A3(csr_n376), .Y(
        csr_n2165) );
  NAND2X0_LVT csr_U2328 ( .A1(csr_n449), .A2(csr_n1461), .Y(csr_net34961) );
  OR2X1_LVT csr_U2327 ( .A1(csr_n376), .A2(csr_N592), .Y(csr_N587) );
  AND2X1_LVT csr_U2326 ( .A1(csr_n1463), .A2(csr_n439), .Y(csr_N592) );
  OR2X1_LVT csr_U2325 ( .A1(csr_n376), .A2(csr_N580), .Y(csr_N575) );
  AND2X1_LVT csr_U2324 ( .A1(csr_n1463), .A2(csr_n437), .Y(csr_N580) );
  AND2X1_LVT csr_U2323 ( .A1(csr_n1463), .A2(csr_n438), .Y(csr_N568) );
  OR2X1_LVT csr_U2322 ( .A1(csr_n376), .A2(csr_N556), .Y(csr_N551) );
  AND2X1_LVT csr_U2321 ( .A1(csr_n1463), .A2(csr_n443), .Y(csr_N556) );
  OR2X1_LVT csr_U2320 ( .A1(csr_n376), .A2(csr_N531), .Y(csr_N527) );
  AND2X1_LVT csr_U2319 ( .A1(csr_n1463), .A2(csr_n440), .Y(csr_N531) );
  NAND2X0_LVT csr_U2318 ( .A1(csr_n590), .A2(csr_n1454), .Y(csr_N1558) );
  NAND3X0_LVT csr_U2317 ( .A1(csr_n1453), .A2(csr_n504), .A3(csr_n1452), .Y(
        csr_n1454) );
  NAND2X0_LVT csr_U2316 ( .A1(csr_io_pc[1]), .A2(csr_n1483), .Y(csr_n1453) );
  NAND2X0_LVT csr_U2315 ( .A1(csr_n1451), .A2(csr_n1461), .Y(csr_N335) );
  OR2X1_LVT csr_U2314 ( .A1(csr_n376), .A2(csr_n1450), .Y(csr_N276) );
  NAND2X0_LVT csr_U2313 ( .A1(csr_n590), .A2(csr_n1449), .Y(csr_N438) );
  NAND2X0_LVT csr_U2312 ( .A1(csr_n450), .A2(csr_n1448), .Y(csr_net35183) );
  OR2X1_LVT csr_U2311 ( .A1(csr_n376), .A2(csr_N487), .Y(csr_N479) );
  AND2X1_LVT csr_U2310 ( .A1(csr_n1481), .A2(csr_n1464), .Y(csr_N487) );
  OA21X1_LVT csr_U2309 ( .A1(csr_io_status_debug), .A2(csr_n457), .A3(csr_n504), .Y(csr_n1464) );
  NAND2X0_LVT csr_U2308 ( .A1(csr_n1447), .A2(csr_n1446), .Y(csr_N1890) );
  MUX21X1_LVT csr_U2307 ( .A1(csr_n_1930_), .A2(io_ptw_status_prv[0]), .S0(
        csr_n1444), .Y(csr_N1691) );
  MUX21X1_LVT csr_U2306 ( .A1(csr_n_1929_), .A2(io_ptw_status_prv[1]), .S0(
        csr_n1444), .Y(csr_N1692) );
  NAND2X0_LVT csr_U2305 ( .A1(csr_n1927), .A2(n9516), .Y(csr_n1444) );
  NAND4X0_LVT csr_U2304 ( .A1(csr_n1440), .A2(csr_n1439), .A3(csr_n1438), .A4(
        csr_n1437), .Y(csr_io_decode_0_read_illegal) );
  NAND3X0_LVT csr_U2303 ( .A1(csr_n1436), .A2(csr_n1435), .A3(csr_n1434), .Y(
        csr_n1437) );
  NAND2X0_LVT csr_U2302 ( .A1(csr_n1433), .A2(ibuf_io_inst_0_bits_raw[24]), 
        .Y(csr_n1434) );
  NAND3X0_LVT csr_U2301 ( .A1(csr_n1431), .A2(csr_n1430), .A3(csr_n1429), .Y(
        csr_n1435) );
  NAND3X0_LVT csr_U2300 ( .A1(csr_n1428), .A2(ibuf_io_inst_0_bits_raw[22]), 
        .A3(csr_n1427), .Y(csr_n1429) );
  AO21X1_LVT csr_U2299 ( .A1(csr_n1426), .A2(csr_n1425), .A3(csr_n1424), .Y(
        csr_n1428) );
  NAND3X0_LVT csr_U2298 ( .A1(csr_n1423), .A2(csr_n1422), .A3(
        csr_io_decode_0_write_flush), .Y(csr_n1431) );
  AND4X1_LVT csr_U2297 ( .A1(csr_n1421), .A2(ibuf_io_inst_0_bits_raw[20]), 
        .A3(csr_n1425), .A4(ibuf_io_inst_0_bits_raw[21]), .Y(csr_n1422) );
  NAND2X0_LVT csr_U2296 ( .A1(csr_n1420), .A2(ibuf_io_inst_0_bits_raw[24]), 
        .Y(csr_n1425) );
  NAND3X0_LVT csr_U2295 ( .A1(csr_n1418), .A2(ibuf_io_inst_0_bits_inst_rs3_2_), 
        .A3(csr_n1417), .Y(csr_n1423) );
  NAND4X0_LVT csr_U2294 ( .A1(csr_n1415), .A2(csr_n1414), .A3(csr_n1413), .A4(
        csr_n1412), .Y(csr_n1438) );
  OA21X1_LVT csr_U2293 ( .A1(csr_n1409), .A2(csr_n1408), .A3(csr_n1407), .Y(
        csr_n1410) );
  NAND4X0_LVT csr_U2292 ( .A1(csr_n1406), .A2(ibuf_io_inst_0_bits_raw[28]), 
        .A3(ibuf_io_inst_0_bits_inst_rs3_2_), .A4(csr_n490), .Y(csr_n1408) );
  NAND3X0_LVT csr_U2291 ( .A1(csr_n1405), .A2(ibuf_io_inst_0_bits_raw[27]), 
        .A3(ibuf_io_inst_0_bits_raw[26]), .Y(csr_n1409) );
  AND3X1_LVT csr_U2290 ( .A1(csr_n1404), .A2(ibuf_io_inst_0_bits_raw[21]), 
        .A3(csr_n1432), .Y(csr_n1411) );
  OA21X1_LVT csr_U2289 ( .A1(io_ptw_status_prv[1]), .A2(csr_n1403), .A3(
        csr_n1402), .Y(csr_n1439) );
  AND3X1_LVT csr_U2288 ( .A1(csr_n1401), .A2(csr_n1400), .A3(csr_n1399), .Y(
        csr_n1402) );
  NAND2X0_LVT csr_U2287 ( .A1(csr_io_decode_0_fp_csr), .A2(
        csr_io_decode_0_fp_illegal), .Y(csr_n1399) );
  NAND4X0_LVT csr_U2286 ( .A1(csr_n1405), .A2(csr_n490), .A3(
        ibuf_io_inst_0_bits_raw[24]), .A4(n9516), .Y(csr_n1400) );
  OA22X1_LVT csr_U2285 ( .A1(csr_n1398), .A2(csr_n1397), .A3(csr_n447), .A4(
        csr_n1396), .Y(csr_n1403) );
  AND3X1_LVT csr_U2284 ( .A1(csr_n1395), .A2(csr_n1412), .A3(csr_n1394), .Y(
        csr_n1397) );
  OAI22X1_LVT csr_U2283 ( .A1(ibuf_io_inst_0_bits_raw[20]), .A2(csr_n1393), 
        .A3(csr_n470), .A4(csr_n1424), .Y(csr_n1394) );
  NAND2X0_LVT csr_U2282 ( .A1(ibuf_io_inst_0_bits_raw[21]), .A2(
        csr_read_mcounteren_2_), .Y(csr_n1393) );
  NOR2X0_LVT csr_U2281 ( .A1(ibuf_io_inst_0_bits_raw[22]), .A2(csr_n1392), .Y(
        csr_n1412) );
  NAND2X0_LVT csr_U2280 ( .A1(csr_n1391), .A2(csr_n429), .Y(csr_n1395) );
  OAI22X1_LVT csr_U2279 ( .A1(csr_read_scounteren_2_), .A2(csr_n1407), .A3(
        csr_read_scounteren_0_), .A4(csr_n1424), .Y(csr_n1391) );
  INVX1_LVT csr_U2278 ( .A(csr_n1390), .Y(csr_n1424) );
  AO21X1_LVT csr_U2277 ( .A1(csr_n1389), .A2(csr_n1416), .A3(csr_n1388), .Y(
        csr_n1440) );
  NAND4X0_LVT csr_U2276 ( .A1(csr_n1387), .A2(csr_n1414), .A3(csr_n1417), .A4(
        csr_n1432), .Y(csr_n1388) );
  OR3X1_LVT csr_U2275 ( .A1(csr_n490), .A2(csr_n1386), .A3(csr_n1385), .Y(
        csr_n1432) );
  OA21X1_LVT csr_U2274 ( .A1(csr_n1383), .A2(csr_n1427), .A3(csr_n1426), .Y(
        csr_n1414) );
  AO22X1_LVT csr_U2273 ( .A1(csr_n1427), .A2(csr_n1390), .A3(csr_n1413), .A4(
        csr_n1382), .Y(csr_n1387) );
  AND2X1_LVT csr_U2272 ( .A1(csr_n1419), .A2(ibuf_io_inst_0_bits_raw[24]), .Y(
        csr_n1382) );
  AND2X1_LVT csr_U2271 ( .A1(csr_n1421), .A2(csr_n1381), .Y(csr_n1413) );
  NAND4X0_LVT csr_U2270 ( .A1(csr_n1380), .A2(csr_n1379), .A3(
        csr_io_decode_0_fp_csr), .A4(csr_n1386), .Y(csr_n1421) );
  NOR2X0_LVT csr_U2269 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(n2576), .Y(
        csr_io_decode_0_fp_csr) );
  NAND3X0_LVT csr_U2268 ( .A1(csr_n1377), .A2(csr_n1376), .A3(csr_n1386), .Y(
        csr_n1427) );
  OR2X1_LVT csr_U2267 ( .A1(csr_n1392), .A2(csr_n1373), .Y(csr_n1389) );
  AND3X1_LVT csr_U2266 ( .A1(csr_n1372), .A2(csr_n1404), .A3(csr_n1396), .Y(
        csr_n1374) );
  NAND4X0_LVT csr_U2265 ( .A1(csr_n1379), .A2(csr_io_decode_0_write_illegal), 
        .A3(csr_n1371), .A4(csr_n1406), .Y(csr_n1398) );
  NAND3X0_LVT csr_U2264 ( .A1(csr_n1406), .A2(n2576), .A3(csr_n1386), .Y(
        csr_n1370) );
  NAND4X0_LVT csr_U2263 ( .A1(csr_n1367), .A2(csr_n1407), .A3(csr_n1430), .A4(
        csr_n1417), .Y(csr_n1372) );
  NAND3X0_LVT csr_U2262 ( .A1(csr_n1384), .A2(ibuf_io_inst_0_bits_raw[27]), 
        .A3(csr_n490), .Y(csr_n1381) );
  AND3X1_LVT csr_U2261 ( .A1(csr_n1376), .A2(ibuf_io_inst_0_bits_inst_rs3_2_), 
        .A3(ibuf_io_inst_0_bits_raw[28]), .Y(csr_n1368) );
  NAND2X0_LVT csr_U2260 ( .A1(csr_n1923), .A2(csr_n1928), .Y(
        csr_io_decode_0_fp_illegal) );
  AND2X1_LVT csr_U2259 ( .A1(csr_n490), .A2(n2576), .Y(
        csr_io_decode_0_write_illegal) );
  OR2X1_LVT csr_U2258 ( .A1(ibuf_io_inst_0_bits_raw[22]), .A2(csr_n1426), .Y(
        csr_io_decode_0_write_flush) );
  NAND3X0_LVT csr_U2257 ( .A1(csr_n1366), .A2(csr_n1401), .A3(csr_n1365), .Y(
        csr_io_decode_0_system_illegal) );
  NAND2X0_LVT csr_U2256 ( .A1(csr_n490), .A2(n9516), .Y(csr_n1365) );
  OA22X1_LVT csr_U2255 ( .A1(io_ptw_status_prv[1]), .A2(csr_n1383), .A3(
        csr_n1364), .A4(csr_n1363), .Y(csr_n1401) );
  NOR2X0_LVT csr_U2254 ( .A1(csr_n381), .A2(ibuf_io_inst_0_bits_inst_rs3_2_), 
        .Y(csr_n1363) );
  NAND2X0_LVT csr_U2253 ( .A1(csr_n429), .A2(ibuf_io_inst_0_bits_raw[28]), .Y(
        csr_n1364) );
  INVX1_LVT csr_U2252 ( .A(ibuf_io_inst_0_bits_inst_rs3_2_), .Y(csr_n1383) );
  AO21X1_LVT csr_U2251 ( .A1(csr_n1362), .A2(csr_n1361), .A3(
        io_ptw_status_prv[1]), .Y(csr_n1366) );
  MUX21X1_LVT csr_U2250 ( .A1(csr_n1360), .A2(csr_n1359), .S0(csr_n1406), .Y(
        csr_n1361) );
  NAND2X0_LVT csr_U2249 ( .A1(csr_n1358), .A2(ibuf_io_inst_0_bits_raw[28]), 
        .Y(csr_n1359) );
  AO22X1_LVT csr_U2248 ( .A1(csr_n1407), .A2(csr_n1925), .A3(csr_n1924), .A4(
        csr_n1417), .Y(csr_n1358) );
  OR2X1_LVT csr_U2247 ( .A1(csr_n447), .A2(csr_n490), .Y(csr_n1360) );
  NAND2X0_LVT csr_U2246 ( .A1(csr_n490), .A2(csr_n1924), .Y(csr_n1362) );
  NAND3X0_LVT csr_U2245 ( .A1(csr_n1357), .A2(csr_n1354), .A3(csr_n1353), .Y(
        csr_io_evec[38]) );
  NAND2X0_LVT csr_U2244 ( .A1(csr_n502), .A2(csr_reg_mepc_38_), .Y(csr_n1353)
         );
  AOI22X1_LVT csr_U2243 ( .A1(csr_n1356), .A2(csr_reg_dpc_38_), .A3(csr_n500), 
        .A4(csr_reg_sepc_38_), .Y(csr_n1354) );
  OR2X1_LVT csr_U2242 ( .A1(csr_n465), .A2(csr_n1352), .Y(csr_n1357) );
  NAND3X0_LVT csr_U2241 ( .A1(csr_n1351), .A2(csr_n1350), .A3(csr_n1349), .Y(
        csr_io_evec[37]) );
  NAND2X0_LVT csr_U2240 ( .A1(csr_n502), .A2(csr_reg_mepc_37_), .Y(csr_n1349)
         );
  AOI22X1_LVT csr_U2239 ( .A1(csr_n1356), .A2(csr_reg_dpc_37_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_37_), .Y(csr_n1350) );
  NAND2X0_LVT csr_U2238 ( .A1(csr_n499), .A2(csr_reg_stvec_37_), .Y(csr_n1351)
         );
  NAND3X0_LVT csr_U2237 ( .A1(csr_n1347), .A2(csr_n1345), .A3(csr_n1344), .Y(
        csr_io_evec[35]) );
  NAND2X0_LVT csr_U2236 ( .A1(csr_n502), .A2(csr_reg_mepc_35_), .Y(csr_n1344)
         );
  AOI22X1_LVT csr_U2235 ( .A1(csr_n1356), .A2(csr_reg_dpc_35_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_35_), .Y(csr_n1345) );
  NAND2X0_LVT csr_U2234 ( .A1(csr_n499), .A2(csr_reg_stvec_35_), .Y(csr_n1347)
         );
  NAND3X0_LVT csr_U2233 ( .A1(csr_n1343), .A2(csr_n1342), .A3(csr_n1341), .Y(
        csr_io_evec[33]) );
  NAND2X0_LVT csr_U2232 ( .A1(csr_n502), .A2(csr_reg_mepc_33_), .Y(csr_n1341)
         );
  AOI22X1_LVT csr_U2231 ( .A1(csr_n1356), .A2(csr_reg_dpc_33_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_33_), .Y(csr_n1342) );
  NAND2X0_LVT csr_U2230 ( .A1(csr_n499), .A2(csr_reg_stvec_33_), .Y(csr_n1343)
         );
  NAND3X0_LVT csr_U2229 ( .A1(csr_n1340), .A2(csr_n1339), .A3(csr_n1338), .Y(
        csr_io_evec[32]) );
  NAND2X0_LVT csr_U2228 ( .A1(csr_n502), .A2(csr_reg_mepc_32_), .Y(csr_n1338)
         );
  AOI22X1_LVT csr_U2227 ( .A1(csr_n1356), .A2(csr_reg_dpc_32_), .A3(csr_n500), 
        .A4(csr_reg_sepc_32_), .Y(csr_n1339) );
  NAND2X0_LVT csr_U2226 ( .A1(csr_n499), .A2(csr_reg_stvec_32_), .Y(csr_n1340)
         );
  NAND4X0_LVT csr_U2225 ( .A1(csr_n1337), .A2(csr_n1336), .A3(csr_n1335), .A4(
        csr_n1334), .Y(csr_io_evec[31]) );
  NAND2X0_LVT csr_U2224 ( .A1(csr_n502), .A2(csr_reg_mepc_31_), .Y(csr_n1334)
         );
  NAND2X0_LVT csr_U2223 ( .A1(csr_n1333), .A2(csr_reg_mtvec_31_), .Y(csr_n1335) );
  AOI22X1_LVT csr_U2222 ( .A1(csr_n1356), .A2(csr_reg_dpc_31_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_31_), .Y(csr_n1336) );
  NAND2X0_LVT csr_U2221 ( .A1(csr_n499), .A2(csr_reg_stvec_31_), .Y(csr_n1337)
         );
  NAND4X0_LVT csr_U2220 ( .A1(csr_n1332), .A2(csr_n1331), .A3(csr_n1330), .A4(
        csr_n1329), .Y(csr_io_evec[29]) );
  NAND2X0_LVT csr_U2219 ( .A1(csr_n502), .A2(csr_reg_mepc_29_), .Y(csr_n1329)
         );
  NAND2X0_LVT csr_U2218 ( .A1(csr_n1333), .A2(csr_reg_mtvec_29_), .Y(csr_n1330) );
  AOI22X1_LVT csr_U2217 ( .A1(csr_n1356), .A2(csr_reg_dpc_29_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_29_), .Y(csr_n1331) );
  NAND2X0_LVT csr_U2216 ( .A1(csr_n499), .A2(csr_reg_stvec_29_), .Y(csr_n1332)
         );
  NAND4X0_LVT csr_U2215 ( .A1(csr_n1328), .A2(csr_n1327), .A3(csr_n1326), .A4(
        csr_n1325), .Y(csr_io_evec[28]) );
  NAND2X0_LVT csr_U2214 ( .A1(csr_n502), .A2(csr_reg_mepc_28_), .Y(csr_n1325)
         );
  NAND2X0_LVT csr_U2213 ( .A1(csr_n1333), .A2(csr_reg_mtvec_28_), .Y(csr_n1326) );
  AOI22X1_LVT csr_U2212 ( .A1(csr_n1356), .A2(csr_reg_dpc_28_), .A3(csr_n500), 
        .A4(csr_reg_sepc_28_), .Y(csr_n1327) );
  NAND2X0_LVT csr_U2211 ( .A1(csr_n499), .A2(csr_reg_stvec_28_), .Y(csr_n1328)
         );
  NAND4X0_LVT csr_U2210 ( .A1(csr_n1324), .A2(csr_n1323), .A3(csr_n1322), .A4(
        csr_n1321), .Y(csr_io_evec[27]) );
  NAND2X0_LVT csr_U2209 ( .A1(csr_n502), .A2(csr_reg_mepc_27_), .Y(csr_n1321)
         );
  NAND2X0_LVT csr_U2208 ( .A1(csr_n1333), .A2(csr_reg_mtvec_27_), .Y(csr_n1322) );
  AOI22X1_LVT csr_U2207 ( .A1(csr_n1356), .A2(csr_reg_dpc_27_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_27_), .Y(csr_n1323) );
  NAND2X0_LVT csr_U2206 ( .A1(csr_n499), .A2(csr_reg_stvec_27_), .Y(csr_n1324)
         );
  NAND4X0_LVT csr_U2205 ( .A1(csr_n1320), .A2(csr_n1319), .A3(csr_n1318), .A4(
        csr_n1317), .Y(csr_io_evec[26]) );
  NAND2X0_LVT csr_U2204 ( .A1(csr_n502), .A2(csr_reg_mepc_26_), .Y(csr_n1317)
         );
  NAND2X0_LVT csr_U2203 ( .A1(csr_n1333), .A2(csr_reg_mtvec_26_), .Y(csr_n1318) );
  AOI22X1_LVT csr_U2202 ( .A1(csr_n1356), .A2(csr_reg_dpc_26_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_26_), .Y(csr_n1319) );
  NAND2X0_LVT csr_U2201 ( .A1(csr_n499), .A2(csr_reg_stvec_26_), .Y(csr_n1320)
         );
  NAND4X0_LVT csr_U2200 ( .A1(csr_n1316), .A2(csr_n1315), .A3(csr_n1314), .A4(
        csr_n1313), .Y(csr_io_evec[25]) );
  NAND2X0_LVT csr_U2199 ( .A1(csr_n502), .A2(csr_reg_mepc_25_), .Y(csr_n1313)
         );
  NAND2X0_LVT csr_U2198 ( .A1(csr_n1333), .A2(csr_reg_mtvec_25_), .Y(csr_n1314) );
  AOI22X1_LVT csr_U2197 ( .A1(csr_n1356), .A2(csr_reg_dpc_25_), .A3(csr_n500), 
        .A4(csr_reg_sepc_25_), .Y(csr_n1315) );
  NAND2X0_LVT csr_U2196 ( .A1(csr_n499), .A2(csr_reg_stvec_25_), .Y(csr_n1316)
         );
  NAND4X0_LVT csr_U2195 ( .A1(csr_n1312), .A2(csr_n1311), .A3(csr_n1310), .A4(
        csr_n1309), .Y(csr_io_evec[24]) );
  NAND2X0_LVT csr_U2194 ( .A1(csr_n502), .A2(csr_reg_mepc_24_), .Y(csr_n1309)
         );
  NAND2X0_LVT csr_U2193 ( .A1(csr_n1333), .A2(csr_reg_mtvec_24_), .Y(csr_n1310) );
  AOI22X1_LVT csr_U2192 ( .A1(csr_n1356), .A2(csr_reg_dpc_24_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_24_), .Y(csr_n1311) );
  NAND2X0_LVT csr_U2191 ( .A1(csr_n499), .A2(csr_reg_stvec_24_), .Y(csr_n1312)
         );
  NAND4X0_LVT csr_U2190 ( .A1(csr_n1308), .A2(csr_n1307), .A3(csr_n1306), .A4(
        csr_n1305), .Y(csr_io_evec[23]) );
  NAND2X0_LVT csr_U2189 ( .A1(csr_n502), .A2(csr_reg_mepc_23_), .Y(csr_n1305)
         );
  NAND2X0_LVT csr_U2188 ( .A1(csr_n1333), .A2(csr_reg_mtvec_23_), .Y(csr_n1306) );
  AOI22X1_LVT csr_U2187 ( .A1(csr_n1356), .A2(csr_reg_dpc_23_), .A3(csr_n500), 
        .A4(csr_reg_sepc_23_), .Y(csr_n1307) );
  NAND2X0_LVT csr_U2186 ( .A1(csr_n499), .A2(csr_reg_stvec_23_), .Y(csr_n1308)
         );
  NAND4X0_LVT csr_U2185 ( .A1(csr_n1304), .A2(csr_n1303), .A3(csr_n1302), .A4(
        csr_n1301), .Y(csr_io_evec[22]) );
  NAND2X0_LVT csr_U2184 ( .A1(csr_n502), .A2(csr_reg_mepc_22_), .Y(csr_n1301)
         );
  NAND2X0_LVT csr_U2183 ( .A1(csr_n1333), .A2(csr_reg_mtvec_22_), .Y(csr_n1302) );
  AOI22X1_LVT csr_U2182 ( .A1(csr_n1356), .A2(csr_reg_dpc_22_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_22_), .Y(csr_n1303) );
  NAND2X0_LVT csr_U2181 ( .A1(csr_n499), .A2(csr_reg_stvec_22_), .Y(csr_n1304)
         );
  NAND4X0_LVT csr_U2180 ( .A1(csr_n1300), .A2(csr_n1299), .A3(csr_n1298), .A4(
        csr_n1297), .Y(csr_io_evec[21]) );
  NAND2X0_LVT csr_U2179 ( .A1(csr_n502), .A2(csr_reg_mepc_21_), .Y(csr_n1297)
         );
  NAND2X0_LVT csr_U2178 ( .A1(csr_n1333), .A2(csr_reg_mtvec_21_), .Y(csr_n1298) );
  AOI22X1_LVT csr_U2177 ( .A1(csr_n1356), .A2(csr_reg_dpc_21_), .A3(csr_n500), 
        .A4(csr_reg_sepc_21_), .Y(csr_n1299) );
  NAND2X0_LVT csr_U2176 ( .A1(csr_n1348), .A2(csr_reg_stvec_21_), .Y(csr_n1300) );
  NAND4X0_LVT csr_U2175 ( .A1(csr_n1296), .A2(csr_n1295), .A3(csr_n1294), .A4(
        csr_n1293), .Y(csr_io_evec[20]) );
  NAND2X0_LVT csr_U2174 ( .A1(csr_n502), .A2(csr_reg_mepc_20_), .Y(csr_n1293)
         );
  NAND2X0_LVT csr_U2173 ( .A1(csr_n1333), .A2(csr_reg_mtvec_20_), .Y(csr_n1294) );
  AOI22X1_LVT csr_U2172 ( .A1(csr_n1356), .A2(csr_reg_dpc_20_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_20_), .Y(csr_n1295) );
  NAND2X0_LVT csr_U2171 ( .A1(csr_n1348), .A2(csr_reg_stvec_20_), .Y(csr_n1296) );
  NAND4X0_LVT csr_U2170 ( .A1(csr_n1292), .A2(csr_n1291), .A3(csr_n1290), .A4(
        csr_n1289), .Y(csr_io_evec[19]) );
  NAND2X0_LVT csr_U2169 ( .A1(csr_n502), .A2(csr_reg_mepc_19_), .Y(csr_n1289)
         );
  NAND2X0_LVT csr_U2168 ( .A1(csr_n1333), .A2(csr_reg_mtvec_19_), .Y(csr_n1290) );
  AOI22X1_LVT csr_U2167 ( .A1(csr_n1356), .A2(csr_reg_dpc_19_), .A3(csr_n500), 
        .A4(csr_reg_sepc_19_), .Y(csr_n1291) );
  NAND2X0_LVT csr_U2166 ( .A1(csr_n1348), .A2(csr_reg_stvec_19_), .Y(csr_n1292) );
  NAND4X0_LVT csr_U2165 ( .A1(csr_n1288), .A2(csr_n1287), .A3(csr_n1286), .A4(
        csr_n1285), .Y(csr_io_evec[18]) );
  NAND2X0_LVT csr_U2164 ( .A1(csr_n502), .A2(csr_reg_mepc_18_), .Y(csr_n1285)
         );
  NAND2X0_LVT csr_U2163 ( .A1(csr_n1333), .A2(csr_reg_mtvec_18_), .Y(csr_n1286) );
  AOI22X1_LVT csr_U2162 ( .A1(csr_n1356), .A2(csr_reg_dpc_18_), .A3(csr_n500), 
        .A4(csr_reg_sepc_18_), .Y(csr_n1287) );
  NAND2X0_LVT csr_U2161 ( .A1(csr_n1348), .A2(csr_reg_stvec_18_), .Y(csr_n1288) );
  NAND4X0_LVT csr_U2160 ( .A1(csr_n1284), .A2(csr_n1283), .A3(csr_n1282), .A4(
        csr_n1281), .Y(csr_io_evec[17]) );
  NAND2X0_LVT csr_U2159 ( .A1(csr_n502), .A2(csr_reg_mepc_17_), .Y(csr_n1281)
         );
  NAND2X0_LVT csr_U2158 ( .A1(csr_n1333), .A2(csr_reg_mtvec_17_), .Y(csr_n1282) );
  AOI22X1_LVT csr_U2157 ( .A1(csr_n1356), .A2(csr_reg_dpc_17_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_17_), .Y(csr_n1283) );
  NAND2X0_LVT csr_U2156 ( .A1(csr_n1348), .A2(csr_reg_stvec_17_), .Y(csr_n1284) );
  NAND4X0_LVT csr_U2155 ( .A1(csr_n1280), .A2(csr_n1279), .A3(csr_n1278), .A4(
        csr_n1277), .Y(csr_io_evec[16]) );
  NAND2X0_LVT csr_U2154 ( .A1(csr_n502), .A2(csr_reg_mepc_16_), .Y(csr_n1277)
         );
  NAND2X0_LVT csr_U2153 ( .A1(csr_n1333), .A2(csr_reg_mtvec_16_), .Y(csr_n1278) );
  AOI22X1_LVT csr_U2152 ( .A1(csr_n1356), .A2(csr_reg_dpc_16_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_16_), .Y(csr_n1279) );
  NAND2X0_LVT csr_U2151 ( .A1(csr_n1348), .A2(csr_reg_stvec_16_), .Y(csr_n1280) );
  NAND4X0_LVT csr_U2150 ( .A1(csr_n1276), .A2(csr_n1275), .A3(csr_n1274), .A4(
        csr_n1273), .Y(csr_io_evec[15]) );
  NAND2X0_LVT csr_U2149 ( .A1(csr_n502), .A2(csr_reg_mepc_15_), .Y(csr_n1273)
         );
  NAND2X0_LVT csr_U2148 ( .A1(csr_n1333), .A2(csr_reg_mtvec_15_), .Y(csr_n1274) );
  AOI22X1_LVT csr_U2147 ( .A1(csr_n1356), .A2(csr_reg_dpc_15_), .A3(csr_n500), 
        .A4(csr_reg_sepc_15_), .Y(csr_n1275) );
  NAND2X0_LVT csr_U2146 ( .A1(csr_n1348), .A2(csr_reg_stvec_15_), .Y(csr_n1276) );
  NAND4X0_LVT csr_U2145 ( .A1(csr_n1272), .A2(csr_n1271), .A3(csr_n1270), .A4(
        csr_n1269), .Y(csr_io_evec[14]) );
  NAND2X0_LVT csr_U2144 ( .A1(csr_n502), .A2(csr_reg_mepc_14_), .Y(csr_n1269)
         );
  NAND2X0_LVT csr_U2143 ( .A1(csr_n1333), .A2(csr_reg_mtvec_14_), .Y(csr_n1270) );
  AOI22X1_LVT csr_U2142 ( .A1(csr_n1356), .A2(csr_reg_dpc_14_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_14_), .Y(csr_n1271) );
  NAND2X0_LVT csr_U2141 ( .A1(csr_n1348), .A2(csr_reg_stvec_14_), .Y(csr_n1272) );
  NAND4X0_LVT csr_U2140 ( .A1(csr_n1268), .A2(csr_n1267), .A3(csr_n1266), .A4(
        csr_n1265), .Y(csr_io_evec[13]) );
  NAND2X0_LVT csr_U2139 ( .A1(csr_n502), .A2(csr_reg_mepc_13_), .Y(csr_n1265)
         );
  NAND2X0_LVT csr_U2138 ( .A1(csr_n1333), .A2(csr_reg_mtvec_13_), .Y(csr_n1266) );
  AOI22X1_LVT csr_U2137 ( .A1(csr_n1356), .A2(csr_reg_dpc_13_), .A3(csr_n500), 
        .A4(csr_reg_sepc_13_), .Y(csr_n1267) );
  NAND2X0_LVT csr_U2136 ( .A1(csr_n1348), .A2(csr_reg_stvec_13_), .Y(csr_n1268) );
  NAND4X0_LVT csr_U2135 ( .A1(csr_n1264), .A2(csr_n1263), .A3(csr_n1262), .A4(
        csr_n1261), .Y(csr_io_evec[12]) );
  NAND2X0_LVT csr_U2134 ( .A1(csr_n502), .A2(csr_reg_mepc_12_), .Y(csr_n1261)
         );
  NAND2X0_LVT csr_U2133 ( .A1(csr_n1333), .A2(csr_reg_mtvec_12_), .Y(csr_n1262) );
  AOI22X1_LVT csr_U2132 ( .A1(csr_n1356), .A2(csr_reg_dpc_12_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_12_), .Y(csr_n1263) );
  NAND2X0_LVT csr_U2131 ( .A1(csr_n1348), .A2(csr_reg_stvec_12_), .Y(csr_n1264) );
  OR3X1_LVT csr_U2130 ( .A1(csr_n1260), .A2(csr_n1259), .A3(csr_n1258), .Y(
        csr_io_evec[11]) );
  OA21X1_LVT csr_U2129 ( .A1(csr_n1257), .A2(csr_n1256), .A3(csr_n1903), .Y(
        csr_n1258) );
  MUX21X1_LVT csr_U2128 ( .A1(csr_reg_stvec_11_), .A2(csr_reg_mtvec_11_), .S0(
        csr_n1255), .Y(csr_n1256) );
  AO22X1_LVT csr_U2127 ( .A1(csr_n1356), .A2(csr_reg_dpc_11_), .A3(csr_n500), 
        .A4(csr_reg_sepc_11_), .Y(csr_n1259) );
  AND2X1_LVT csr_U2126 ( .A1(csr_n502), .A2(csr_reg_mepc_11_), .Y(csr_n1260)
         );
  NAND4X0_LVT csr_U2125 ( .A1(csr_n1254), .A2(csr_n1253), .A3(csr_n1252), .A4(
        csr_n1251), .Y(csr_io_evec[10]) );
  NAND2X0_LVT csr_U2124 ( .A1(csr_n502), .A2(csr_reg_mepc_10_), .Y(csr_n1251)
         );
  NAND2X0_LVT csr_U2123 ( .A1(csr_n1333), .A2(csr_reg_mtvec_10_), .Y(csr_n1252) );
  AOI22X1_LVT csr_U2122 ( .A1(csr_n1356), .A2(csr_reg_dpc_10_), .A3(csr_n500), 
        .A4(csr_reg_sepc_10_), .Y(csr_n1253) );
  NAND2X0_LVT csr_U2121 ( .A1(csr_n1348), .A2(csr_reg_stvec_10_), .Y(csr_n1254) );
  NAND4X0_LVT csr_U2120 ( .A1(csr_n1250), .A2(csr_n1249), .A3(csr_n1248), .A4(
        csr_n1247), .Y(csr_io_evec[9]) );
  NAND2X0_LVT csr_U2119 ( .A1(csr_n502), .A2(csr_reg_mepc_9_), .Y(csr_n1247)
         );
  NAND2X0_LVT csr_U2118 ( .A1(csr_n1333), .A2(csr_reg_mtvec_9_), .Y(csr_n1248)
         );
  AOI22X1_LVT csr_U2117 ( .A1(csr_n1356), .A2(csr_reg_dpc_9_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_9_), .Y(csr_n1249) );
  NAND2X0_LVT csr_U2116 ( .A1(csr_n1348), .A2(csr_reg_stvec_9_), .Y(csr_n1250)
         );
  NAND4X0_LVT csr_U2115 ( .A1(csr_n1246), .A2(csr_n1245), .A3(csr_n1244), .A4(
        csr_n1243), .Y(csr_io_evec[8]) );
  NAND2X0_LVT csr_U2114 ( .A1(csr_n502), .A2(csr_reg_mepc_8_), .Y(csr_n1243)
         );
  NAND2X0_LVT csr_U2113 ( .A1(csr_n1333), .A2(csr_reg_mtvec_8_), .Y(csr_n1244)
         );
  AOI22X1_LVT csr_U2112 ( .A1(csr_n1356), .A2(csr_reg_dpc_8_), .A3(csr_n500), 
        .A4(csr_reg_sepc_8_), .Y(csr_n1245) );
  NAND2X0_LVT csr_U2111 ( .A1(csr_n1348), .A2(csr_reg_stvec_8_), .Y(csr_n1246)
         );
  NAND2X0_LVT csr_U2110 ( .A1(csr_n1239), .A2(csr_reg_mtvec_7_), .Y(csr_n1240)
         );
  NAND2X0_LVT csr_U2109 ( .A1(csr_n1238), .A2(csr_reg_stvec_7_), .Y(csr_n1241)
         );
  AOI21X1_LVT csr_U2108 ( .A1(csr_n502), .A2(csr_reg_mepc_7_), .A3(csr_n1237), 
        .Y(csr_n1242) );
  AO22X1_LVT csr_U2107 ( .A1(csr_n1356), .A2(csr_reg_dpc_7_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_7_), .Y(csr_n1237) );
  NAND2X0_LVT csr_U2106 ( .A1(csr_n1239), .A2(csr_reg_mtvec_6_), .Y(csr_n1233)
         );
  NAND2X0_LVT csr_U2105 ( .A1(csr_n1238), .A2(csr_reg_stvec_6_), .Y(csr_n1234)
         );
  AOI21X1_LVT csr_U2104 ( .A1(csr_n502), .A2(csr_reg_mepc_6_), .A3(csr_n1232), 
        .Y(csr_n1235) );
  AO22X1_LVT csr_U2103 ( .A1(csr_n1356), .A2(csr_reg_dpc_6_), .A3(csr_n500), 
        .A4(csr_reg_sepc_6_), .Y(csr_n1232) );
  NAND4X0_LVT csr_U2102 ( .A1(csr_n1231), .A2(csr_n1230), .A3(csr_n1229), .A4(
        csr_n1228), .Y(csr_io_evec[5]) );
  NAND2X0_LVT csr_U2101 ( .A1(csr_n1239), .A2(csr_reg_mtvec_5_), .Y(csr_n1228)
         );
  NAND2X0_LVT csr_U2100 ( .A1(csr_n1238), .A2(csr_reg_stvec_5_), .Y(csr_n1229)
         );
  AOI21X1_LVT csr_U2099 ( .A1(csr_n502), .A2(csr_reg_mepc_5_), .A3(csr_n1227), 
        .Y(csr_n1230) );
  AO22X1_LVT csr_U2098 ( .A1(csr_n1356), .A2(csr_reg_dpc_5_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_5_), .Y(csr_n1227) );
  NAND2X0_LVT csr_U2097 ( .A1(csr_n1236), .A2(csr_n1226), .Y(csr_n1231) );
  NAND4X0_LVT csr_U2096 ( .A1(csr_n1225), .A2(csr_n1224), .A3(csr_n1223), .A4(
        csr_n1222), .Y(csr_io_evec[4]) );
  NAND2X0_LVT csr_U2095 ( .A1(csr_n1239), .A2(csr_reg_mtvec_4_), .Y(csr_n1222)
         );
  NAND2X0_LVT csr_U2094 ( .A1(csr_n1238), .A2(csr_reg_stvec_4_), .Y(csr_n1223)
         );
  AOI21X1_LVT csr_U2093 ( .A1(csr_n502), .A2(csr_reg_mepc_4_), .A3(csr_n1221), 
        .Y(csr_n1224) );
  AO22X1_LVT csr_U2092 ( .A1(csr_n1356), .A2(csr_reg_dpc_4_), .A3(csr_n500), 
        .A4(csr_reg_sepc_4_), .Y(csr_n1221) );
  NAND2X0_LVT csr_U2091 ( .A1(csr_n1236), .A2(csr_n1220), .Y(csr_n1225) );
  NAND4X0_LVT csr_U2090 ( .A1(csr_n1219), .A2(csr_n1218), .A3(csr_n1217), .A4(
        csr_n1216), .Y(csr_io_evec[3]) );
  NAND2X0_LVT csr_U2089 ( .A1(csr_n1239), .A2(csr_reg_mtvec_3_), .Y(csr_n1216)
         );
  NAND2X0_LVT csr_U2088 ( .A1(csr_n1238), .A2(csr_reg_stvec_3_), .Y(csr_n1217)
         );
  AND4X1_LVT csr_U2087 ( .A1(csr_n1215), .A2(csr_n1214), .A3(csr_n1213), .A4(
        csr_n1212), .Y(csr_n1218) );
  NAND3X0_LVT csr_U2086 ( .A1(csr_n1211), .A2(csr_io_status_debug), .A3(
        csr_n1903), .Y(csr_n1212) );
  NAND2X0_LVT csr_U2085 ( .A1(csr_n1356), .A2(csr_reg_dpc_3_), .Y(csr_n1213)
         );
  NAND2X0_LVT csr_U2084 ( .A1(csr_reg_mepc_3_), .A2(csr_n502), .Y(csr_n1214)
         );
  NAND2X0_LVT csr_U2083 ( .A1(csr_reg_sepc_3_), .A2(csr_n500), .Y(csr_n1215)
         );
  NAND2X0_LVT csr_U2082 ( .A1(csr_n1236), .A2(csr_n1209), .Y(csr_n1219) );
  NAND4X0_LVT csr_U2081 ( .A1(csr_n1208), .A2(csr_n1207), .A3(csr_n1206), .A4(
        csr_n1205), .Y(csr_io_evec[2]) );
  NAND2X0_LVT csr_U2080 ( .A1(csr_n1239), .A2(csr_reg_mtvec_2_), .Y(csr_n1205)
         );
  AND2X1_LVT csr_U2079 ( .A1(csr_n1333), .A2(csr_n659), .Y(csr_n1239) );
  NAND2X0_LVT csr_U2078 ( .A1(csr_n1238), .A2(csr_reg_stvec_2_), .Y(csr_n1206)
         );
  AND2X1_LVT csr_U2077 ( .A1(csr_n1348), .A2(csr_n658), .Y(csr_n1238) );
  AOI21X1_LVT csr_U2076 ( .A1(csr_n502), .A2(csr_reg_mepc_2_), .A3(csr_n1203), 
        .Y(csr_n1207) );
  AO22X1_LVT csr_U2075 ( .A1(csr_n1356), .A2(csr_reg_dpc_2_), .A3(csr_n1355), 
        .A4(csr_reg_sepc_2_), .Y(csr_n1203) );
  NAND2X0_LVT csr_U2074 ( .A1(csr_n1236), .A2(csr_n1202), .Y(csr_n1208) );
  AND2X1_LVT csr_U2073 ( .A1(csr_n1201), .A2(csr_n1200), .Y(csr_n1236) );
  OAI22X1_LVT csr_U2072 ( .A1(csr_n659), .A2(csr_n1204), .A3(csr_n658), .A4(
        csr_n1352), .Y(csr_n1200) );
  NAND3X0_LVT csr_U2071 ( .A1(csr_n1255), .A2(csr_n1198), .A3(csr_n1903), .Y(
        csr_n1204) );
  AND2X1_LVT csr_U2070 ( .A1(csr_io_status_isa[2]), .A2(csr_n1197), .Y(
        csr_io_evec[1]) );
  AO222X1_LVT csr_U2069 ( .A1(csr_n502), .A2(csr_reg_mepc_1_), .A3(csr_n1356), 
        .A4(csr_reg_dpc_1_), .A5(csr_n1355), .A6(csr_reg_sepc_1_), .Y(
        csr_n1197) );
  OA21X1_LVT csr_U2068 ( .A1(csr_n426), .A2(csr_n1196), .A3(csr_n1195), .Y(
        csr_io_interrupt) );
  NOR2X0_LVT csr_U2067 ( .A1(csr_io_status_debug), .A2(csr_n1918), .Y(
        csr_n1195) );
  OA21X1_LVT csr_U2066 ( .A1(io_interrupts_debug), .A2(csr_n1194), .A3(
        csr_n452), .Y(csr_n1196) );
  OR3X1_LVT csr_U2065 ( .A1(io_interrupts_debug), .A2(csr_n1184), .A3(
        csr_n1180), .Y(csr_io_interrupt_cause[1]) );
  NAND3X0_LVT csr_U2064 ( .A1(csr_n1177), .A2(csr_n407), .A3(csr_n1176), .Y(
        csr_n1190) );
  NAND2X0_LVT csr_U2063 ( .A1(csr_n1176), .A2(csr_n1173), .Y(csr_n1192) );
  NOR3X0_LVT csr_U2062 ( .A1(csr_read_mideleg_9_), .A2(csr_n1187), .A3(
        csr_n1171), .Y(csr_n1189) );
  AND2X1_LVT csr_U2061 ( .A1(csr_n1181), .A2(csr_n1170), .Y(csr_n1191) );
  AND2X1_LVT csr_U2060 ( .A1(csr_n1174), .A2(csr_n1175), .Y(csr_n1181) );
  OA21X1_LVT csr_U2059 ( .A1(csr_n1935), .A2(csr_n429), .A3(csr_n381), .Y(
        csr_n1175) );
  NAND3X0_LVT csr_U2058 ( .A1(csr_n1169), .A2(csr_n427), .A3(csr_n1176), .Y(
        csr_n1174) );
  NAND2X0_LVT csr_U2057 ( .A1(csr_n383), .A2(io_ptw_status_prv[1]), .Y(
        csr_n1176) );
  NOR2X0_LVT csr_U2056 ( .A1(csr_n_T_241[12]), .A2(csr_n406), .Y(
        io_ptw_pmp_0_mask[14]) );
  NOR2X0_LVT csr_U2055 ( .A1(csr_n_T_241[10]), .A2(csr_n419), .Y(
        io_ptw_pmp_0_mask[12]) );
  NOR2X0_LVT csr_U2054 ( .A1(csr_n_T_241[8]), .A2(csr_n398), .Y(
        io_ptw_pmp_0_mask[10]) );
  NOR2X0_LVT csr_U2053 ( .A1(csr_n_T_241[4]), .A2(csr_n415), .Y(
        io_ptw_pmp_0_mask[6]) );
  NOR2X0_LVT csr_U2052 ( .A1(csr_n_T_250[12]), .A2(csr_n402), .Y(
        io_ptw_pmp_1_mask[14]) );
  NOR2X0_LVT csr_U2051 ( .A1(csr_n_T_250[10]), .A2(csr_n425), .Y(
        io_ptw_pmp_1_mask[12]) );
  NOR2X0_LVT csr_U2050 ( .A1(csr_n_T_250[8]), .A2(csr_n397), .Y(
        io_ptw_pmp_1_mask[10]) );
  NOR2X0_LVT csr_U2049 ( .A1(csr_n_T_250[4]), .A2(csr_n411), .Y(
        io_ptw_pmp_1_mask[6]) );
  NOR2X0_LVT csr_U2048 ( .A1(csr_n_T_259[12]), .A2(csr_n405), .Y(
        io_ptw_pmp_2_mask[14]) );
  NOR2X0_LVT csr_U2047 ( .A1(csr_n_T_259[10]), .A2(csr_n421), .Y(
        io_ptw_pmp_2_mask[12]) );
  NOR2X0_LVT csr_U2046 ( .A1(csr_n_T_259[8]), .A2(csr_n393), .Y(
        io_ptw_pmp_2_mask[10]) );
  NOR2X0_LVT csr_U2045 ( .A1(csr_n_T_259[4]), .A2(csr_n410), .Y(
        io_ptw_pmp_2_mask[6]) );
  NOR2X0_LVT csr_U2044 ( .A1(csr_n_T_268[12]), .A2(csr_n401), .Y(
        io_ptw_pmp_3_mask[14]) );
  NOR2X0_LVT csr_U2043 ( .A1(csr_n_T_268[10]), .A2(csr_n418), .Y(
        io_ptw_pmp_3_mask[12]) );
  NOR2X0_LVT csr_U2042 ( .A1(csr_n_T_268[8]), .A2(csr_n396), .Y(
        io_ptw_pmp_3_mask[10]) );
  NOR2X0_LVT csr_U2041 ( .A1(csr_n_T_268[4]), .A2(csr_n409), .Y(
        io_ptw_pmp_3_mask[6]) );
  NOR2X0_LVT csr_U2040 ( .A1(csr_n_T_277[12]), .A2(csr_n400), .Y(
        io_ptw_pmp_4_mask[14]) );
  NOR2X0_LVT csr_U2039 ( .A1(csr_n_T_277[10]), .A2(csr_n423), .Y(
        io_ptw_pmp_4_mask[12]) );
  NOR2X0_LVT csr_U2038 ( .A1(csr_n_T_277[8]), .A2(csr_n395), .Y(
        io_ptw_pmp_4_mask[10]) );
  NOR2X0_LVT csr_U2037 ( .A1(csr_n_T_277[4]), .A2(csr_n408), .Y(
        io_ptw_pmp_4_mask[6]) );
  NOR2X0_LVT csr_U2036 ( .A1(csr_n_T_286[12]), .A2(csr_n399), .Y(
        io_ptw_pmp_5_mask[14]) );
  NOR2X0_LVT csr_U2035 ( .A1(csr_n_T_286[10]), .A2(csr_n422), .Y(
        io_ptw_pmp_5_mask[12]) );
  NOR2X0_LVT csr_U2034 ( .A1(csr_n_T_286[8]), .A2(csr_n392), .Y(
        io_ptw_pmp_5_mask[10]) );
  NOR2X0_LVT csr_U2033 ( .A1(csr_n_T_286[4]), .A2(csr_n414), .Y(
        io_ptw_pmp_5_mask[6]) );
  NOR2X0_LVT csr_U2032 ( .A1(csr_n_T_295[12]), .A2(csr_n404), .Y(
        io_ptw_pmp_6_mask[14]) );
  NOR2X0_LVT csr_U2031 ( .A1(csr_n_T_295[10]), .A2(csr_n420), .Y(
        io_ptw_pmp_6_mask[12]) );
  NOR2X0_LVT csr_U2030 ( .A1(csr_n_T_295[8]), .A2(csr_n391), .Y(
        io_ptw_pmp_6_mask[10]) );
  NOR2X0_LVT csr_U2029 ( .A1(csr_n_T_295[4]), .A2(csr_n413), .Y(
        io_ptw_pmp_6_mask[6]) );
  NOR2X0_LVT csr_U2028 ( .A1(csr_n_T_304[12]), .A2(csr_n403), .Y(
        io_ptw_pmp_7_mask[14]) );
  NOR2X0_LVT csr_U2027 ( .A1(csr_n_T_304[10]), .A2(csr_n424), .Y(
        io_ptw_pmp_7_mask[12]) );
  NOR2X0_LVT csr_U2026 ( .A1(csr_n_T_304[8]), .A2(csr_n394), .Y(
        io_ptw_pmp_7_mask[10]) );
  NOR2X0_LVT csr_U2025 ( .A1(csr_n_T_304[4]), .A2(csr_n412), .Y(
        io_ptw_pmp_7_mask[6]) );
  INVX1_LVT csr_U2024 ( .A(csr_n_T_304[7]), .Y(csr_n1897) );
  INVX1_LVT csr_U2023 ( .A(csr_n_T_304[6]), .Y(csr_n1896) );
  INVX1_LVT csr_U2022 ( .A(csr_n_T_304[5]), .Y(csr_n1895) );
  INVX1_LVT csr_U2021 ( .A(csr_n_T_304[3]), .Y(csr_n1894) );
  INVX1_LVT csr_U2020 ( .A(csr_n_T_304[2]), .Y(csr_n1893) );
  INVX1_LVT csr_U2019 ( .A(csr_n_T_304[1]), .Y(csr_n1892) );
  INVX1_LVT csr_U2018 ( .A(csr_n_T_304[29]), .Y(csr_n1891) );
  INVX1_LVT csr_U2017 ( .A(csr_n_T_304[28]), .Y(csr_n1890) );
  INVX1_LVT csr_U2016 ( .A(csr_n_T_304[27]), .Y(csr_n1889) );
  INVX1_LVT csr_U2015 ( .A(csr_n_T_304[26]), .Y(csr_n1888) );
  INVX1_LVT csr_U2014 ( .A(csr_n_T_304[25]), .Y(csr_n1887) );
  INVX1_LVT csr_U2013 ( .A(csr_n_T_304[24]), .Y(csr_n1886) );
  INVX1_LVT csr_U2012 ( .A(csr_n_T_304[23]), .Y(csr_n1885) );
  INVX1_LVT csr_U2011 ( .A(csr_n_T_304[22]), .Y(csr_n1884) );
  INVX1_LVT csr_U2010 ( .A(csr_n_T_304[21]), .Y(csr_n1883) );
  INVX1_LVT csr_U2009 ( .A(csr_n_T_304[20]), .Y(csr_n1882) );
  INVX1_LVT csr_U2008 ( .A(csr_n_T_304[19]), .Y(csr_n1881) );
  INVX1_LVT csr_U2007 ( .A(csr_n_T_304[18]), .Y(csr_n1880) );
  INVX1_LVT csr_U2006 ( .A(csr_n_T_304[17]), .Y(csr_n1879) );
  INVX1_LVT csr_U2005 ( .A(csr_n_T_304[16]), .Y(csr_n1878) );
  INVX1_LVT csr_U2004 ( .A(csr_n_T_304[15]), .Y(csr_n1877) );
  INVX1_LVT csr_U2003 ( .A(csr_n_T_304[14]), .Y(csr_n1876) );
  INVX1_LVT csr_U2002 ( .A(csr_n_T_304[13]), .Y(csr_n1875) );
  INVX1_LVT csr_U2001 ( .A(csr_n_T_304[11]), .Y(csr_n1874) );
  INVX1_LVT csr_U2000 ( .A(csr_n_T_304[9]), .Y(csr_n1873) );
  INVX1_LVT csr_U1999 ( .A(csr_n_T_295[7]), .Y(csr_n1872) );
  INVX1_LVT csr_U1998 ( .A(csr_n_T_295[6]), .Y(csr_n1871) );
  INVX1_LVT csr_U1997 ( .A(csr_n_T_295[5]), .Y(csr_n1870) );
  INVX1_LVT csr_U1996 ( .A(csr_n_T_295[3]), .Y(csr_n1869) );
  INVX1_LVT csr_U1995 ( .A(csr_n_T_295[2]), .Y(csr_n1868) );
  INVX1_LVT csr_U1994 ( .A(csr_n_T_295[1]), .Y(csr_n1867) );
  INVX1_LVT csr_U1993 ( .A(csr_n_T_295[29]), .Y(csr_n1866) );
  INVX1_LVT csr_U1992 ( .A(csr_n_T_295[28]), .Y(csr_n1865) );
  INVX1_LVT csr_U1991 ( .A(csr_n_T_295[27]), .Y(csr_n1864) );
  INVX1_LVT csr_U1990 ( .A(csr_n_T_295[26]), .Y(csr_n1863) );
  INVX1_LVT csr_U1989 ( .A(csr_n_T_295[25]), .Y(csr_n1862) );
  INVX1_LVT csr_U1988 ( .A(csr_n_T_295[24]), .Y(csr_n1861) );
  INVX1_LVT csr_U1987 ( .A(csr_n_T_295[23]), .Y(csr_n1860) );
  INVX1_LVT csr_U1986 ( .A(csr_n_T_295[22]), .Y(csr_n1859) );
  INVX1_LVT csr_U1985 ( .A(csr_n_T_295[21]), .Y(csr_n1858) );
  INVX1_LVT csr_U1984 ( .A(csr_n_T_295[20]), .Y(csr_n1857) );
  INVX1_LVT csr_U1983 ( .A(csr_n_T_295[19]), .Y(csr_n1856) );
  INVX1_LVT csr_U1982 ( .A(csr_n_T_295[18]), .Y(csr_n1855) );
  INVX1_LVT csr_U1981 ( .A(csr_n_T_295[17]), .Y(csr_n1854) );
  INVX1_LVT csr_U1980 ( .A(csr_n_T_295[16]), .Y(csr_n1853) );
  INVX1_LVT csr_U1979 ( .A(csr_n_T_295[15]), .Y(csr_n1852) );
  INVX1_LVT csr_U1978 ( .A(csr_n_T_295[14]), .Y(csr_n1851) );
  INVX1_LVT csr_U1977 ( .A(csr_n_T_295[13]), .Y(csr_n1850) );
  INVX1_LVT csr_U1976 ( .A(csr_n_T_295[11]), .Y(csr_n1849) );
  INVX1_LVT csr_U1975 ( .A(csr_n_T_295[9]), .Y(csr_n1848) );
  INVX1_LVT csr_U1974 ( .A(csr_n_T_286[7]), .Y(csr_n1847) );
  INVX1_LVT csr_U1973 ( .A(csr_n_T_286[6]), .Y(csr_n1846) );
  INVX1_LVT csr_U1972 ( .A(csr_n_T_286[5]), .Y(csr_n1845) );
  INVX1_LVT csr_U1971 ( .A(csr_n_T_286[3]), .Y(csr_n1844) );
  INVX1_LVT csr_U1970 ( .A(csr_n_T_286[2]), .Y(csr_n1843) );
  INVX1_LVT csr_U1969 ( .A(csr_n_T_286[1]), .Y(csr_n1842) );
  INVX1_LVT csr_U1968 ( .A(csr_n_T_286[29]), .Y(csr_n1841) );
  INVX1_LVT csr_U1967 ( .A(csr_n_T_286[28]), .Y(csr_n1840) );
  INVX1_LVT csr_U1966 ( .A(csr_n_T_286[27]), .Y(csr_n1839) );
  INVX1_LVT csr_U1965 ( .A(csr_n_T_286[26]), .Y(csr_n1838) );
  INVX1_LVT csr_U1964 ( .A(csr_n_T_286[25]), .Y(csr_n1837) );
  INVX1_LVT csr_U1963 ( .A(csr_n_T_286[24]), .Y(csr_n1836) );
  INVX1_LVT csr_U1962 ( .A(csr_n_T_286[23]), .Y(csr_n1835) );
  INVX1_LVT csr_U1961 ( .A(csr_n_T_286[22]), .Y(csr_n1834) );
  INVX1_LVT csr_U1960 ( .A(csr_n_T_286[21]), .Y(csr_n1833) );
  INVX1_LVT csr_U1959 ( .A(csr_n_T_286[20]), .Y(csr_n1832) );
  INVX1_LVT csr_U1958 ( .A(csr_n_T_286[19]), .Y(csr_n1831) );
  INVX1_LVT csr_U1957 ( .A(csr_n_T_286[18]), .Y(csr_n1830) );
  INVX1_LVT csr_U1956 ( .A(csr_n_T_286[17]), .Y(csr_n1829) );
  INVX1_LVT csr_U1955 ( .A(csr_n_T_286[16]), .Y(csr_n1828) );
  INVX1_LVT csr_U1954 ( .A(csr_n_T_286[15]), .Y(csr_n1827) );
  INVX1_LVT csr_U1953 ( .A(csr_n_T_286[14]), .Y(csr_n1826) );
  INVX1_LVT csr_U1952 ( .A(csr_n_T_286[13]), .Y(csr_n1825) );
  INVX1_LVT csr_U1951 ( .A(csr_n_T_286[11]), .Y(csr_n1824) );
  INVX1_LVT csr_U1950 ( .A(csr_n_T_286[9]), .Y(csr_n1823) );
  INVX1_LVT csr_U1949 ( .A(csr_n_T_277[7]), .Y(csr_n1822) );
  INVX1_LVT csr_U1948 ( .A(csr_n_T_277[6]), .Y(csr_n1821) );
  INVX1_LVT csr_U1947 ( .A(csr_n_T_277[5]), .Y(csr_n1820) );
  INVX1_LVT csr_U1946 ( .A(csr_n_T_277[3]), .Y(csr_n1819) );
  INVX1_LVT csr_U1945 ( .A(csr_n_T_277[2]), .Y(csr_n1818) );
  INVX1_LVT csr_U1944 ( .A(csr_n_T_277[1]), .Y(csr_n1817) );
  INVX1_LVT csr_U1943 ( .A(csr_n_T_277[29]), .Y(csr_n1816) );
  INVX1_LVT csr_U1942 ( .A(csr_n_T_277[28]), .Y(csr_n1815) );
  INVX1_LVT csr_U1941 ( .A(csr_n_T_277[27]), .Y(csr_n1814) );
  INVX1_LVT csr_U1940 ( .A(csr_n_T_277[26]), .Y(csr_n1813) );
  INVX1_LVT csr_U1939 ( .A(csr_n_T_277[25]), .Y(csr_n1812) );
  INVX1_LVT csr_U1938 ( .A(csr_n_T_277[24]), .Y(csr_n1811) );
  INVX1_LVT csr_U1937 ( .A(csr_n_T_277[23]), .Y(csr_n1810) );
  INVX1_LVT csr_U1936 ( .A(csr_n_T_277[22]), .Y(csr_n1809) );
  INVX1_LVT csr_U1935 ( .A(csr_n_T_277[21]), .Y(csr_n1808) );
  INVX1_LVT csr_U1934 ( .A(csr_n_T_277[20]), .Y(csr_n1807) );
  INVX1_LVT csr_U1933 ( .A(csr_n_T_277[19]), .Y(csr_n1806) );
  INVX1_LVT csr_U1932 ( .A(csr_n_T_277[18]), .Y(csr_n1805) );
  INVX1_LVT csr_U1931 ( .A(csr_n_T_277[17]), .Y(csr_n1804) );
  INVX1_LVT csr_U1930 ( .A(csr_n_T_277[16]), .Y(csr_n1803) );
  INVX1_LVT csr_U1929 ( .A(csr_n_T_277[15]), .Y(csr_n1802) );
  INVX1_LVT csr_U1928 ( .A(csr_n_T_277[14]), .Y(csr_n1801) );
  INVX1_LVT csr_U1927 ( .A(csr_n_T_277[13]), .Y(csr_n1800) );
  INVX1_LVT csr_U1926 ( .A(csr_n_T_277[11]), .Y(csr_n1799) );
  INVX1_LVT csr_U1925 ( .A(csr_n_T_277[9]), .Y(csr_n1798) );
  INVX1_LVT csr_U1924 ( .A(csr_n_T_268[7]), .Y(csr_n1797) );
  INVX1_LVT csr_U1923 ( .A(csr_n_T_268[6]), .Y(csr_n1796) );
  INVX1_LVT csr_U1922 ( .A(csr_n_T_268[5]), .Y(csr_n1795) );
  INVX1_LVT csr_U1921 ( .A(csr_n_T_268[3]), .Y(csr_n1794) );
  INVX1_LVT csr_U1920 ( .A(csr_n_T_268[2]), .Y(csr_n1793) );
  INVX1_LVT csr_U1919 ( .A(csr_n_T_268[1]), .Y(csr_n1792) );
  INVX1_LVT csr_U1918 ( .A(csr_n_T_268[29]), .Y(csr_n1791) );
  INVX1_LVT csr_U1917 ( .A(csr_n_T_268[28]), .Y(csr_n1790) );
  INVX1_LVT csr_U1916 ( .A(csr_n_T_268[27]), .Y(csr_n1789) );
  INVX1_LVT csr_U1915 ( .A(csr_n_T_268[26]), .Y(csr_n1788) );
  INVX1_LVT csr_U1914 ( .A(csr_n_T_268[25]), .Y(csr_n1787) );
  INVX1_LVT csr_U1913 ( .A(csr_n_T_268[24]), .Y(csr_n1786) );
  INVX1_LVT csr_U1912 ( .A(csr_n_T_268[23]), .Y(csr_n1785) );
  INVX1_LVT csr_U1911 ( .A(csr_n_T_268[22]), .Y(csr_n1784) );
  INVX1_LVT csr_U1910 ( .A(csr_n_T_268[21]), .Y(csr_n1783) );
  INVX1_LVT csr_U1909 ( .A(csr_n_T_268[20]), .Y(csr_n1782) );
  INVX1_LVT csr_U1908 ( .A(csr_n_T_268[19]), .Y(csr_n1781) );
  INVX1_LVT csr_U1907 ( .A(csr_n_T_268[18]), .Y(csr_n1780) );
  INVX1_LVT csr_U1906 ( .A(csr_n_T_268[17]), .Y(csr_n1779) );
  INVX1_LVT csr_U1905 ( .A(csr_n_T_268[16]), .Y(csr_n1778) );
  INVX1_LVT csr_U1904 ( .A(csr_n_T_268[15]), .Y(csr_n1777) );
  INVX1_LVT csr_U1903 ( .A(csr_n_T_268[14]), .Y(csr_n1776) );
  INVX1_LVT csr_U1902 ( .A(csr_n_T_268[13]), .Y(csr_n1775) );
  INVX1_LVT csr_U1901 ( .A(csr_n_T_268[11]), .Y(csr_n1774) );
  INVX1_LVT csr_U1900 ( .A(csr_n_T_268[9]), .Y(csr_n1773) );
  INVX1_LVT csr_U1899 ( .A(csr_n_T_259[7]), .Y(csr_n1772) );
  INVX1_LVT csr_U1898 ( .A(csr_n_T_259[6]), .Y(csr_n1771) );
  INVX1_LVT csr_U1897 ( .A(csr_n_T_259[5]), .Y(csr_n1770) );
  INVX1_LVT csr_U1896 ( .A(csr_n_T_259[3]), .Y(csr_n1769) );
  INVX1_LVT csr_U1895 ( .A(csr_n_T_259[2]), .Y(csr_n1768) );
  INVX1_LVT csr_U1894 ( .A(csr_n_T_259[1]), .Y(csr_n1767) );
  INVX1_LVT csr_U1893 ( .A(csr_n_T_259[29]), .Y(csr_n1766) );
  INVX1_LVT csr_U1892 ( .A(csr_n_T_259[28]), .Y(csr_n1765) );
  INVX1_LVT csr_U1891 ( .A(csr_n_T_259[27]), .Y(csr_n1764) );
  INVX1_LVT csr_U1890 ( .A(csr_n_T_259[26]), .Y(csr_n1763) );
  INVX1_LVT csr_U1889 ( .A(csr_n_T_259[25]), .Y(csr_n1762) );
  INVX1_LVT csr_U1888 ( .A(csr_n_T_259[24]), .Y(csr_n1761) );
  INVX1_LVT csr_U1887 ( .A(csr_n_T_259[23]), .Y(csr_n1760) );
  INVX1_LVT csr_U1886 ( .A(csr_n_T_259[22]), .Y(csr_n1759) );
  INVX1_LVT csr_U1885 ( .A(csr_n_T_259[21]), .Y(csr_n1758) );
  INVX1_LVT csr_U1884 ( .A(csr_n_T_259[20]), .Y(csr_n1757) );
  INVX1_LVT csr_U1883 ( .A(csr_n_T_259[19]), .Y(csr_n1756) );
  INVX1_LVT csr_U1882 ( .A(csr_n_T_259[18]), .Y(csr_n1755) );
  INVX1_LVT csr_U1881 ( .A(csr_n_T_259[17]), .Y(csr_n1754) );
  INVX1_LVT csr_U1880 ( .A(csr_n_T_259[16]), .Y(csr_n1753) );
  INVX1_LVT csr_U1879 ( .A(csr_n_T_259[15]), .Y(csr_n1752) );
  INVX1_LVT csr_U1878 ( .A(csr_n_T_259[14]), .Y(csr_n1751) );
  INVX1_LVT csr_U1877 ( .A(csr_n_T_259[13]), .Y(csr_n1750) );
  INVX1_LVT csr_U1876 ( .A(csr_n_T_259[11]), .Y(csr_n1749) );
  INVX1_LVT csr_U1875 ( .A(csr_n_T_259[9]), .Y(csr_n1748) );
  INVX1_LVT csr_U1874 ( .A(csr_n_T_250[7]), .Y(csr_n1747) );
  INVX1_LVT csr_U1873 ( .A(csr_n_T_250[6]), .Y(csr_n1746) );
  INVX1_LVT csr_U1872 ( .A(csr_n_T_250[5]), .Y(csr_n1745) );
  INVX1_LVT csr_U1871 ( .A(csr_n_T_250[3]), .Y(csr_n1744) );
  INVX1_LVT csr_U1870 ( .A(csr_n_T_250[2]), .Y(csr_n1743) );
  INVX1_LVT csr_U1869 ( .A(csr_n_T_250[1]), .Y(csr_n1742) );
  INVX1_LVT csr_U1868 ( .A(csr_n_T_250[29]), .Y(csr_n1741) );
  INVX1_LVT csr_U1867 ( .A(csr_n_T_250[28]), .Y(csr_n1740) );
  INVX1_LVT csr_U1866 ( .A(csr_n_T_250[27]), .Y(csr_n1739) );
  INVX1_LVT csr_U1865 ( .A(csr_n_T_250[26]), .Y(csr_n1738) );
  INVX1_LVT csr_U1864 ( .A(csr_n_T_250[25]), .Y(csr_n1737) );
  INVX1_LVT csr_U1863 ( .A(csr_n_T_250[24]), .Y(csr_n1736) );
  INVX1_LVT csr_U1862 ( .A(csr_n_T_250[23]), .Y(csr_n1735) );
  INVX1_LVT csr_U1861 ( .A(csr_n_T_250[22]), .Y(csr_n1734) );
  INVX1_LVT csr_U1860 ( .A(csr_n_T_250[21]), .Y(csr_n1733) );
  INVX1_LVT csr_U1859 ( .A(csr_n_T_250[20]), .Y(csr_n1732) );
  INVX1_LVT csr_U1858 ( .A(csr_n_T_250[19]), .Y(csr_n1731) );
  INVX1_LVT csr_U1857 ( .A(csr_n_T_250[18]), .Y(csr_n1730) );
  INVX1_LVT csr_U1856 ( .A(csr_n_T_250[17]), .Y(csr_n1729) );
  INVX1_LVT csr_U1855 ( .A(csr_n_T_250[16]), .Y(csr_n1728) );
  INVX1_LVT csr_U1854 ( .A(csr_n_T_250[15]), .Y(csr_n1727) );
  INVX1_LVT csr_U1853 ( .A(csr_n_T_250[14]), .Y(csr_n1726) );
  INVX1_LVT csr_U1852 ( .A(csr_n_T_250[13]), .Y(csr_n1725) );
  INVX1_LVT csr_U1851 ( .A(csr_n_T_250[11]), .Y(csr_n1724) );
  INVX1_LVT csr_U1850 ( .A(csr_n_T_250[9]), .Y(csr_n1723) );
  INVX1_LVT csr_U1849 ( .A(csr_n_T_241[7]), .Y(csr_n1722) );
  INVX1_LVT csr_U1848 ( .A(csr_n_T_241[6]), .Y(csr_n1721) );
  INVX1_LVT csr_U1847 ( .A(csr_n_T_241[5]), .Y(csr_n1720) );
  INVX1_LVT csr_U1846 ( .A(csr_n_T_241[3]), .Y(csr_n1719) );
  INVX1_LVT csr_U1845 ( .A(csr_n_T_241[2]), .Y(csr_n1718) );
  INVX1_LVT csr_U1844 ( .A(csr_n_T_241[1]), .Y(csr_n1717) );
  INVX1_LVT csr_U1843 ( .A(csr_n_T_241[29]), .Y(csr_n1716) );
  INVX1_LVT csr_U1842 ( .A(csr_n_T_241[28]), .Y(csr_n1715) );
  INVX1_LVT csr_U1841 ( .A(csr_n_T_241[27]), .Y(csr_n1714) );
  INVX1_LVT csr_U1840 ( .A(csr_n_T_241[26]), .Y(csr_n1713) );
  INVX1_LVT csr_U1839 ( .A(csr_n_T_241[25]), .Y(csr_n1712) );
  INVX1_LVT csr_U1838 ( .A(csr_n_T_241[24]), .Y(csr_n1711) );
  INVX1_LVT csr_U1837 ( .A(csr_n_T_241[23]), .Y(csr_n1710) );
  INVX1_LVT csr_U1836 ( .A(csr_n_T_241[22]), .Y(csr_n1709) );
  INVX1_LVT csr_U1835 ( .A(csr_n_T_241[21]), .Y(csr_n1708) );
  INVX1_LVT csr_U1834 ( .A(csr_n_T_241[20]), .Y(csr_n1707) );
  INVX1_LVT csr_U1833 ( .A(csr_n_T_241[19]), .Y(csr_n1706) );
  INVX1_LVT csr_U1832 ( .A(csr_n_T_241[18]), .Y(csr_n1705) );
  INVX1_LVT csr_U1831 ( .A(csr_n_T_241[17]), .Y(csr_n1704) );
  INVX1_LVT csr_U1830 ( .A(csr_n_T_241[16]), .Y(csr_n1703) );
  INVX1_LVT csr_U1829 ( .A(csr_n_T_241[15]), .Y(csr_n1702) );
  INVX1_LVT csr_U1828 ( .A(csr_n_T_241[14]), .Y(csr_n1701) );
  INVX1_LVT csr_U1827 ( .A(csr_n_T_241[13]), .Y(csr_n1700) );
  INVX1_LVT csr_U1826 ( .A(csr_n_T_241[11]), .Y(csr_n1699) );
  INVX1_LVT csr_U1825 ( .A(csr_n_T_241[9]), .Y(csr_n1698) );
  INVX1_LVT csr_U1824 ( .A(csr_n1553), .Y(csr_n1691) );
  MUX21X1_LVT csr_U1823 ( .A1(csr_io_pc[6]), .A2(csr_wdata_6_), .S0(csr_n514), 
        .Y(csr_net35064) );
  MUX21X1_LVT csr_U1822 ( .A1(csr_io_pc[6]), .A2(csr_wdata_6_), .S0(csr_n515), 
        .Y(csr_net35286) );
  MUX21X1_LVT csr_U1821 ( .A1(csr_io_pc[4]), .A2(csr_wdata_4_), .S0(csr_n513), 
        .Y(csr_net34868) );
  MUX21X1_LVT csr_U1820 ( .A1(csr_io_pc[4]), .A2(csr_wdata_4_), .S0(csr_n515), 
        .Y(csr_net35292) );
  MUX21X1_LVT csr_U1819 ( .A1(csr_io_pc[4]), .A2(csr_wdata_4_), .S0(csr_n514), 
        .Y(csr_net35070) );
  AO22X1_LVT csr_U1818 ( .A1(csr_n1481), .A2(csr_io_bp_0_control_x), .A3(
        csr_n1495), .A4(csr_n_T_389_2), .Y(csr_n1666) );
  AO22X1_LVT csr_U1817 ( .A1(csr_read_fcsr_2_), .A2(csr_n1167), .A3(csr_n1465), 
        .A4(csr_read_scounteren_2_), .Y(csr_n1663) );
  NAND2X0_LVT csr_U1816 ( .A1(csr_n1166), .A2(csr_n1165), .Y(csr_n_GEN_345[2])
         );
  NAND2X0_LVT csr_U1815 ( .A1(csr_n1164), .A2(io_fpu_fcsr_flags_bits[2]), .Y(
        csr_n1165) );
  MUX21X1_LVT csr_U1814 ( .A1(csr_n1483), .A2(csr_n477), .S0(csr_n1163), .Y(
        csr_n1166) );
  MUX21X1_LVT csr_U1813 ( .A1(csr_io_pc[2]), .A2(csr_wdata_2_), .S0(csr_n514), 
        .Y(csr_net35076) );
  MUX21X1_LVT csr_U1812 ( .A1(csr_io_pc[2]), .A2(csr_wdata_2_), .S0(csr_n513), 
        .Y(csr_net34874) );
  MUX21X1_LVT csr_U1811 ( .A1(csr_io_pc[39]), .A2(csr_wdata_39_), .S0(csr_n513), .Y(csr_net34763) );
  MUX21X1_LVT csr_U1810 ( .A1(csr_io_pc[39]), .A2(csr_wdata_39_), .S0(csr_n514), .Y(csr_net34965) );
  MUX21X1_LVT csr_U1809 ( .A1(csr_io_pc[37]), .A2(csr_wdata_37_), .S0(csr_n513), .Y(csr_net34769) );
  MUX21X1_LVT csr_U1808 ( .A1(csr_io_pc[37]), .A2(csr_wdata_37_), .S0(csr_n515), .Y(csr_net35193) );
  MUX21X1_LVT csr_U1807 ( .A1(csr_io_pc[37]), .A2(csr_wdata_37_), .S0(csr_n514), .Y(csr_net34971) );
  AO22X1_LVT csr_U1806 ( .A1(csr_n1689), .A2(csr_n_T_45_36_), .A3(csr_n1487), 
        .A4(csr_reg_stvec_36_), .Y(csr_n1640) );
  MUX21X1_LVT csr_U1805 ( .A1(csr_io_pc[36]), .A2(csr_wdata_36_), .S0(csr_n515), .Y(csr_net35196) );
  MUX21X1_LVT csr_U1804 ( .A1(csr_io_pc[36]), .A2(csr_wdata_36_), .S0(csr_n514), .Y(csr_net34974) );
  MUX21X1_LVT csr_U1803 ( .A1(csr_io_pc[35]), .A2(csr_wdata_35_), .S0(csr_n513), .Y(csr_net34775) );
  MUX21X1_LVT csr_U1802 ( .A1(csr_io_pc[34]), .A2(csr_wdata_34_), .S0(csr_n514), .Y(csr_net34980) );
  AO22X1_LVT csr_U1801 ( .A1(csr_n1162), .A2(csr_n1965), .A3(csr_n1487), .A4(
        csr_reg_stvec_34_), .Y(csr_n1635) );
  MUX21X1_LVT csr_U1800 ( .A1(csr_io_pc[34]), .A2(csr_wdata_34_), .S0(csr_n515), .Y(csr_net35202) );
  AO22X1_LVT csr_U1799 ( .A1(csr_n1162), .A2(csr_n1967), .A3(csr_n1487), .A4(
        csr_reg_stvec_32_), .Y(csr_n1630) );
  MUX21X1_LVT csr_U1798 ( .A1(csr_io_pc[32]), .A2(csr_wdata_32_), .S0(csr_n514), .Y(csr_net34986) );
  MUX21X1_LVT csr_U1797 ( .A1(csr_io_pc[31]), .A2(csr_wdata_31_), .S0(csr_n515), .Y(csr_net35211) );
  MUX21X1_LVT csr_U1796 ( .A1(csr_io_pc[31]), .A2(csr_wdata_31_), .S0(csr_n513), .Y(csr_net34787) );
  MUX21X1_LVT csr_U1795 ( .A1(csr_io_pc[31]), .A2(csr_wdata_31_), .S0(csr_n514), .Y(csr_net34989) );
  MUX21X1_LVT csr_U1794 ( .A1(csr_io_pc[30]), .A2(csr_wdata_30_), .S0(csr_n514), .Y(csr_net34992) );
  MUX21X1_LVT csr_U1793 ( .A1(csr_io_pc[29]), .A2(csr_wdata_29_), .S0(csr_n513), .Y(csr_net34793) );
  MUX21X1_LVT csr_U1792 ( .A1(csr_io_pc[28]), .A2(csr_wdata_28_), .S0(csr_n513), .Y(csr_net34796) );
  MUX21X1_LVT csr_U1791 ( .A1(csr_io_pc[28]), .A2(csr_wdata_28_), .S0(csr_n514), .Y(csr_net34998) );
  MUX21X1_LVT csr_U1790 ( .A1(csr_io_pc[27]), .A2(csr_wdata_27_), .S0(csr_n513), .Y(csr_net34799) );
  MUX21X1_LVT csr_U1789 ( .A1(csr_io_pc[27]), .A2(csr_wdata_27_), .S0(csr_n514), .Y(csr_net35001) );
  MUX21X1_LVT csr_U1788 ( .A1(csr_io_pc[26]), .A2(csr_wdata_26_), .S0(csr_n515), .Y(csr_net35226) );
  MUX21X1_LVT csr_U1787 ( .A1(csr_io_pc[26]), .A2(csr_wdata_26_), .S0(csr_n513), .Y(csr_net34802) );
  MUX21X1_LVT csr_U1786 ( .A1(csr_io_pc[25]), .A2(csr_wdata_25_), .S0(csr_n515), .Y(csr_net35229) );
  MUX21X1_LVT csr_U1785 ( .A1(csr_io_pc[25]), .A2(csr_wdata_25_), .S0(csr_n514), .Y(csr_net35007) );
  MUX21X1_LVT csr_U1784 ( .A1(csr_io_pc[24]), .A2(csr_wdata_24_), .S0(csr_n514), .Y(csr_net35010) );
  MUX21X1_LVT csr_U1783 ( .A1(csr_io_pc[24]), .A2(csr_wdata_24_), .S0(csr_n513), .Y(csr_net34808) );
  AO22X1_LVT csr_U1782 ( .A1(csr_n1160), .A2(csr_n_T_444[23]), .A3(csr_n1506), 
        .A4(csr_reg_sepc_23_), .Y(csr_n1603) );
  MUX21X1_LVT csr_U1781 ( .A1(csr_io_pc[23]), .A2(csr_wdata_23_), .S0(csr_n513), .Y(csr_net34811) );
  AO22X1_LVT csr_U1780 ( .A1(csr_n1159), .A2(csr_io_tval[23]), .A3(
        csr_wdata_23_), .A4(csr_n1158), .Y(csr_N1405) );
  MUX21X1_LVT csr_U1779 ( .A1(csr_io_pc[23]), .A2(csr_wdata_23_), .S0(csr_n515), .Y(csr_net35235) );
  MUX21X1_LVT csr_U1778 ( .A1(csr_io_pc[22]), .A2(csr_wdata_22_), .S0(csr_n514), .Y(csr_net35016) );
  MUX21X1_LVT csr_U1777 ( .A1(csr_io_pc[22]), .A2(csr_wdata_22_), .S0(csr_n513), .Y(csr_net34814) );
  MUX21X1_LVT csr_U1776 ( .A1(csr_io_pc[21]), .A2(csr_wdata_21_), .S0(csr_n513), .Y(csr_net34817) );
  MUX21X1_LVT csr_U1775 ( .A1(csr_io_pc[21]), .A2(csr_wdata_21_), .S0(csr_n515), .Y(csr_net35241) );
  AO22X1_LVT csr_U1774 ( .A1(csr_n1689), .A2(csr_n_T_45_20_), .A3(csr_n1487), 
        .A4(csr_reg_stvec_20_), .Y(csr_n1596) );
  AO22X1_LVT csr_U1773 ( .A1(csr_n1689), .A2(csr_n_T_45_19_), .A3(csr_n1487), 
        .A4(csr_reg_stvec_19_), .Y(csr_n1591) );
  MUX21X1_LVT csr_U1772 ( .A1(csr_io_pc[19]), .A2(csr_wdata_19_), .S0(csr_n515), .Y(csr_net35247) );
  MUX21X1_LVT csr_U1771 ( .A1(csr_io_pc[19]), .A2(csr_wdata_19_), .S0(csr_n513), .Y(csr_net34823) );
  MUX21X1_LVT csr_U1770 ( .A1(csr_io_pc[19]), .A2(csr_wdata_19_), .S0(csr_n514), .Y(csr_net35025) );
  MUX21X1_LVT csr_U1769 ( .A1(csr_io_pc[18]), .A2(csr_wdata_18_), .S0(csr_n515), .Y(csr_net35250) );
  MUX21X1_LVT csr_U1768 ( .A1(csr_io_pc[18]), .A2(csr_wdata_18_), .S0(csr_n514), .Y(csr_net35028) );
  MUX21X1_LVT csr_U1767 ( .A1(csr_io_pc[18]), .A2(csr_wdata_18_), .S0(csr_n513), .Y(csr_net34826) );
  AO22X1_LVT csr_U1766 ( .A1(csr_n1159), .A2(csr_io_tval[17]), .A3(
        csr_wdata_17_), .A4(csr_n1158), .Y(csr_N1399) );
  MUX21X1_LVT csr_U1765 ( .A1(csr_io_pc[17]), .A2(csr_wdata_17_), .S0(csr_n515), .Y(csr_net35253) );
  MUX21X1_LVT csr_U1764 ( .A1(csr_io_pc[17]), .A2(csr_wdata_17_), .S0(csr_n513), .Y(csr_net34829) );
  AO22X1_LVT csr_U1763 ( .A1(csr_n1157), .A2(csr_n1927), .A3(csr_n1480), .A4(
        io_ptw_pmp_0_addr[17]), .Y(csr_n1573) );
  MUX21X1_LVT csr_U1762 ( .A1(csr_io_pc[16]), .A2(csr_wdata_16_), .S0(csr_n513), .Y(csr_net34832) );
  MUX21X1_LVT csr_U1761 ( .A1(csr_io_pc[16]), .A2(csr_wdata_16_), .S0(csr_n514), .Y(csr_net35034) );
  MUX21X1_LVT csr_U1760 ( .A1(csr_io_pc[15]), .A2(csr_wdata_15_), .S0(csr_n513), .Y(csr_net34835) );
  MUX21X1_LVT csr_U1759 ( .A1(csr_io_pc[14]), .A2(csr_wdata_14_), .S0(csr_n513), .Y(csr_net34838) );
  MUX21X1_LVT csr_U1758 ( .A1(csr_io_pc[14]), .A2(csr_wdata_14_), .S0(csr_n515), .Y(csr_net35262) );
  MUX21X1_LVT csr_U1757 ( .A1(csr_io_pc[13]), .A2(csr_wdata_13_), .S0(csr_n514), .Y(csr_net35043) );
  MUX21X1_LVT csr_U1756 ( .A1(csr_io_pc[13]), .A2(csr_wdata_13_), .S0(csr_n513), .Y(csr_net34841) );
  MUX21X1_LVT csr_U1755 ( .A1(csr_io_pc[13]), .A2(csr_wdata_13_), .S0(csr_n515), .Y(csr_net35265) );
  MUX21X1_LVT csr_U1754 ( .A1(csr_io_pc[12]), .A2(csr_wdata_12_), .S0(csr_n513), .Y(csr_net34844) );
  MUX21X1_LVT csr_U1753 ( .A1(csr_io_pc[12]), .A2(csr_wdata_12_), .S0(csr_n514), .Y(csr_net35046) );
  MUX21X1_LVT csr_U1752 ( .A1(csr_io_pc[12]), .A2(csr_wdata_12_), .S0(csr_n515), .Y(csr_net35268) );
  MUX21X1_LVT csr_U1751 ( .A1(csr_io_pc[10]), .A2(csr_wdata_10_), .S0(csr_n513), .Y(csr_net34850) );
  MUX21X1_LVT csr_U1750 ( .A1(csr_io_pc[10]), .A2(csr_wdata_10_), .S0(csr_n515), .Y(csr_net35274) );
  AO22X1_LVT csr_U1749 ( .A1(csr_n1154), .A2(csr_n1933), .A3(csr_n1480), .A4(
        io_ptw_pmp_0_addr[5]), .Y(csr_n1541) );
  AO22X1_LVT csr_U1748 ( .A1(csr_n1152), .A2(csr_io_tval[5]), .A3(csr_wdata_5_), .A4(csr_n1151), .Y(csr_N998) );
  MUX21X1_LVT csr_U1747 ( .A1(csr_io_pc[5]), .A2(csr_wdata_5_), .S0(csr_n515), 
        .Y(csr_net35289) );
  AO22X1_LVT csr_U1746 ( .A1(csr_io_tval[5]), .A2(csr_n1159), .A3(csr_wdata_5_), .A4(csr_n1158), .Y(csr_N1387) );
  MUX21X1_LVT csr_U1745 ( .A1(csr_io_pc[5]), .A2(csr_wdata_5_), .S0(csr_n514), 
        .Y(csr_net35067) );
  MUX21X1_LVT csr_U1744 ( .A1(csr_io_pc[5]), .A2(csr_wdata_5_), .S0(csr_n513), 
        .Y(csr_net34865) );
  MUX21X1_LVT csr_U1743 ( .A1(csr_io_pc[8]), .A2(csr_wdata_8_), .S0(csr_n515), 
        .Y(csr_net35280) );
  MUX21X1_LVT csr_U1742 ( .A1(csr_io_pc[8]), .A2(csr_wdata_8_), .S0(csr_n514), 
        .Y(csr_net35058) );
  MUX21X1_LVT csr_U1741 ( .A1(csr_io_pc[8]), .A2(csr_wdata_8_), .S0(csr_n513), 
        .Y(csr_net34856) );
  AO21X1_LVT csr_U1740 ( .A1(csr_n1922), .A2(csr_n504), .A3(csr_n376), .Y(
        csr_N1567) );
  AO22X1_LVT csr_U1739 ( .A1(csr_n1159), .A2(csr_io_tval[8]), .A3(csr_wdata_8_), .A4(csr_n1158), .Y(csr_N1390) );
  AO22X1_LVT csr_U1738 ( .A1(csr_n1152), .A2(csr_io_tval[8]), .A3(csr_wdata_8_), .A4(csr_n1151), .Y(csr_N1001) );
  AO22X1_LVT csr_U1737 ( .A1(csr_n1150), .A2(csr_n_T_52[2]), .A3(csr_wdata_8_), 
        .A4(csr_n1149), .Y(csr_N1893) );
  AO22X1_LVT csr_U1736 ( .A1(csr_n498), .A2(csr_n_T_52[26]), .A3(csr_wdata_32_), .A4(csr_n1149), .Y(csr_N1917) );
  AO22X1_LVT csr_U1735 ( .A1(csr_n498), .A2(csr_n_T_52[28]), .A3(csr_wdata_34_), .A4(csr_n1149), .Y(csr_N1919) );
  AO22X1_LVT csr_U1734 ( .A1(csr_n1149), .A2(csr_wdata_63_), .A3(
        csr_n_T_52[57]), .A4(csr_n496), .Y(csr_N1948) );
  AO22X1_LVT csr_U1733 ( .A1(csr_n1446), .A2(csr_n1148), .A3(csr_wdata_5_), 
        .A4(csr_n1149), .Y(csr_N1827) );
  AO22X1_LVT csr_U1732 ( .A1(csr_n1446), .A2(csr_n1146), .A3(csr_wdata_4_), 
        .A4(csr_n1149), .Y(csr_N1826) );
  AOI21X1_LVT csr_U1731 ( .A1(csr_n1145), .A2(csr_n454), .A3(csr_n1147), .Y(
        csr_n1146) );
  NAND2X0_LVT csr_U1730 ( .A1(csr_n1144), .A2(csr_io_time[3]), .Y(csr_n1145)
         );
  AO22X1_LVT csr_U1729 ( .A1(csr_n1446), .A2(csr_n1143), .A3(csr_wdata_2_), 
        .A4(csr_n1149), .Y(csr_N1824) );
  OA21X1_LVT csr_U1728 ( .A1(csr_n1142), .A2(csr_io_time[2]), .A3(csr_n1141), 
        .Y(csr_n1143) );
  NAND4X0_LVT csr_U1727 ( .A1(csr_n1138), .A2(csr_n1183), .A3(csr_n1182), .A4(
        csr_n1137), .Y(csr_n1140) );
  AND4X1_LVT csr_U1726 ( .A1(csr_n1179), .A2(csr_n1172), .A3(csr_n590), .A4(
        csr_n1186), .Y(csr_n1137) );
  NAND2X0_LVT csr_U1725 ( .A1(csr_reg_mie_7_), .A2(io_interrupts_mtip), .Y(
        csr_n1172) );
  NAND2X0_LVT csr_U1724 ( .A1(csr_n_T_61_5_), .A2(csr_reg_mie_5_), .Y(
        csr_n1179) );
  AND2X1_LVT csr_U1723 ( .A1(csr_n1171), .A2(csr_n1178), .Y(csr_n1182) );
  NAND2X0_LVT csr_U1722 ( .A1(csr_n_T_61_1), .A2(csr_reg_mie_1_), .Y(csr_n1178) );
  NAND2X0_LVT csr_U1721 ( .A1(csr_n1136), .A2(csr_reg_mie_9_), .Y(csr_n1171)
         );
  AND2X1_LVT csr_U1720 ( .A1(csr_n1188), .A2(csr_n1193), .Y(csr_n1183) );
  NAND2X0_LVT csr_U1719 ( .A1(csr_reg_mie_3_), .A2(io_interrupts_msip), .Y(
        csr_n1193) );
  NAND2X0_LVT csr_U1718 ( .A1(csr_reg_mie_11_), .A2(io_interrupts_meip), .Y(
        csr_n1188) );
  NAND2X0_LVT csr_U1717 ( .A1(csr_n1135), .A2(csr_n472), .Y(csr_n1138) );
  NAND4X0_LVT csr_U1716 ( .A1(csr_n1134), .A2(csr_n1133), .A3(csr_n1519), .A4(
        csr_n1517), .Y(csr_n1135) );
  NOR3X0_LVT csr_U1715 ( .A1(csr_io_status_debug), .A2(csr_n_T_389_2), .A3(
        csr_io_rw_addr[9]), .Y(csr_n1133) );
  AO22X1_LVT csr_U1714 ( .A1(csr_n1695), .A2(csr_n1504), .A3(csr_n427), .A4(
        csr_n1132), .Y(csr_N611) );
  INVX1_LVT csr_U1713 ( .A(csr_n1694), .Y(csr_n1132) );
  AO22X1_LVT csr_U1712 ( .A1(csr_n1474), .A2(csr_n1131), .A3(csr_n_T_61_5_), 
        .A4(csr_n1906), .Y(csr_n199) );
  AND2X1_LVT csr_U1711 ( .A1(io_imem_sfence_bits_addr[5]), .A2(csr_n516), .Y(
        csr_n1131) );
  AO222X1_LVT csr_U1710 ( .A1(csr_wdata_1_), .A2(csr_n1901), .A3(csr_n1902), 
        .A4(csr_n_T_61_1), .A5(csr_n1474), .A6(csr_n1900), .Y(csr_n2162) );
  AO22X1_LVT csr_U1709 ( .A1(csr_n1693), .A2(csr_n1504), .A3(csr_n407), .A4(
        csr_n1130), .Y(csr_N607) );
  INVX1_LVT csr_U1708 ( .A(csr_n1692), .Y(csr_n1130) );
  AO22X1_LVT csr_U1707 ( .A1(csr_reg_mie_11_), .A2(csr_n1503), .A3(
        csr_wdata_11_), .A4(csr_n1502), .Y(csr_N617) );
  MUX21X1_LVT csr_U1706 ( .A1(csr_io_pc[11]), .A2(csr_wdata_11_), .S0(csr_n514), .Y(csr_net35049) );
  MUX21X1_LVT csr_U1705 ( .A1(io_ptw_pmp_7_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n512), .Y(csr_n_GEN_307[11]) );
  MUX21X1_LVT csr_U1704 ( .A1(io_ptw_pmp_0_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n505), .Y(csr_n_GEN_258[11]) );
  MUX21X1_LVT csr_U1703 ( .A1(io_ptw_pmp_4_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n509), .Y(csr_n_GEN_286[11]) );
  MUX21X1_LVT csr_U1702 ( .A1(io_ptw_pmp_5_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n510), .Y(csr_n_GEN_293[11]) );
  MUX21X1_LVT csr_U1701 ( .A1(io_ptw_pmp_3_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n508), .Y(csr_n_GEN_279[11]) );
  MUX21X1_LVT csr_U1700 ( .A1(io_ptw_pmp_2_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n507), .Y(csr_n_GEN_272[11]) );
  MUX21X1_LVT csr_U1699 ( .A1(io_ptw_pmp_6_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n511), .Y(csr_n_GEN_300[11]) );
  MUX21X1_LVT csr_U1698 ( .A1(io_ptw_pmp_1_addr[11]), .A2(csr_wdata_11_), .S0(
        csr_n506), .Y(csr_n_GEN_265[11]) );
  AO22X1_LVT csr_U1697 ( .A1(csr_n493), .A2(csr_n_T_44[9]), .A3(csr_wdata_15_), 
        .A4(csr_n1128), .Y(csr_N1506) );
  AO22X1_LVT csr_U1696 ( .A1(csr_n493), .A2(csr_n_T_44[2]), .A3(csr_wdata_8_), 
        .A4(csr_n1128), .Y(csr_N1499) );
  AO22X1_LVT csr_U1695 ( .A1(csr_n493), .A2(csr_n_T_44[4]), .A3(csr_wdata_10_), 
        .A4(csr_n491), .Y(csr_N1501) );
  MUX21X1_LVT csr_U1694 ( .A1(csr_io_pc[10]), .A2(csr_wdata_10_), .S0(csr_n514), .Y(csr_net35052) );
  AO22X1_LVT csr_U1693 ( .A1(csr_n1159), .A2(csr_io_tval[10]), .A3(
        csr_wdata_10_), .A4(csr_n1158), .Y(csr_N1392) );
  AO22X1_LVT csr_U1692 ( .A1(csr_n1152), .A2(csr_io_tval[10]), .A3(
        csr_wdata_10_), .A4(csr_n1151), .Y(csr_N1003) );
  AO22X1_LVT csr_U1691 ( .A1(csr_n498), .A2(csr_n_T_52[4]), .A3(csr_wdata_10_), 
        .A4(csr_n1149), .Y(csr_N1895) );
  AO22X1_LVT csr_U1690 ( .A1(csr_n494), .A2(csr_n_T_44[5]), .A3(csr_wdata_11_), 
        .A4(csr_n491), .Y(csr_N1502) );
  AO22X1_LVT csr_U1689 ( .A1(csr_n493), .A2(csr_n_T_44[10]), .A3(csr_wdata_16_), .A4(csr_n492), .Y(csr_N1507) );
  MUX21X1_LVT csr_U1688 ( .A1(csr_io_pc[16]), .A2(csr_wdata_16_), .S0(csr_n515), .Y(csr_net35256) );
  AO22X1_LVT csr_U1687 ( .A1(csr_n1159), .A2(csr_io_tval[16]), .A3(
        csr_wdata_16_), .A4(csr_n1158), .Y(csr_N1398) );
  AO22X1_LVT csr_U1686 ( .A1(csr_n1152), .A2(csr_io_tval[16]), .A3(
        csr_wdata_16_), .A4(csr_n1151), .Y(csr_N1009) );
  AO22X1_LVT csr_U1685 ( .A1(csr_n498), .A2(csr_n_T_52[10]), .A3(csr_wdata_16_), .A4(csr_n1149), .Y(csr_N1901) );
  NAND2X0_LVT csr_U1684 ( .A1(csr_n1127), .A2(csr_n1570), .Y(
        csr_io_rw_rdata[16]) );
  NOR4X1_LVT csr_U1683 ( .A1(csr_n1562), .A2(csr_n1561), .A3(csr_n1126), .A4(
        csr_n1569), .Y(csr_n1127) );
  OR2X1_LVT csr_U1682 ( .A1(csr_n1125), .A2(csr_n1563), .Y(csr_n1126) );
  NAND4X0_LVT csr_U1681 ( .A1(csr_n1124), .A2(csr_n1123), .A3(csr_n1122), .A4(
        csr_n1121), .Y(csr_n1125) );
  NAND2X0_LVT csr_U1680 ( .A1(csr_n1153), .A2(csr_n_T_383[16]), .Y(csr_n1121)
         );
  AOI21X1_LVT csr_U1679 ( .A1(csr_n1493), .A2(csr_reg_dpc_16_), .A3(csr_n1120), 
        .Y(csr_n1122) );
  AO22X1_LVT csr_U1678 ( .A1(csr_n1689), .A2(csr_n_T_45_16_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[16]), .Y(csr_n1120) );
  AO22X1_LVT csr_U1677 ( .A1(csr_n493), .A2(csr_n_T_44[11]), .A3(csr_wdata_17_), .A4(csr_n1128), .Y(csr_N1508) );
  MUX21X1_LVT csr_U1676 ( .A1(csr_io_pc[17]), .A2(csr_wdata_17_), .S0(csr_n514), .Y(csr_net35031) );
  AO22X1_LVT csr_U1675 ( .A1(csr_n1152), .A2(csr_io_tval[17]), .A3(
        csr_wdata_17_), .A4(csr_n1151), .Y(csr_N1010) );
  AO22X1_LVT csr_U1674 ( .A1(csr_n498), .A2(csr_n_T_52[11]), .A3(csr_wdata_17_), .A4(csr_n1149), .Y(csr_N1902) );
  NAND3X0_LVT csr_U1673 ( .A1(csr_n1580), .A2(csr_n1581), .A3(csr_n1119), .Y(
        csr_io_rw_rdata[17]) );
  NOR4X1_LVT csr_U1672 ( .A1(csr_n1118), .A2(csr_n1117), .A3(csr_n1116), .A4(
        csr_n1115), .Y(csr_n1119) );
  AO22X1_LVT csr_U1671 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[17]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[17]), .Y(csr_n1115) );
  AO22X1_LVT csr_U1670 ( .A1(csr_n1489), .A2(csr_reg_mepc_17_), .A3(csr_n1162), 
        .A4(csr_io_time[17]), .Y(csr_n1116) );
  AND2X1_LVT csr_U1669 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[17]), .Y(
        csr_n1117) );
  AO21X1_LVT csr_U1668 ( .A1(csr_n1153), .A2(csr_n_T_383[17]), .A3(csr_n1114), 
        .Y(csr_n1118) );
  NAND4X0_LVT csr_U1667 ( .A1(csr_n1113), .A2(csr_n1579), .A3(csr_n1112), .A4(
        csr_n1111), .Y(csr_n1114) );
  NAND2X0_LVT csr_U1666 ( .A1(csr_n1689), .A2(csr_n_T_45_17_), .Y(csr_n1111)
         );
  NAND2X0_LVT csr_U1665 ( .A1(csr_n1488), .A2(io_ptw_ptbr_ppn[17]), .Y(
        csr_n1112) );
  NAND2X0_LVT csr_U1664 ( .A1(io_ptw_pmp_2_cfg_w), .A2(csr_n1507), .Y(
        csr_n1113) );
  AO22X1_LVT csr_U1663 ( .A1(csr_n493), .A2(csr_n_T_44[12]), .A3(csr_wdata_18_), .A4(csr_n492), .Y(csr_N1509) );
  AO21X1_LVT csr_U1662 ( .A1(csr_n1921), .A2(csr_n504), .A3(csr_n376), .Y(
        csr_N1577) );
  AO22X1_LVT csr_U1661 ( .A1(csr_n1159), .A2(csr_io_tval[18]), .A3(
        csr_wdata_18_), .A4(csr_n1158), .Y(csr_N1400) );
  AO22X1_LVT csr_U1660 ( .A1(csr_n1152), .A2(csr_io_tval[18]), .A3(
        csr_wdata_18_), .A4(csr_n1151), .Y(csr_N1011) );
  AO22X1_LVT csr_U1659 ( .A1(csr_n498), .A2(csr_n_T_52[12]), .A3(csr_wdata_18_), .A4(csr_n1149), .Y(csr_N1903) );
  NAND4X0_LVT csr_U1658 ( .A1(csr_n1110), .A2(csr_n1109), .A3(csr_n1108), .A4(
        csr_n1107), .Y(csr_io_rw_rdata[18]) );
  NOR4X1_LVT csr_U1657 ( .A1(csr_n1106), .A2(csr_n1105), .A3(csr_n1104), .A4(
        csr_n1103), .Y(csr_n1108) );
  AO22X1_LVT csr_U1656 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[18]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[18]), .Y(csr_n1103) );
  AO22X1_LVT csr_U1655 ( .A1(csr_n1162), .A2(csr_io_time[18]), .A3(csr_n1480), 
        .A4(io_ptw_pmp_0_addr[18]), .Y(csr_n1104) );
  NOR4X1_LVT csr_U1654 ( .A1(csr_n1102), .A2(csr_n1101), .A3(csr_n1100), .A4(
        csr_n1582), .Y(csr_n1110) );
  AO22X1_LVT csr_U1653 ( .A1(csr_n1153), .A2(csr_n_T_383[18]), .A3(csr_n1452), 
        .A4(csr_n1921), .Y(csr_n1100) );
  NAND4X0_LVT csr_U1652 ( .A1(csr_n1099), .A2(csr_n1098), .A3(csr_n1097), .A4(
        csr_n1096), .Y(csr_n1101) );
  NAND2X0_LVT csr_U1651 ( .A1(io_ptw_pmp_2_cfg_x), .A2(csr_n1507), .Y(
        csr_n1096) );
  AOI22X1_LVT csr_U1650 ( .A1(csr_n1689), .A2(csr_n_T_45_18_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[18]), .Y(csr_n1097) );
  NAND2X0_LVT csr_U1649 ( .A1(io_ptw_status_sum), .A2(csr_n1154), .Y(csr_n1098) );
  NAND2X0_LVT csr_U1648 ( .A1(csr_reg_stvec_18_), .A2(csr_n1487), .Y(csr_n1099) );
  AO22X1_LVT csr_U1647 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[18]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[18]), .Y(csr_n1102) );
  AO22X1_LVT csr_U1646 ( .A1(csr_n493), .A2(csr_n_T_44[13]), .A3(csr_wdata_19_), .A4(csr_n1128), .Y(csr_N1510) );
  AO22X1_LVT csr_U1645 ( .A1(csr_n1159), .A2(csr_io_tval[19]), .A3(
        csr_wdata_19_), .A4(csr_n1158), .Y(csr_N1401) );
  AO22X1_LVT csr_U1644 ( .A1(csr_n1152), .A2(csr_io_tval[19]), .A3(
        csr_wdata_19_), .A4(csr_n1151), .Y(csr_N1012) );
  AO22X1_LVT csr_U1643 ( .A1(csr_n498), .A2(csr_n_T_52[13]), .A3(csr_wdata_19_), .A4(csr_n1149), .Y(csr_N1904) );
  NAND3X0_LVT csr_U1642 ( .A1(csr_n1095), .A2(csr_n1094), .A3(csr_n1093), .Y(
        csr_io_rw_rdata[19]) );
  NOR4X1_LVT csr_U1641 ( .A1(csr_n1092), .A2(csr_n1091), .A3(csr_n1090), .A4(
        csr_n1089), .Y(csr_n1093) );
  NAND4X0_LVT csr_U1640 ( .A1(csr_n1088), .A2(csr_n1087), .A3(csr_n1086), .A4(
        csr_n1085), .Y(csr_n1089) );
  NAND2X0_LVT csr_U1639 ( .A1(io_ptw_status_mxr), .A2(csr_n1154), .Y(csr_n1085) );
  NAND2X0_LVT csr_U1638 ( .A1(csr_n_T_383[19]), .A2(csr_n1153), .Y(csr_n1086)
         );
  AND4X1_LVT csr_U1637 ( .A1(csr_n1084), .A2(csr_n1083), .A3(csr_n1082), .A4(
        csr_n478), .Y(csr_n1087) );
  NAND2X0_LVT csr_U1636 ( .A1(csr_n488), .A2(io_ptw_ptbr_ppn[19]), .Y(
        csr_n1082) );
  NAND2X0_LVT csr_U1635 ( .A1(io_ptw_pmp_2_cfg_a[0]), .A2(csr_n1507), .Y(
        csr_n1084) );
  NAND2X0_LVT csr_U1634 ( .A1(io_ptw_pmp_6_addr[19]), .A2(csr_n1494), .Y(
        csr_n1088) );
  AO22X1_LVT csr_U1633 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[19]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[19]), .Y(csr_n1090) );
  AO22X1_LVT csr_U1632 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[19]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[19]), .Y(csr_n1091) );
  NOR4X1_LVT csr_U1631 ( .A1(csr_n1587), .A2(csr_n1081), .A3(csr_n1080), .A4(
        csr_n1588), .Y(csr_n1095) );
  AO22X1_LVT csr_U1630 ( .A1(csr_n1160), .A2(csr_n_T_444[19]), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_19_), .Y(csr_n1080) );
  AO22X1_LVT csr_U1629 ( .A1(csr_n493), .A2(csr_n_T_44[14]), .A3(csr_wdata_20_), .A4(csr_n491), .Y(csr_N1511) );
  MUX21X1_LVT csr_U1628 ( .A1(csr_io_pc[20]), .A2(csr_wdata_20_), .S0(csr_n514), .Y(csr_net35022) );
  MUX21X1_LVT csr_U1627 ( .A1(csr_io_pc[20]), .A2(csr_wdata_20_), .S0(csr_n515), .Y(csr_net35244) );
  MUX21X1_LVT csr_U1626 ( .A1(csr_io_pc[20]), .A2(csr_wdata_20_), .S0(csr_n513), .Y(csr_net34820) );
  AO21X1_LVT csr_U1625 ( .A1(csr_n1920), .A2(csr_n504), .A3(csr_n376), .Y(
        csr_N1579) );
  AO22X1_LVT csr_U1624 ( .A1(csr_n1159), .A2(csr_io_tval[20]), .A3(
        csr_wdata_20_), .A4(csr_n1158), .Y(csr_N1402) );
  AO22X1_LVT csr_U1623 ( .A1(csr_n1152), .A2(csr_io_tval[20]), .A3(
        csr_wdata_20_), .A4(csr_n1151), .Y(csr_N1013) );
  AO22X1_LVT csr_U1622 ( .A1(csr_n496), .A2(csr_n_T_52[14]), .A3(csr_wdata_20_), .A4(csr_n1149), .Y(csr_N1905) );
  NAND2X0_LVT csr_U1621 ( .A1(csr_n1079), .A2(csr_n1078), .Y(
        csr_io_rw_rdata[20]) );
  NOR3X0_LVT csr_U1620 ( .A1(csr_n1594), .A2(csr_n1597), .A3(csr_n1593), .Y(
        csr_n1078) );
  NOR4X1_LVT csr_U1619 ( .A1(csr_n1077), .A2(csr_n1076), .A3(csr_n1592), .A4(
        csr_n1595), .Y(csr_n1079) );
  NAND4X0_LVT csr_U1618 ( .A1(csr_n1075), .A2(csr_n1074), .A3(csr_n1073), .A4(
        csr_n1072), .Y(csr_n1076) );
  AOI22X1_LVT csr_U1617 ( .A1(csr_n1160), .A2(csr_n_T_444[20]), .A3(csr_n1489), 
        .A4(csr_reg_mepc_20_), .Y(csr_n1074) );
  AOI22X1_LVT csr_U1616 ( .A1(csr_n1485), .A2(csr_reg_mscratch[20]), .A3(
        csr_n1157), .A4(csr_n1926), .Y(csr_n1075) );
  NAND4X0_LVT csr_U1615 ( .A1(csr_n1071), .A2(csr_n1070), .A3(csr_n1069), .A4(
        csr_n1068), .Y(csr_n1077) );
  NAND2X0_LVT csr_U1614 ( .A1(io_ptw_pmp_2_addr[20]), .A2(csr_n1492), .Y(
        csr_n1068) );
  NAND2X0_LVT csr_U1613 ( .A1(csr_n1920), .A2(csr_n1452), .Y(csr_n1069) );
  AND4X1_LVT csr_U1612 ( .A1(csr_n1067), .A2(csr_n1083), .A3(csr_n1066), .A4(
        csr_n1065), .Y(csr_n1070) );
  NAND2X0_LVT csr_U1611 ( .A1(csr_n1510), .A2(csr_reg_dscratch[20]), .Y(
        csr_n1065) );
  NAND2X0_LVT csr_U1610 ( .A1(csr_n1493), .A2(csr_reg_dpc_20_), .Y(csr_n1066)
         );
  NAND2X0_LVT csr_U1609 ( .A1(io_ptw_pmp_2_cfg_a[1]), .A2(csr_n1507), .Y(
        csr_n1067) );
  AOI22X1_LVT csr_U1608 ( .A1(csr_n1162), .A2(csr_io_time[20]), .A3(csr_n1506), 
        .A4(csr_reg_sepc_20_), .Y(csr_n1071) );
  AO22X1_LVT csr_U1607 ( .A1(csr_n493), .A2(csr_n_T_44[15]), .A3(csr_wdata_21_), .A4(csr_n1128), .Y(csr_N1512) );
  MUX21X1_LVT csr_U1606 ( .A1(csr_io_pc[21]), .A2(csr_wdata_21_), .S0(csr_n514), .Y(csr_net35019) );
  AO22X1_LVT csr_U1605 ( .A1(csr_n1159), .A2(csr_io_tval[21]), .A3(
        csr_wdata_21_), .A4(csr_n1158), .Y(csr_N1403) );
  AO22X1_LVT csr_U1604 ( .A1(csr_n1152), .A2(csr_io_tval[21]), .A3(
        csr_wdata_21_), .A4(csr_n1151), .Y(csr_N1014) );
  AO22X1_LVT csr_U1603 ( .A1(csr_n497), .A2(csr_n_T_52[15]), .A3(csr_wdata_21_), .A4(csr_n1149), .Y(csr_N1906) );
  AO22X1_LVT csr_U1602 ( .A1(csr_n493), .A2(csr_n_T_44[16]), .A3(csr_wdata_22_), .A4(csr_n491), .Y(csr_N1513) );
  MUX21X1_LVT csr_U1601 ( .A1(csr_io_pc[22]), .A2(csr_wdata_22_), .S0(csr_n515), .Y(csr_net35238) );
  AO22X1_LVT csr_U1600 ( .A1(csr_n1159), .A2(csr_io_tval[22]), .A3(
        csr_wdata_22_), .A4(csr_n1158), .Y(csr_N1404) );
  AO22X1_LVT csr_U1599 ( .A1(csr_n1152), .A2(csr_io_tval[22]), .A3(
        csr_wdata_22_), .A4(csr_n1151), .Y(csr_N1015) );
  AO22X1_LVT csr_U1598 ( .A1(csr_n498), .A2(csr_n_T_52[16]), .A3(csr_wdata_22_), .A4(csr_n1149), .Y(csr_N1907) );
  AO22X1_LVT csr_U1597 ( .A1(csr_n493), .A2(csr_n_T_44[18]), .A3(csr_wdata_24_), .A4(csr_n491), .Y(csr_N1515) );
  MUX21X1_LVT csr_U1596 ( .A1(csr_io_pc[24]), .A2(csr_wdata_24_), .S0(csr_n515), .Y(csr_net35232) );
  AO22X1_LVT csr_U1595 ( .A1(csr_n1159), .A2(csr_io_tval[24]), .A3(
        csr_wdata_24_), .A4(csr_n1158), .Y(csr_N1406) );
  AO22X1_LVT csr_U1594 ( .A1(csr_n1152), .A2(csr_io_tval[24]), .A3(
        csr_wdata_24_), .A4(csr_n1151), .Y(csr_N1017) );
  AO22X1_LVT csr_U1593 ( .A1(csr_n496), .A2(csr_n_T_52[18]), .A3(csr_wdata_24_), .A4(csr_n1149), .Y(csr_N1909) );
  NAND2X0_LVT csr_U1592 ( .A1(csr_n1613), .A2(csr_n1064), .Y(
        csr_io_rw_rdata[24]) );
  NOR4X1_LVT csr_U1591 ( .A1(csr_n1612), .A2(csr_n1063), .A3(csr_n1606), .A4(
        csr_n1607), .Y(csr_n1064) );
  NAND4X0_LVT csr_U1590 ( .A1(csr_n1061), .A2(csr_n1060), .A3(csr_n1059), .A4(
        csr_n1058), .Y(csr_n1063) );
  NAND2X0_LVT csr_U1589 ( .A1(csr_n1162), .A2(csr_io_time[24]), .Y(csr_n1058)
         );
  AND4X1_LVT csr_U1588 ( .A1(csr_n1057), .A2(csr_n1056), .A3(csr_n1055), .A4(
        csr_n1054), .Y(csr_n1059) );
  NAND2X0_LVT csr_U1587 ( .A1(csr_n1507), .A2(io_ptw_pmp_3_cfg_r), .Y(
        csr_n1054) );
  NAND2X0_LVT csr_U1586 ( .A1(csr_n1487), .A2(csr_reg_stvec_24_), .Y(csr_n1055) );
  AOI22X1_LVT csr_U1585 ( .A1(csr_n1689), .A2(csr_n_T_45_24_), .A3(csr_n1493), 
        .A4(csr_reg_dpc_24_), .Y(csr_n1056) );
  NAND2X0_LVT csr_U1584 ( .A1(csr_n1153), .A2(csr_n_T_383[24]), .Y(csr_n1057)
         );
  AO22X1_LVT csr_U1583 ( .A1(csr_n494), .A2(csr_n_T_44[19]), .A3(csr_wdata_25_), .A4(csr_n491), .Y(csr_N1516) );
  MUX21X1_LVT csr_U1582 ( .A1(csr_io_pc[25]), .A2(csr_wdata_25_), .S0(csr_n513), .Y(csr_net34805) );
  AO22X1_LVT csr_U1581 ( .A1(csr_n1159), .A2(csr_io_tval[25]), .A3(
        csr_wdata_25_), .A4(csr_n1158), .Y(csr_N1407) );
  AO22X1_LVT csr_U1580 ( .A1(csr_n1152), .A2(csr_io_tval[25]), .A3(
        csr_wdata_25_), .A4(csr_n1151), .Y(csr_N1018) );
  AO22X1_LVT csr_U1579 ( .A1(csr_n497), .A2(csr_n_T_52[19]), .A3(csr_wdata_25_), .A4(csr_n1149), .Y(csr_N1910) );
  AO22X1_LVT csr_U1578 ( .A1(csr_n1129), .A2(csr_n_T_44[20]), .A3(
        csr_wdata_26_), .A4(csr_n491), .Y(csr_N1517) );
  MUX21X1_LVT csr_U1577 ( .A1(csr_io_pc[26]), .A2(csr_wdata_26_), .S0(csr_n514), .Y(csr_net35004) );
  AO22X1_LVT csr_U1576 ( .A1(csr_n1159), .A2(csr_io_tval[26]), .A3(
        csr_wdata_26_), .A4(csr_n1158), .Y(csr_N1408) );
  AO22X1_LVT csr_U1575 ( .A1(csr_n1152), .A2(csr_io_tval[26]), .A3(
        csr_wdata_26_), .A4(csr_n1151), .Y(csr_N1019) );
  AO22X1_LVT csr_U1574 ( .A1(csr_n498), .A2(csr_n_T_52[20]), .A3(csr_wdata_26_), .A4(csr_n1149), .Y(csr_N1911) );
  AO22X1_LVT csr_U1573 ( .A1(csr_n494), .A2(csr_n_T_44[23]), .A3(csr_wdata_29_), .A4(csr_n491), .Y(csr_N1520) );
  MUX21X1_LVT csr_U1572 ( .A1(csr_io_pc[29]), .A2(csr_wdata_29_), .S0(csr_n514), .Y(csr_net34995) );
  MUX21X1_LVT csr_U1571 ( .A1(csr_io_pc[29]), .A2(csr_wdata_29_), .S0(csr_n515), .Y(csr_net35217) );
  AO22X1_LVT csr_U1570 ( .A1(csr_n1159), .A2(csr_io_tval[29]), .A3(
        csr_wdata_29_), .A4(csr_n1158), .Y(csr_N1411) );
  AO22X1_LVT csr_U1569 ( .A1(csr_n1152), .A2(csr_io_tval[29]), .A3(
        csr_wdata_29_), .A4(csr_n1151), .Y(csr_N1022) );
  AO22X1_LVT csr_U1568 ( .A1(csr_n496), .A2(csr_n_T_52[23]), .A3(csr_wdata_29_), .A4(csr_n1149), .Y(csr_N1914) );
  NAND3X0_LVT csr_U1567 ( .A1(csr_n1053), .A2(csr_n1052), .A3(csr_n1051), .Y(
        csr_io_rw_rdata[29]) );
  NOR4X1_LVT csr_U1566 ( .A1(csr_n1626), .A2(csr_n1050), .A3(csr_n1049), .A4(
        csr_n1623), .Y(csr_n1051) );
  AO21X1_LVT csr_U1565 ( .A1(csr_n1153), .A2(csr_n_T_383[29]), .A3(csr_n1048), 
        .Y(csr_n1050) );
  AO21X1_LVT csr_U1564 ( .A1(csr_n1487), .A2(csr_reg_stvec_29_), .A3(csr_n1047), .Y(csr_n1048) );
  AO22X1_LVT csr_U1563 ( .A1(csr_n1689), .A2(csr_n_T_45_29_), .A3(csr_n1493), 
        .A4(csr_reg_dpc_29_), .Y(csr_n1047) );
  NOR3X0_LVT csr_U1562 ( .A1(csr_n1622), .A2(csr_n1620), .A3(csr_n1046), .Y(
        csr_n1053) );
  OR3X1_LVT csr_U1561 ( .A1(csr_n1045), .A2(csr_n1044), .A3(csr_n1625), .Y(
        csr_n1046) );
  AO22X1_LVT csr_U1560 ( .A1(csr_n1162), .A2(csr_io_time[29]), .A3(csr_n1480), 
        .A4(io_ptw_pmp_0_addr[29]), .Y(csr_n1044) );
  AO22X1_LVT csr_U1559 ( .A1(csr_n494), .A2(csr_n_T_44[24]), .A3(csr_wdata_30_), .A4(csr_n491), .Y(csr_N1521) );
  MUX21X1_LVT csr_U1558 ( .A1(csr_io_pc[30]), .A2(csr_wdata_30_), .S0(csr_n515), .Y(csr_net35214) );
  MUX21X1_LVT csr_U1557 ( .A1(csr_io_pc[30]), .A2(csr_wdata_30_), .S0(csr_n513), .Y(csr_net34790) );
  AO22X1_LVT csr_U1556 ( .A1(csr_wdata_30_), .A2(csr_n1158), .A3(csr_n1159), 
        .A4(csr_io_tval[30]), .Y(csr_N1412) );
  AO22X1_LVT csr_U1555 ( .A1(csr_wdata_30_), .A2(csr_n1151), .A3(csr_n1152), 
        .A4(csr_io_tval[30]), .Y(csr_N1023) );
  AO22X1_LVT csr_U1554 ( .A1(csr_n498), .A2(csr_n_T_52[24]), .A3(csr_wdata_30_), .A4(csr_n1149), .Y(csr_N1915) );
  OR2X1_LVT csr_U1553 ( .A1(csr_n1043), .A2(csr_n1628), .Y(csr_io_rw_rdata[30]) );
  NAND4X0_LVT csr_U1552 ( .A1(csr_n1042), .A2(csr_n1040), .A3(csr_n1039), .A4(
        csr_n1038), .Y(csr_n1043) );
  NAND2X0_LVT csr_U1551 ( .A1(csr_n1162), .A2(csr_io_time[30]), .Y(csr_n1038)
         );
  AOI21X1_LVT csr_U1550 ( .A1(csr_n1153), .A2(csr_n_T_383[30]), .A3(csr_n1037), 
        .Y(csr_n1039) );
  NAND4X0_LVT csr_U1549 ( .A1(csr_n1036), .A2(csr_n1035), .A3(csr_n1034), .A4(
        csr_n1033), .Y(csr_n1037) );
  NAND2X0_LVT csr_U1548 ( .A1(csr_n1510), .A2(csr_reg_dscratch[30]), .Y(
        csr_n1033) );
  NAND2X0_LVT csr_U1547 ( .A1(csr_n1493), .A2(csr_reg_dpc_30_), .Y(csr_n1034)
         );
  AOI21X1_LVT csr_U1546 ( .A1(csr_n_T_45_30_), .A2(csr_n1689), .A3(csr_n1627), 
        .Y(csr_n1035) );
  NAND2X0_LVT csr_U1545 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[30]), .Y(
        csr_n1036) );
  AOI22X1_LVT csr_U1544 ( .A1(csr_n1160), .A2(csr_n_T_444[30]), .A3(csr_n1506), 
        .A4(csr_reg_sepc_30_), .Y(csr_n1042) );
  AO22X1_LVT csr_U1543 ( .A1(csr_n495), .A2(csr_n_T_44[26]), .A3(csr_wdata_32_), .A4(csr_n491), .Y(csr_N1523) );
  MUX21X1_LVT csr_U1542 ( .A1(csr_io_pc[32]), .A2(csr_wdata_32_), .S0(csr_n515), .Y(csr_net35208) );
  MUX21X1_LVT csr_U1541 ( .A1(csr_io_pc[32]), .A2(csr_wdata_32_), .S0(csr_n513), .Y(csr_net34784) );
  AO22X1_LVT csr_U1540 ( .A1(csr_n1159), .A2(csr_io_tval[32]), .A3(
        csr_wdata_32_), .A4(csr_n1158), .Y(csr_N1414) );
  AO22X1_LVT csr_U1539 ( .A1(csr_n1152), .A2(csr_io_tval[32]), .A3(
        csr_wdata_32_), .A4(csr_n1151), .Y(csr_N1025) );
  OR3X1_LVT csr_U1538 ( .A1(csr_n1032), .A2(csr_n1031), .A3(csr_n1633), .Y(
        csr_io_rw_rdata[32]) );
  NAND4X0_LVT csr_U1537 ( .A1(csr_n1030), .A2(csr_n1029), .A3(csr_n1028), .A4(
        csr_n1027), .Y(csr_n1031) );
  NAND2X0_LVT csr_U1536 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[32]), .Y(
        csr_n1027) );
  AOI22X1_LVT csr_U1535 ( .A1(csr_n1689), .A2(csr_n_T_45_32_), .A3(csr_n1493), 
        .A4(csr_reg_dpc_32_), .Y(csr_n1028) );
  NAND2X0_LVT csr_U1534 ( .A1(csr_n1153), .A2(csr_n_T_383[32]), .Y(csr_n1029)
         );
  NAND2X0_LVT csr_U1533 ( .A1(csr_n1506), .A2(csr_reg_sepc_32_), .Y(csr_n1030)
         );
  AO22X1_LVT csr_U1532 ( .A1(csr_n1160), .A2(csr_n_T_444[32]), .A3(csr_n1485), 
        .A4(csr_reg_mscratch[32]), .Y(csr_n1032) );
  AO22X1_LVT csr_U1531 ( .A1(csr_n1128), .A2(csr_wdata_33_), .A3(
        csr_n_T_44[27]), .A4(csr_n495), .Y(csr_N1524) );
  MUX21X1_LVT csr_U1530 ( .A1(csr_io_pc[33]), .A2(csr_wdata_33_), .S0(csr_n514), .Y(csr_net34983) );
  MUX21X1_LVT csr_U1529 ( .A1(csr_io_pc[33]), .A2(csr_wdata_33_), .S0(csr_n515), .Y(csr_net35205) );
  MUX21X1_LVT csr_U1528 ( .A1(csr_io_pc[33]), .A2(csr_wdata_33_), .S0(csr_n513), .Y(csr_net34781) );
  AO22X1_LVT csr_U1527 ( .A1(csr_n1158), .A2(csr_wdata_33_), .A3(
        csr_io_tval[33]), .A4(csr_n1159), .Y(csr_N1415) );
  AO22X1_LVT csr_U1526 ( .A1(csr_n1151), .A2(csr_wdata_33_), .A3(
        csr_io_tval[33]), .A4(csr_n1152), .Y(csr_N1026) );
  AO22X1_LVT csr_U1525 ( .A1(csr_n1149), .A2(csr_wdata_33_), .A3(
        csr_n_T_52[27]), .A4(csr_n496), .Y(csr_N1918) );
  AO22X1_LVT csr_U1524 ( .A1(csr_n1129), .A2(csr_n_T_44[28]), .A3(
        csr_wdata_34_), .A4(csr_n491), .Y(csr_N1525) );
  MUX21X1_LVT csr_U1523 ( .A1(csr_io_pc[34]), .A2(csr_wdata_34_), .S0(csr_n513), .Y(csr_net34778) );
  AO22X1_LVT csr_U1522 ( .A1(csr_n1159), .A2(csr_io_tval[34]), .A3(
        csr_wdata_34_), .A4(csr_n1158), .Y(csr_N1416) );
  AO22X1_LVT csr_U1521 ( .A1(csr_n1152), .A2(csr_io_tval[34]), .A3(
        csr_wdata_34_), .A4(csr_n1151), .Y(csr_N1027) );
  OR3X1_LVT csr_U1520 ( .A1(csr_n1025), .A2(csr_n1024), .A3(csr_n1638), .Y(
        csr_io_rw_rdata[34]) );
  NAND4X0_LVT csr_U1519 ( .A1(csr_n1023), .A2(csr_n1022), .A3(csr_n1021), .A4(
        csr_n1020), .Y(csr_n1024) );
  NAND2X0_LVT csr_U1518 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[34]), .Y(
        csr_n1020) );
  AOI22X1_LVT csr_U1517 ( .A1(csr_n1689), .A2(csr_n_T_45_34_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[34]), .Y(csr_n1021) );
  NAND2X0_LVT csr_U1516 ( .A1(csr_n1153), .A2(csr_n_T_383[34]), .Y(csr_n1022)
         );
  NAND2X0_LVT csr_U1515 ( .A1(csr_n1506), .A2(csr_reg_sepc_34_), .Y(csr_n1023)
         );
  AO22X1_LVT csr_U1514 ( .A1(csr_n1160), .A2(csr_n_T_444[34]), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[34]), .Y(csr_n1025) );
  AO22X1_LVT csr_U1513 ( .A1(csr_n_T_44[30]), .A2(csr_n495), .A3(csr_wdata_36_), .A4(csr_n491), .Y(csr_N1527) );
  AO22X1_LVT csr_U1512 ( .A1(csr_n495), .A2(csr_n_T_44[31]), .A3(csr_wdata_37_), .A4(csr_n491), .Y(csr_N1528) );
  AO22X1_LVT csr_U1511 ( .A1(csr_n1159), .A2(csr_io_tval[37]), .A3(
        csr_wdata_37_), .A4(csr_n1158), .Y(csr_N1419) );
  AO22X1_LVT csr_U1510 ( .A1(csr_n1152), .A2(csr_io_tval[37]), .A3(
        csr_wdata_37_), .A4(csr_n1151), .Y(csr_N1030) );
  AO22X1_LVT csr_U1509 ( .A1(csr_n498), .A2(csr_n_T_52[31]), .A3(csr_wdata_37_), .A4(csr_n1149), .Y(csr_N1922) );
  OR2X1_LVT csr_U1508 ( .A1(csr_n1019), .A2(csr_n1648), .Y(csr_io_rw_rdata[37]) );
  NAND4X0_LVT csr_U1507 ( .A1(csr_n1018), .A2(csr_n1017), .A3(csr_n1016), .A4(
        csr_n1015), .Y(csr_n1019) );
  NAND2X0_LVT csr_U1506 ( .A1(csr_n1162), .A2(csr_n1962), .Y(csr_n1015) );
  NAND2X0_LVT csr_U1505 ( .A1(csr_n1153), .A2(csr_n_T_383[37]), .Y(csr_n1016)
         );
  AOI22X1_LVT csr_U1504 ( .A1(csr_n1689), .A2(csr_n_T_45_37_), .A3(csr_n1487), 
        .A4(csr_reg_stvec_37_), .Y(csr_n1017) );
  AOI22X1_LVT csr_U1503 ( .A1(csr_n1160), .A2(csr_n_T_444[37]), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[37]), .Y(csr_n1018) );
  MUX21X1_LVT csr_U1502 ( .A1(csr_io_pc[38]), .A2(csr_wdata_38_), .S0(csr_n514), .Y(csr_net34968) );
  MUX21X1_LVT csr_U1501 ( .A1(csr_io_pc[38]), .A2(csr_wdata_38_), .S0(csr_n515), .Y(csr_net35190) );
  MUX21X1_LVT csr_U1500 ( .A1(csr_io_pc[38]), .A2(csr_wdata_38_), .S0(csr_n513), .Y(csr_net34766) );
  AO22X1_LVT csr_U1499 ( .A1(csr_wdata_38_), .A2(csr_n1158), .A3(csr_n1159), 
        .A4(csr_io_tval[38]), .Y(csr_N1420) );
  AO22X1_LVT csr_U1498 ( .A1(csr_wdata_38_), .A2(csr_n1151), .A3(csr_n1152), 
        .A4(csr_io_tval[38]), .Y(csr_N1031) );
  AO22X1_LVT csr_U1497 ( .A1(csr_n1128), .A2(csr_wdata_40_), .A3(
        csr_n_T_44[34]), .A4(csr_n495), .Y(csr_N1531) );
  AO22X1_LVT csr_U1496 ( .A1(csr_n1149), .A2(csr_wdata_40_), .A3(
        csr_n_T_52[34]), .A4(csr_n496), .Y(csr_N1925) );
  NAND3X0_LVT csr_U1495 ( .A1(csr_n481), .A2(csr_n1675), .A3(csr_n1014), .Y(
        csr_io_rw_rdata[40]) );
  NAND2X0_LVT csr_U1494 ( .A1(csr_n1162), .A2(csr_n1959), .Y(csr_n1011) );
  AOI22X1_LVT csr_U1493 ( .A1(csr_n1689), .A2(csr_n_T_45_40_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[40]), .Y(csr_n1012) );
  AO22X1_LVT csr_U1492 ( .A1(csr_n1128), .A2(csr_wdata_41_), .A3(
        csr_n_T_44[35]), .A4(csr_n494), .Y(csr_N1532) );
  AO22X1_LVT csr_U1491 ( .A1(csr_n1149), .A2(csr_wdata_41_), .A3(
        csr_n_T_52[35]), .A4(csr_n496), .Y(csr_N1926) );
  NAND3X0_LVT csr_U1490 ( .A1(csr_n481), .A2(csr_n1676), .A3(csr_n1010), .Y(
        csr_io_rw_rdata[41]) );
  NOR3X0_LVT csr_U1489 ( .A1(csr_n1009), .A2(csr_n1008), .A3(csr_n1007), .Y(
        csr_n1010) );
  AO22X1_LVT csr_U1488 ( .A1(csr_n1508), .A2(csr_reg_sscratch[41]), .A3(
        csr_n1162), .A4(csr_n1958), .Y(csr_n1007) );
  AO22X1_LVT csr_U1487 ( .A1(csr_n1128), .A2(csr_wdata_42_), .A3(
        csr_n_T_44[36]), .A4(csr_n495), .Y(csr_N1533) );
  AO22X1_LVT csr_U1486 ( .A1(csr_n1149), .A2(csr_wdata_42_), .A3(
        csr_n_T_52[36]), .A4(csr_n497), .Y(csr_N1927) );
  NAND3X0_LVT csr_U1485 ( .A1(csr_n481), .A2(csr_n1677), .A3(csr_n1006), .Y(
        csr_io_rw_rdata[42]) );
  NAND2X0_LVT csr_U1484 ( .A1(csr_n1162), .A2(csr_n1957), .Y(csr_n1003) );
  AOI22X1_LVT csr_U1483 ( .A1(csr_n1689), .A2(csr_n_T_45_42_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_5_cfg_x), .Y(csr_n1004) );
  AO22X1_LVT csr_U1482 ( .A1(csr_n1128), .A2(csr_wdata_45_), .A3(
        csr_n_T_44[39]), .A4(csr_n495), .Y(csr_N1536) );
  AO22X1_LVT csr_U1481 ( .A1(csr_n1149), .A2(csr_wdata_45_), .A3(
        csr_n_T_52[39]), .A4(csr_n496), .Y(csr_N1930) );
  OR2X1_LVT csr_U1480 ( .A1(csr_n1002), .A2(csr_n1690), .Y(csr_io_rw_rdata[45]) );
  AOI22X1_LVT csr_U1479 ( .A1(csr_n1689), .A2(csr_n_T_45_45_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[45]), .Y(csr_n999) );
  AOI22X1_LVT csr_U1478 ( .A1(csr_n1508), .A2(csr_reg_sscratch[45]), .A3(
        csr_n1162), .A4(csr_n1954), .Y(csr_n1001) );
  AO22X1_LVT csr_U1477 ( .A1(csr_n_T_44[40]), .A2(csr_n1129), .A3(csr_n492), 
        .A4(csr_wdata_46_), .Y(csr_N1537) );
  AO22X1_LVT csr_U1476 ( .A1(csr_n_T_52[40]), .A2(csr_n1150), .A3(csr_n1149), 
        .A4(csr_wdata_46_), .Y(csr_N1931) );
  OR3X1_LVT csr_U1475 ( .A1(csr_n998), .A2(csr_n997), .A3(csr_n1679), .Y(
        csr_io_rw_rdata[46]) );
  AO22X1_LVT csr_U1474 ( .A1(csr_n1485), .A2(csr_reg_mscratch[46]), .A3(
        csr_n1162), .A4(csr_n1953), .Y(csr_n997) );
  AO22X1_LVT csr_U1473 ( .A1(csr_n1128), .A2(csr_wdata_49_), .A3(
        csr_n_T_44[43]), .A4(csr_n495), .Y(csr_N1540) );
  AO22X1_LVT csr_U1472 ( .A1(csr_n1128), .A2(csr_wdata_48_), .A3(
        csr_n_T_44[42]), .A4(csr_n1129), .Y(csr_N1539) );
  AO22X1_LVT csr_U1471 ( .A1(csr_n1149), .A2(csr_wdata_48_), .A3(
        csr_n_T_52[42]), .A4(csr_n497), .Y(csr_N1933) );
  NAND3X0_LVT csr_U1470 ( .A1(csr_n481), .A2(csr_n1681), .A3(csr_n996), .Y(
        csr_io_rw_rdata[48]) );
  NAND2X0_LVT csr_U1469 ( .A1(csr_n1162), .A2(csr_n1951), .Y(csr_n993) );
  AOI22X1_LVT csr_U1468 ( .A1(csr_n1689), .A2(csr_n_T_45_48_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_6_cfg_r), .Y(csr_n994) );
  AO22X1_LVT csr_U1467 ( .A1(csr_n1149), .A2(csr_wdata_49_), .A3(
        csr_n_T_52[43]), .A4(csr_n496), .Y(csr_N1934) );
  NAND3X0_LVT csr_U1466 ( .A1(csr_n481), .A2(csr_n1682), .A3(csr_n992), .Y(
        csr_io_rw_rdata[49]) );
  NAND2X0_LVT csr_U1465 ( .A1(csr_n1162), .A2(csr_n1950), .Y(csr_n989) );
  AOI22X1_LVT csr_U1464 ( .A1(csr_n1689), .A2(csr_n_T_45_49_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_6_cfg_w), .Y(csr_n990) );
  NAND3X0_LVT csr_U1463 ( .A1(csr_n481), .A2(csr_n1683), .A3(csr_n988), .Y(
        csr_io_rw_rdata[50]) );
  NAND2X0_LVT csr_U1462 ( .A1(csr_n1162), .A2(csr_n1949), .Y(csr_n985) );
  AOI22X1_LVT csr_U1461 ( .A1(csr_n1689), .A2(csr_n_T_45_50_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[50]), .Y(csr_n986) );
  AO22X1_LVT csr_U1460 ( .A1(csr_n1128), .A2(csr_wdata_53_), .A3(
        csr_n_T_44[47]), .A4(csr_n1129), .Y(csr_N1544) );
  AO22X1_LVT csr_U1459 ( .A1(csr_n1149), .A2(csr_wdata_53_), .A3(
        csr_n_T_52[47]), .A4(csr_n497), .Y(csr_N1938) );
  OR2X1_LVT csr_U1458 ( .A1(csr_n984), .A2(csr_n1690), .Y(csr_io_rw_rdata[53])
         );
  AOI22X1_LVT csr_U1457 ( .A1(csr_n1689), .A2(csr_n_T_45_53_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[53]), .Y(csr_n981) );
  AOI22X1_LVT csr_U1456 ( .A1(csr_n1508), .A2(csr_reg_sscratch[53]), .A3(
        csr_n1162), .A4(csr_n1946), .Y(csr_n983) );
  AO22X1_LVT csr_U1455 ( .A1(csr_n1128), .A2(csr_wdata_54_), .A3(
        csr_n_T_44[48]), .A4(csr_n494), .Y(csr_N1545) );
  OR2X1_LVT csr_U1454 ( .A1(csr_n980), .A2(csr_n1690), .Y(csr_io_rw_rdata[54])
         );
  AOI22X1_LVT csr_U1453 ( .A1(csr_n1689), .A2(csr_n_T_45_54_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[54]), .Y(csr_n977) );
  AOI22X1_LVT csr_U1452 ( .A1(csr_n1508), .A2(csr_reg_sscratch[54]), .A3(
        csr_n1162), .A4(csr_n1945), .Y(csr_n979) );
  AO22X1_LVT csr_U1451 ( .A1(csr_n1128), .A2(csr_wdata_57_), .A3(
        csr_n_T_44[51]), .A4(csr_n495), .Y(csr_N1548) );
  AO22X1_LVT csr_U1450 ( .A1(csr_n1128), .A2(csr_wdata_56_), .A3(
        csr_n_T_44[50]), .A4(csr_n494), .Y(csr_N1547) );
  AO22X1_LVT csr_U1449 ( .A1(csr_n1149), .A2(csr_wdata_56_), .A3(
        csr_n_T_52[50]), .A4(csr_n497), .Y(csr_N1941) );
  NAND3X0_LVT csr_U1448 ( .A1(csr_n481), .A2(csr_n1686), .A3(csr_n976), .Y(
        csr_io_rw_rdata[56]) );
  NAND2X0_LVT csr_U1447 ( .A1(csr_n1162), .A2(csr_n1943), .Y(csr_n973) );
  AOI22X1_LVT csr_U1446 ( .A1(csr_n1689), .A2(csr_n_T_45_56_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[56]), .Y(csr_n974) );
  AO22X1_LVT csr_U1445 ( .A1(csr_n1149), .A2(csr_wdata_57_), .A3(
        csr_n_T_52[51]), .A4(csr_n497), .Y(csr_N1942) );
  NAND4X0_LVT csr_U1444 ( .A1(csr_n481), .A2(csr_n1687), .A3(csr_n475), .A4(
        csr_n972), .Y(csr_io_rw_rdata[57]) );
  AO22X1_LVT csr_U1443 ( .A1(csr_n1689), .A2(csr_n_T_45_57_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[57]), .Y(csr_n971) );
  NAND4X0_LVT csr_U1442 ( .A1(csr_n481), .A2(csr_n1688), .A3(csr_n474), .A4(
        csr_n970), .Y(csr_io_rw_rdata[58]) );
  AO22X1_LVT csr_U1441 ( .A1(csr_n1689), .A2(csr_n_T_45_58_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[58]), .Y(csr_n969) );
  AO22X1_LVT csr_U1440 ( .A1(csr_n1128), .A2(csr_wdata_61_), .A3(
        csr_n_T_44[55]), .A4(csr_n1129), .Y(csr_N1552) );
  AO22X1_LVT csr_U1439 ( .A1(csr_n1149), .A2(csr_wdata_61_), .A3(
        csr_n_T_52[55]), .A4(csr_n1150), .Y(csr_N1946) );
  NAND4X0_LVT csr_U1438 ( .A1(csr_n968), .A2(csr_n967), .A3(csr_n467), .A4(
        csr_n966), .Y(csr_io_rw_rdata[61]) );
  AOI22X1_LVT csr_U1437 ( .A1(csr_n1508), .A2(csr_reg_sscratch[61]), .A3(
        csr_n1162), .A4(csr_n1938), .Y(csr_n967) );
  AO22X1_LVT csr_U1436 ( .A1(csr_n1128), .A2(csr_wdata_62_), .A3(
        csr_n_T_44[56]), .A4(csr_n494), .Y(csr_N1553) );
  AO22X1_LVT csr_U1435 ( .A1(csr_n1149), .A2(csr_wdata_62_), .A3(
        csr_n_T_52[56]), .A4(csr_n1150), .Y(csr_N1947) );
  OR2X1_LVT csr_U1434 ( .A1(csr_n965), .A2(csr_n1690), .Y(csr_io_rw_rdata[62])
         );
  AOI22X1_LVT csr_U1433 ( .A1(csr_n1689), .A2(csr_n_T_45_62_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[62]), .Y(csr_n962) );
  AOI22X1_LVT csr_U1432 ( .A1(csr_n1508), .A2(csr_reg_sscratch[62]), .A3(
        csr_n1162), .A4(csr_n1937), .Y(csr_n964) );
  AO22X1_LVT csr_U1431 ( .A1(csr_n1128), .A2(csr_wdata_63_), .A3(
        csr_n_T_44[57]), .A4(csr_n1129), .Y(csr_N1554) );
  OAI22X1_LVT csr_U1430 ( .A1(csr_n959), .A2(csr_n958), .A3(csr_n957), .A4(
        csr_n1483), .Y(csr_N1430) );
  AO22X1_LVT csr_U1429 ( .A1(csr_io_tval[0]), .A2(csr_n1159), .A3(csr_wdata_0_), .A4(csr_n1158), .Y(csr_N1382) );
  AO22X1_LVT csr_U1428 ( .A1(csr_io_tval[0]), .A2(csr_n1152), .A3(csr_wdata_0_), .A4(csr_n1151), .Y(csr_N993) );
  AO22X1_LVT csr_U1427 ( .A1(csr_n1498), .A2(csr_n1202), .A3(csr_wdata_0_), 
        .A4(csr_n955), .Y(csr_N881) );
  NAND2X0_LVT csr_U1426 ( .A1(csr_n1495), .A2(csr_n_T_389[8]), .Y(csr_n947) );
  NAND2X0_LVT csr_U1425 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[8]), .Y(
        csr_n948) );
  AO22X1_LVT csr_U1424 ( .A1(csr_n946), .A2(csr_n945), .A3(csr_n944), .A4(
        csr_n590), .Y(csr_n2161) );
  MUX21X1_LVT csr_U1423 ( .A1(csr_io_status_debug), .A2(csr_n943), .S0(
        csr_n945), .Y(csr_n944) );
  INVX1_LVT csr_U1422 ( .A(csr_n942), .Y(csr_n943) );
  AO21X1_LVT csr_U1421 ( .A1(csr_n1257), .A2(csr_n1139), .A3(csr_n1356), .Y(
        csr_n945) );
  AND2X1_LVT csr_U1420 ( .A1(csr_n1499), .A2(csr_n941), .Y(csr_n946) );
  NAND2X0_LVT csr_U1419 ( .A1(csr_n950), .A2(io_ptw_status_prv[1]), .Y(
        csr_n938) );
  AND2X1_LVT csr_U1418 ( .A1(io_ptw_status_prv[0]), .A2(csr_n1903), .Y(
        csr_n950) );
  NAND3X0_LVT csr_U1417 ( .A1(csr_n951), .A2(csr_io_rw_addr[9]), .A3(csr_n937), 
        .Y(csr_n939) );
  MUX21X1_LVT csr_U1416 ( .A1(csr_n_1929_), .A2(csr_n_T_389_1), .S0(
        csr_io_rw_addr[10]), .Y(csr_n937) );
  AO21X1_LVT csr_U1415 ( .A1(csr_n1199), .A2(csr_n936), .A3(csr_n500), .Y(
        csr_n951) );
  MUX21X1_LVT csr_U1414 ( .A1(csr_n_1930_), .A2(csr_n_T_389_0), .S0(
        csr_io_rw_addr[10]), .Y(csr_n936) );
  NAND2X0_LVT csr_U1413 ( .A1(csr_n1441), .A2(csr_n952), .Y(csr_n940) );
  AND3X1_LVT csr_U1412 ( .A1(csr_n1139), .A2(csr_n1903), .A3(n9516), .Y(
        csr_n952) );
  OR2X1_LVT csr_U1411 ( .A1(csr_n1257), .A2(csr_n1255), .Y(csr_n1441) );
  OA22X1_LVT csr_U1410 ( .A1(csr_n_T_389_0), .A2(csr_n935), .A3(csr_n934), 
        .A4(csr_n933), .Y(csr_n2156) );
  MUX21X1_LVT csr_U1409 ( .A1(io_ptw_status_prv[0]), .A2(csr_wdata_0_), .S0(
        csr_n932), .Y(csr_n933) );
  NAND2X0_LVT csr_U1408 ( .A1(csr_wdata_11_), .A2(csr_n1450), .Y(csr_n931) );
  NAND2X0_LVT csr_U1407 ( .A1(csr_n928), .A2(csr_n501), .Y(csr_n929) );
  NAND2X0_LVT csr_U1406 ( .A1(csr_n925), .A2(csr_n451), .Y(csr_n926) );
  NAND2X0_LVT csr_U1405 ( .A1(csr_n1041), .A2(csr_io_exception), .Y(csr_n927)
         );
  AO22X1_LVT csr_U1404 ( .A1(csr_n493), .A2(csr_n455), .A3(csr_wdata_6_), .A4(
        csr_n492), .Y(csr_N1497) );
  MUX21X1_LVT csr_U1403 ( .A1(csr_io_pc[6]), .A2(csr_wdata_6_), .S0(csr_n513), 
        .Y(csr_net34862) );
  AO22X1_LVT csr_U1402 ( .A1(csr_n1159), .A2(csr_io_tval[6]), .A3(csr_wdata_6_), .A4(csr_n1158), .Y(csr_N1388) );
  AO22X1_LVT csr_U1401 ( .A1(csr_n1152), .A2(csr_io_tval[6]), .A3(csr_wdata_6_), .A4(csr_n1151), .Y(csr_N999) );
  AO22X1_LVT csr_U1400 ( .A1(csr_n498), .A2(csr_n456), .A3(csr_wdata_6_), .A4(
        csr_n1149), .Y(csr_N1891) );
  NAND2X0_LVT csr_U1399 ( .A1(csr_n_T_383[6]), .A2(csr_n1153), .Y(csr_n924) );
  AO22X1_LVT csr_U1398 ( .A1(csr_n1159), .A2(csr_io_tval[4]), .A3(csr_wdata_4_), .A4(csr_n1158), .Y(csr_N1386) );
  AO22X1_LVT csr_U1397 ( .A1(csr_n1152), .A2(csr_io_tval[4]), .A3(csr_wdata_4_), .A4(csr_n1151), .Y(csr_N997) );
  AO21X1_LVT csr_U1396 ( .A1(csr_n1164), .A2(io_fpu_fcsr_flags_bits[4]), .A3(
        csr_n922), .Y(csr_n_GEN_345[4]) );
  MUX21X1_LVT csr_U1395 ( .A1(csr_wdata_4_), .A2(csr_read_fcsr_4_), .S0(
        csr_n1163), .Y(csr_n922) );
  AO22X1_LVT csr_U1394 ( .A1(csr_n1129), .A2(csr_n_T_44[3]), .A3(csr_wdata_9_), 
        .A4(csr_n492), .Y(csr_N1500) );
  AO22X1_LVT csr_U1393 ( .A1(csr_n494), .A2(csr_n_T_44[1]), .A3(csr_wdata_7_), 
        .A4(csr_n492), .Y(csr_N1498) );
  NAND4X0_LVT csr_U1392 ( .A1(csr_n921), .A2(csr_n920), .A3(csr_n919), .A4(
        csr_n918), .Y(csr_N360) );
  AO21X1_LVT csr_U1391 ( .A1(csr_n1442), .A2(csr_n917), .A3(csr_n916), .Y(
        csr_n918) );
  NAND2X0_LVT csr_U1390 ( .A1(csr_n502), .A2(csr_n590), .Y(csr_n919) );
  NAND2X0_LVT csr_U1389 ( .A1(csr_n1450), .A2(csr_wdata_7_), .Y(csr_n920) );
  NOR2X0_LVT csr_U1388 ( .A1(csr_n389), .A2(csr_n1041), .Y(csr_n1450) );
  MUX21X1_LVT csr_U1387 ( .A1(csr_n1932), .A2(csr_n1934), .S0(csr_n925), .Y(
        csr_n915) );
  AND2X1_LVT csr_U1386 ( .A1(csr_n914), .A2(csr_n913), .Y(csr_n194) );
  NAND3X0_LVT csr_U1385 ( .A1(csr_n912), .A2(csr_n1934), .A3(csr_n590), .Y(
        csr_n913) );
  AO21X1_LVT csr_U1384 ( .A1(csr_n911), .A2(csr_n910), .A3(csr_n930), .Y(
        csr_n912) );
  AND2X1_LVT csr_U1383 ( .A1(csr_n909), .A2(csr_n1461), .Y(csr_n930) );
  AND2X1_LVT csr_U1382 ( .A1(csr_n908), .A2(csr_n1255), .Y(csr_n925) );
  AND3X1_LVT csr_U1381 ( .A1(csr_n451), .A2(csr_n387), .A3(csr_n501), .Y(
        csr_n909) );
  AO21X1_LVT csr_U1380 ( .A1(csr_n1026), .A2(csr_n1903), .A3(csr_n1515), .Y(
        csr_n910) );
  AND2X1_LVT csr_U1379 ( .A1(csr_n1198), .A2(csr_n1139), .Y(csr_n908) );
  INVX1_LVT csr_U1378 ( .A(csr_n1257), .Y(csr_n1198) );
  OA22X1_LVT csr_U1377 ( .A1(csr_n451), .A2(csr_n907), .A3(csr_n916), .A4(
        csr_n1255), .Y(csr_n914) );
  AND3X1_LVT csr_U1376 ( .A1(csr_n903), .A2(csr_n1202), .A3(csr_n902), .Y(
        csr_n904) );
  MUX21X1_LVT csr_U1375 ( .A1(csr_n901), .A2(csr_n900), .S0(csr_n899), .Y(
        csr_n903) );
  MUX21X1_LVT csr_U1374 ( .A1(csr_read_mideleg_1), .A2(csr_read_mideleg_9_), 
        .S0(csr_n1226), .Y(csr_n900) );
  MUX21X1_LVT csr_U1373 ( .A1(csr_n898), .A2(csr_n897), .S0(csr_n899), .Y(
        csr_n905) );
  AO22X1_LVT csr_U1372 ( .A1(csr_n896), .A2(csr_read_medeleg_8), .A3(csr_n895), 
        .A4(csr_n894), .Y(csr_n897) );
  MUX21X1_LVT csr_U1371 ( .A1(csr_n893), .A2(csr_n892), .S0(csr_n1202), .Y(
        csr_n894) );
  AND2X1_LVT csr_U1370 ( .A1(csr_read_medeleg_3_), .A2(csr_n1209), .Y(csr_n892) );
  MUX21X1_LVT csr_U1369 ( .A1(csr_read_medeleg_0), .A2(csr_read_medeleg_2_), 
        .S0(csr_n1209), .Y(csr_n893) );
  NAND2X0_LVT csr_U1368 ( .A1(csr_n890), .A2(csr_n889), .Y(csr_n898) );
  NAND2X0_LVT csr_U1367 ( .A1(csr_n896), .A2(csr_read_medeleg_12), .Y(csr_n889) );
  AND3X1_LVT csr_U1366 ( .A1(csr_n1226), .A2(csr_n891), .A3(csr_n888), .Y(
        csr_n896) );
  MUX21X1_LVT csr_U1365 ( .A1(csr_n887), .A2(csr_n886), .S0(csr_n1226), .Y(
        csr_n890) );
  NAND2X0_LVT csr_U1364 ( .A1(csr_n885), .A2(wb_cause[0]), .Y(csr_n886) );
  MUX21X1_LVT csr_U1363 ( .A1(csr_read_medeleg_13), .A2(csr_read_medeleg_15), 
        .S0(csr_n1209), .Y(csr_n885) );
  NAND2X0_LVT csr_U1362 ( .A1(csr_n884), .A2(csr_n954), .Y(csr_n887) );
  MUX21X1_LVT csr_U1361 ( .A1(csr_read_medeleg_4_), .A2(csr_read_medeleg_6), 
        .S0(csr_n1209), .Y(csr_n884) );
  NAND2X0_LVT csr_U1360 ( .A1(csr_n1451), .A2(csr_n1934), .Y(csr_n916) );
  AO21X1_LVT csr_U1359 ( .A1(csr_n503), .A2(csr_n1041), .A3(csr_n883), .Y(
        csr_n1451) );
  NAND2X0_LVT csr_U1358 ( .A1(csr_n590), .A2(csr_n1932), .Y(csr_n907) );
  NAND2X0_LVT csr_U1357 ( .A1(csr_n1514), .A2(csr_io_rw_addr[9]), .Y(csr_n882)
         );
  MUX21X1_LVT csr_U1356 ( .A1(csr_io_pc[3]), .A2(csr_wdata_3_), .S0(csr_n514), 
        .Y(csr_net35073) );
  MUX21X1_LVT csr_U1355 ( .A1(io_ptw_pmp_7_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n512), .Y(csr_n_GEN_307[3]) );
  MUX21X1_LVT csr_U1354 ( .A1(io_ptw_pmp_0_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n505), .Y(csr_n_GEN_258[3]) );
  MUX21X1_LVT csr_U1353 ( .A1(io_ptw_pmp_4_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n509), .Y(csr_n_GEN_286[3]) );
  MUX21X1_LVT csr_U1352 ( .A1(io_ptw_pmp_5_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n510), .Y(csr_n_GEN_293[3]) );
  MUX21X1_LVT csr_U1351 ( .A1(io_ptw_pmp_3_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n508), .Y(csr_n_GEN_279[3]) );
  MUX21X1_LVT csr_U1350 ( .A1(io_ptw_pmp_2_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n507), .Y(csr_n_GEN_272[3]) );
  MUX21X1_LVT csr_U1349 ( .A1(io_ptw_pmp_6_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n511), .Y(csr_n_GEN_300[3]) );
  MUX21X1_LVT csr_U1348 ( .A1(csr_io_pc[3]), .A2(csr_wdata_3_), .S0(csr_n513), 
        .Y(csr_net34871) );
  AO22X1_LVT csr_U1347 ( .A1(csr_reg_mie_3_), .A2(csr_n1503), .A3(csr_wdata_3_), .A4(csr_n1502), .Y(csr_N609) );
  AO22X1_LVT csr_U1346 ( .A1(csr_wdata_3_), .A2(csr_n1158), .A3(csr_n1159), 
        .A4(csr_io_tval[3]), .Y(csr_N1385) );
  AO22X1_LVT csr_U1345 ( .A1(csr_wdata_3_), .A2(csr_n1151), .A3(csr_n1152), 
        .A4(csr_io_tval[3]), .Y(csr_N996) );
  AO22X1_LVT csr_U1344 ( .A1(csr_n1498), .A2(csr_n1226), .A3(csr_n1468), .A4(
        csr_n1161), .Y(csr_N884) );
  AND2X1_LVT csr_U1343 ( .A1(csr_wdata_3_), .A2(csr_n503), .Y(csr_n1468) );
  AO22X1_LVT csr_U1342 ( .A1(csr_n1501), .A2(csr_n1226), .A3(csr_wdata_3_), 
        .A4(csr_n923), .Y(csr_N1273) );
  AO21X1_LVT csr_U1341 ( .A1(csr_n1164), .A2(io_fpu_fcsr_flags_bits[3]), .A3(
        csr_n881), .Y(csr_n_GEN_345[3]) );
  MUX21X1_LVT csr_U1340 ( .A1(csr_wdata_3_), .A2(csr_read_fcsr_3_), .S0(
        csr_n1163), .Y(csr_n881) );
  AND2X1_LVT csr_U1339 ( .A1(csr_n590), .A2(csr_n1910), .Y(csr_n880) );
  NAND4X0_LVT csr_U1338 ( .A1(csr_n878), .A2(csr_n877), .A3(csr_n876), .A4(
        csr_n875), .Y(csr_io_rw_rdata[3]) );
  NOR4X1_LVT csr_U1337 ( .A1(csr_n874), .A2(csr_n873), .A3(csr_n872), .A4(
        csr_n871), .Y(csr_n875) );
  AO22X1_LVT csr_U1336 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[3]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[3]), .Y(csr_n871) );
  AO22X1_LVT csr_U1335 ( .A1(csr_n1481), .A2(csr_io_bp_0_control_u), .A3(
        csr_n1167), .A4(csr_read_fcsr_3_), .Y(csr_n872) );
  NAND4X0_LVT csr_U1334 ( .A1(csr_n870), .A2(csr_n869), .A3(csr_n868), .A4(
        csr_n867), .Y(csr_n873) );
  NAND2X0_LVT csr_U1333 ( .A1(csr_n1507), .A2(io_ptw_pmp_0_cfg_a[0]), .Y(
        csr_n867) );
  OA21X1_LVT csr_U1332 ( .A1(csr_n1910), .A2(csr_n866), .A3(csr_n865), .Y(
        csr_n868) );
  AOI22X1_LVT csr_U1331 ( .A1(csr_n1689), .A2(csr_n_T_45_3_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[3]), .Y(csr_n865) );
  AOI22X1_LVT csr_U1330 ( .A1(csr_n1493), .A2(csr_reg_dpc_3_), .A3(csr_n488), 
        .A4(io_ptw_ptbr_ppn[3]), .Y(csr_n869) );
  NAND2X0_LVT csr_U1329 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[3]), .Y(
        csr_n870) );
  AND2X1_LVT csr_U1328 ( .A1(csr_n1162), .A2(csr_io_time[3]), .Y(csr_n874) );
  AOI21X1_LVT csr_U1327 ( .A1(csr_reg_mtvec_3_), .A2(csr_n1470), .A3(csr_n864), 
        .Y(csr_n876) );
  AO22X1_LVT csr_U1326 ( .A1(csr_n1502), .A2(csr_reg_mie_3_), .A3(
        csr_reg_stvec_3_), .A4(csr_n1478), .Y(csr_n864) );
  NOR4X1_LVT csr_U1325 ( .A1(csr_n863), .A2(csr_n862), .A3(csr_n861), .A4(
        csr_n859), .Y(csr_n877) );
  AO22X1_LVT csr_U1324 ( .A1(csr_n1508), .A2(csr_reg_sscratch[3]), .A3(
        csr_reg_sepc_3_), .A4(csr_n1506), .Y(csr_n859) );
  AO22X1_LVT csr_U1323 ( .A1(csr_n1160), .A2(csr_n_T_444[3]), .A3(csr_n1168), 
        .A4(csr_reg_scause[3]), .Y(csr_n861) );
  AO22X1_LVT csr_U1322 ( .A1(csr_n1485), .A2(csr_reg_mscratch[3]), .A3(
        csr_reg_mepc_3_), .A4(csr_n1489), .Y(csr_n862) );
  AO22X1_LVT csr_U1321 ( .A1(csr_n1474), .A2(io_interrupts_msip), .A3(
        csr_read_medeleg_3_), .A4(csr_n1469), .Y(csr_n863) );
  NOR4X1_LVT csr_U1320 ( .A1(csr_n856), .A2(csr_n855), .A3(csr_n854), .A4(
        csr_n853), .Y(csr_n878) );
  OR2X1_LVT csr_U1319 ( .A1(csr_n852), .A2(csr_n851), .Y(csr_n853) );
  AO22X1_LVT csr_U1318 ( .A1(csr_n1161), .A2(csr_reg_mcause[3]), .A3(csr_n1157), .A4(csr_n1934), .Y(csr_n851) );
  AO22X1_LVT csr_U1317 ( .A1(csr_n1153), .A2(csr_n_T_383[3]), .A3(csr_n1452), 
        .A4(csr_io_status_isa[3]), .Y(csr_n852) );
  AO22X1_LVT csr_U1316 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[3]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[3]), .Y(csr_n854) );
  AO22X1_LVT csr_U1315 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[3]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[3]), .Y(csr_n855) );
  AO22X1_LVT csr_U1314 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[3]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[3]), .Y(csr_n856) );
  MUX21X1_LVT csr_U1313 ( .A1(csr_wdata_7_), .A2(csr_wdata_2_), .S0(csr_n1696), 
        .Y(csr_n_GEN_155[2]) );
  MUX21X1_LVT csr_U1312 ( .A1(io_ptw_pmp_7_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n512), .Y(csr_n_GEN_307[7]) );
  MUX21X1_LVT csr_U1311 ( .A1(io_ptw_pmp_0_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n505), .Y(csr_n_GEN_258[7]) );
  MUX21X1_LVT csr_U1310 ( .A1(io_ptw_pmp_4_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n509), .Y(csr_n_GEN_286[7]) );
  MUX21X1_LVT csr_U1309 ( .A1(io_ptw_pmp_5_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n510), .Y(csr_n_GEN_293[7]) );
  MUX21X1_LVT csr_U1308 ( .A1(io_ptw_pmp_3_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n508), .Y(csr_n_GEN_279[7]) );
  MUX21X1_LVT csr_U1307 ( .A1(io_ptw_pmp_2_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n507), .Y(csr_n_GEN_272[7]) );
  MUX21X1_LVT csr_U1306 ( .A1(io_ptw_pmp_6_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n511), .Y(csr_n_GEN_300[7]) );
  MUX21X1_LVT csr_U1305 ( .A1(io_ptw_pmp_1_addr[7]), .A2(csr_wdata_7_), .S0(
        csr_n506), .Y(csr_n_GEN_265[7]) );
  AND2X1_LVT csr_U1304 ( .A1(csr_n1467), .A2(csr_n1471), .Y(csr_N469) );
  AND2X1_LVT csr_U1303 ( .A1(csr_n1499), .A2(csr_n860), .Y(csr_n1471) );
  AO22X1_LVT csr_U1302 ( .A1(csr_reg_mie_7_), .A2(csr_n1503), .A3(csr_wdata_7_), .A4(csr_n1502), .Y(csr_N613) );
  AO22X1_LVT csr_U1301 ( .A1(csr_n1158), .A2(csr_wdata_7_), .A3(csr_io_tval[7]), .A4(csr_n1159), .Y(csr_N1389) );
  AO22X1_LVT csr_U1300 ( .A1(csr_n1151), .A2(csr_wdata_7_), .A3(csr_io_tval[7]), .A4(csr_n1152), .Y(csr_N1000) );
  AO22X1_LVT csr_U1299 ( .A1(csr_n498), .A2(csr_n_T_52[1]), .A3(csr_wdata_7_), 
        .A4(csr_n1149), .Y(csr_N1892) );
  NAND3X0_LVT csr_U1298 ( .A1(csr_n850), .A2(csr_n849), .A3(csr_n848), .Y(
        csr_io_rw_rdata[7]) );
  NOR4X1_LVT csr_U1297 ( .A1(csr_n847), .A2(csr_n846), .A3(csr_n845), .A4(
        csr_n844), .Y(csr_n848) );
  AND2X1_LVT csr_U1296 ( .A1(csr_n1470), .A2(csr_reg_mtvec_7_), .Y(csr_n844)
         );
  AND2X1_LVT csr_U1295 ( .A1(csr_n1497), .A2(csr_n659), .Y(csr_n1470) );
  NAND4X0_LVT csr_U1294 ( .A1(csr_n843), .A2(csr_n842), .A3(csr_n841), .A4(
        csr_n840), .Y(csr_n845) );
  NAND2X0_LVT csr_U1293 ( .A1(csr_io_bp_0_address[7]), .A2(csr_n1490), .Y(
        csr_n840) );
  NAND2X0_LVT csr_U1292 ( .A1(csr_io_bp_0_control_tmatch[0]), .A2(csr_n1481), 
        .Y(csr_n841) );
  AND4X1_LVT csr_U1291 ( .A1(csr_n839), .A2(csr_n838), .A3(csr_n837), .A4(
        csr_n836), .Y(csr_n842) );
  NAND2X0_LVT csr_U1290 ( .A1(io_ptw_ptbr_ppn[7]), .A2(csr_n488), .Y(csr_n836)
         );
  AOI22X1_LVT csr_U1289 ( .A1(csr_n1689), .A2(csr_n_T_45_7_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[7]), .Y(csr_n837) );
  AOI22X1_LVT csr_U1288 ( .A1(csr_n1493), .A2(csr_reg_dpc_7_), .A3(csr_n1495), 
        .A4(csr_n_T_389[7]), .Y(csr_n838) );
  NAND2X0_LVT csr_U1287 ( .A1(io_ptw_pmp_0_cfg_l), .A2(csr_n1507), .Y(csr_n839) );
  NAND2X0_LVT csr_U1286 ( .A1(io_ptw_pmp_0_addr[7]), .A2(csr_n1480), .Y(
        csr_n843) );
  AO22X1_LVT csr_U1285 ( .A1(csr_n1506), .A2(csr_reg_sepc_7_), .A3(
        csr_reg_stvec_7_), .A4(csr_n1478), .Y(csr_n846) );
  AO22X1_LVT csr_U1284 ( .A1(csr_n1502), .A2(csr_reg_mie_7_), .A3(csr_n1162), 
        .A4(csr_io_time[7]), .Y(csr_n847) );
  NOR4X1_LVT csr_U1283 ( .A1(csr_n835), .A2(csr_n834), .A3(csr_n833), .A4(
        csr_n832), .Y(csr_n849) );
  AO22X1_LVT csr_U1282 ( .A1(csr_n1160), .A2(csr_n_T_444[7]), .A3(
        csr_reg_mepc_7_), .A4(csr_n1489), .Y(csr_n833) );
  AO22X1_LVT csr_U1281 ( .A1(csr_n1485), .A2(csr_reg_mscratch[7]), .A3(
        csr_n1157), .A4(csr_n1932), .Y(csr_n834) );
  AO22X1_LVT csr_U1280 ( .A1(csr_n1153), .A2(csr_n_T_383[7]), .A3(csr_n1474), 
        .A4(io_interrupts_mtip), .Y(csr_n835) );
  NOR4X1_LVT csr_U1279 ( .A1(csr_n831), .A2(csr_n830), .A3(csr_n829), .A4(
        csr_n828), .Y(csr_n850) );
  AO21X1_LVT csr_U1278 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[7]), .A3(
        csr_n827), .Y(csr_n828) );
  AO22X1_LVT csr_U1277 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[7]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[7]), .Y(csr_n829) );
  AO22X1_LVT csr_U1276 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[7]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[7]), .Y(csr_n830) );
  AO22X1_LVT csr_U1275 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[7]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[7]), .Y(csr_n831) );
  MUX21X1_LVT csr_U1274 ( .A1(io_ptw_pmp_4_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n509), .Y(csr_n_GEN_286[9]) );
  AO22X1_LVT csr_U1273 ( .A1(csr_n1128), .A2(csr_wdata_44_), .A3(
        csr_n_T_44[38]), .A4(csr_n494), .Y(csr_N1535) );
  AO22X1_LVT csr_U1272 ( .A1(csr_n1149), .A2(csr_wdata_44_), .A3(
        csr_n_T_52[38]), .A4(csr_n1150), .Y(csr_N1929) );
  OR2X1_LVT csr_U1271 ( .A1(csr_n826), .A2(csr_n1690), .Y(csr_io_rw_rdata[44])
         );
  AOI21X1_LVT csr_U1270 ( .A1(csr_n1507), .A2(io_ptw_pmp_5_cfg_a[1]), .A3(
        csr_n822), .Y(csr_n823) );
  AO22X1_LVT csr_U1269 ( .A1(csr_n1689), .A2(csr_n_T_45_44_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[44]), .Y(csr_n822) );
  AOI22X1_LVT csr_U1268 ( .A1(csr_n1508), .A2(csr_reg_sscratch[44]), .A3(
        csr_n1162), .A4(csr_n1955), .Y(csr_n825) );
  AO22X1_LVT csr_U1267 ( .A1(csr_n1128), .A2(csr_wdata_43_), .A3(
        csr_n_T_44[37]), .A4(csr_n495), .Y(csr_N1534) );
  AO22X1_LVT csr_U1266 ( .A1(csr_n1149), .A2(csr_wdata_43_), .A3(
        csr_n_T_52[37]), .A4(csr_n497), .Y(csr_N1928) );
  NAND3X0_LVT csr_U1265 ( .A1(csr_n481), .A2(csr_n1678), .A3(csr_n821), .Y(
        csr_io_rw_rdata[43]) );
  NAND2X0_LVT csr_U1264 ( .A1(csr_n1162), .A2(csr_n1956), .Y(csr_n818) );
  AOI22X1_LVT csr_U1263 ( .A1(csr_n1689), .A2(csr_n_T_45_43_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_5_cfg_a[0]), .Y(csr_n819) );
  MUX21X1_LVT csr_U1262 ( .A1(io_ptw_pmp_5_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n510), .Y(csr_n_GEN_293[9]) );
  AO22X1_LVT csr_U1261 ( .A1(csr_n1128), .A2(csr_wdata_52_), .A3(
        csr_n_T_44[46]), .A4(csr_n1129), .Y(csr_N1543) );
  AO22X1_LVT csr_U1260 ( .A1(csr_n1149), .A2(csr_wdata_52_), .A3(
        csr_n_T_52[46]), .A4(csr_n1150), .Y(csr_N1937) );
  NAND3X0_LVT csr_U1259 ( .A1(csr_n481), .A2(csr_n1685), .A3(csr_n817), .Y(
        csr_io_rw_rdata[52]) );
  NAND2X0_LVT csr_U1258 ( .A1(csr_n1162), .A2(csr_n1947), .Y(csr_n814) );
  AOI22X1_LVT csr_U1257 ( .A1(csr_n1689), .A2(csr_n_T_45_52_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_6_cfg_a[1]), .Y(csr_n815) );
  AO22X1_LVT csr_U1256 ( .A1(csr_n1128), .A2(csr_wdata_51_), .A3(
        csr_n_T_44[45]), .A4(csr_n1129), .Y(csr_N1542) );
  AO22X1_LVT csr_U1255 ( .A1(csr_n1149), .A2(csr_wdata_51_), .A3(
        csr_n_T_52[45]), .A4(csr_n497), .Y(csr_N1936) );
  NAND3X0_LVT csr_U1254 ( .A1(csr_n481), .A2(csr_n1684), .A3(csr_n813), .Y(
        csr_io_rw_rdata[51]) );
  NAND2X0_LVT csr_U1253 ( .A1(csr_n1162), .A2(csr_n1948), .Y(csr_n810) );
  AOI22X1_LVT csr_U1252 ( .A1(csr_n1689), .A2(csr_n_T_45_51_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_6_cfg_a[0]), .Y(csr_n811) );
  AO22X1_LVT csr_U1251 ( .A1(csr_n1128), .A2(csr_wdata_47_), .A3(
        csr_n_T_44[41]), .A4(csr_n1129), .Y(csr_N1538) );
  AO22X1_LVT csr_U1250 ( .A1(csr_n1149), .A2(csr_wdata_47_), .A3(
        csr_n_T_52[41]), .A4(csr_n497), .Y(csr_N1932) );
  NAND3X0_LVT csr_U1249 ( .A1(csr_n481), .A2(csr_n1680), .A3(csr_n809), .Y(
        csr_io_rw_rdata[47]) );
  NAND2X0_LVT csr_U1248 ( .A1(csr_n1162), .A2(csr_n1952), .Y(csr_n806) );
  AOI22X1_LVT csr_U1247 ( .A1(csr_n1689), .A2(csr_n_T_45_47_), .A3(csr_n1507), 
        .A4(io_ptw_pmp_5_cfg_l), .Y(csr_n807) );
  MUX21X1_LVT csr_U1246 ( .A1(io_ptw_pmp_3_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n508), .Y(csr_n_GEN_279[9]) );
  MUX21X1_LVT csr_U1245 ( .A1(csr_io_pc[36]), .A2(csr_wdata_36_), .S0(csr_n513), .Y(csr_net34772) );
  AO22X1_LVT csr_U1244 ( .A1(csr_n1159), .A2(csr_io_tval[36]), .A3(
        csr_wdata_36_), .A4(csr_n1158), .Y(csr_N1418) );
  AO22X1_LVT csr_U1243 ( .A1(csr_n1152), .A2(csr_io_tval[36]), .A3(
        csr_wdata_36_), .A4(csr_n1151), .Y(csr_N1029) );
  AO22X1_LVT csr_U1242 ( .A1(csr_n_T_52[30]), .A2(csr_n1150), .A3(csr_n1149), 
        .A4(csr_wdata_36_), .Y(csr_N1921) );
  OR2X1_LVT csr_U1241 ( .A1(csr_n805), .A2(csr_n1643), .Y(csr_io_rw_rdata[36])
         );
  NAND4X0_LVT csr_U1240 ( .A1(csr_n804), .A2(csr_n803), .A3(csr_n802), .A4(
        csr_n801), .Y(csr_n805) );
  NAND2X0_LVT csr_U1239 ( .A1(csr_n1162), .A2(csr_n1963), .Y(csr_n801) );
  AOI22X1_LVT csr_U1238 ( .A1(csr_n1153), .A2(csr_n_T_383[36]), .A3(csr_n1160), 
        .A4(csr_n_T_444[36]), .Y(csr_n803) );
  AO22X1_LVT csr_U1237 ( .A1(csr_n1128), .A2(csr_wdata_35_), .A3(
        csr_n_T_44[29]), .A4(csr_n1129), .Y(csr_N1526) );
  MUX21X1_LVT csr_U1236 ( .A1(csr_io_pc[35]), .A2(csr_wdata_35_), .S0(csr_n514), .Y(csr_net34977) );
  MUX21X1_LVT csr_U1235 ( .A1(csr_io_pc[35]), .A2(csr_wdata_35_), .S0(csr_n515), .Y(csr_net35199) );
  AO22X1_LVT csr_U1234 ( .A1(csr_wdata_35_), .A2(csr_n1158), .A3(csr_n1159), 
        .A4(csr_io_tval[35]), .Y(csr_N1417) );
  AO22X1_LVT csr_U1233 ( .A1(csr_wdata_35_), .A2(csr_n1151), .A3(csr_n1152), 
        .A4(csr_io_tval[35]), .Y(csr_N1028) );
  AO22X1_LVT csr_U1232 ( .A1(csr_n1149), .A2(csr_wdata_35_), .A3(
        csr_n_T_52[29]), .A4(csr_n496), .Y(csr_N1920) );
  AO22X1_LVT csr_U1231 ( .A1(csr_n493), .A2(csr_n_T_44[22]), .A3(csr_wdata_28_), .A4(csr_n492), .Y(csr_N1519) );
  MUX21X1_LVT csr_U1230 ( .A1(csr_io_pc[28]), .A2(csr_wdata_28_), .S0(csr_n515), .Y(csr_net35220) );
  AO22X1_LVT csr_U1229 ( .A1(csr_n1159), .A2(csr_io_tval[28]), .A3(
        csr_wdata_28_), .A4(csr_n1158), .Y(csr_N1410) );
  AO22X1_LVT csr_U1228 ( .A1(csr_n1152), .A2(csr_io_tval[28]), .A3(
        csr_wdata_28_), .A4(csr_n1151), .Y(csr_N1021) );
  AO22X1_LVT csr_U1227 ( .A1(csr_n497), .A2(csr_n_T_52[22]), .A3(csr_wdata_28_), .A4(csr_n1149), .Y(csr_N1913) );
  AO22X1_LVT csr_U1226 ( .A1(csr_n495), .A2(csr_n_T_44[21]), .A3(csr_wdata_27_), .A4(csr_n492), .Y(csr_N1518) );
  MUX21X1_LVT csr_U1225 ( .A1(csr_io_pc[27]), .A2(csr_wdata_27_), .S0(csr_n515), .Y(csr_net35223) );
  AO22X1_LVT csr_U1224 ( .A1(csr_n1159), .A2(csr_io_tval[27]), .A3(
        csr_wdata_27_), .A4(csr_n1158), .Y(csr_N1409) );
  AO22X1_LVT csr_U1223 ( .A1(csr_n1152), .A2(csr_io_tval[27]), .A3(
        csr_wdata_27_), .A4(csr_n1151), .Y(csr_N1020) );
  AO22X1_LVT csr_U1222 ( .A1(csr_n1150), .A2(csr_n_T_52[21]), .A3(
        csr_wdata_27_), .A4(csr_n1149), .Y(csr_N1912) );
  NAND4X0_LVT csr_U1221 ( .A1(csr_n800), .A2(csr_n799), .A3(csr_n798), .A4(
        csr_n466), .Y(csr_io_rw_rdata[27]) );
  NOR2X0_LVT csr_U1220 ( .A1(csr_n1615), .A2(csr_n1616), .Y(csr_n798) );
  NOR3X0_LVT csr_U1219 ( .A1(csr_n797), .A2(csr_n796), .A3(csr_n1614), .Y(
        csr_n799) );
  AO22X1_LVT csr_U1218 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[27]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[27]), .Y(csr_n796) );
  NOR4X1_LVT csr_U1217 ( .A1(csr_n1619), .A2(csr_n795), .A3(csr_n794), .A4(
        csr_n1618), .Y(csr_n800) );
  NAND4X0_LVT csr_U1216 ( .A1(csr_n793), .A2(csr_n792), .A3(csr_n791), .A4(
        csr_n790), .Y(csr_n795) );
  NAND2X0_LVT csr_U1215 ( .A1(csr_n1493), .A2(csr_reg_dpc_27_), .Y(csr_n790)
         );
  NAND2X0_LVT csr_U1214 ( .A1(csr_n1507), .A2(io_ptw_pmp_3_cfg_a[0]), .Y(
        csr_n791) );
  AOI21X1_LVT csr_U1213 ( .A1(csr_n_T_45_27_), .A2(csr_n1689), .A3(csr_n1617), 
        .Y(csr_n792) );
  NAND2X0_LVT csr_U1212 ( .A1(csr_n1153), .A2(csr_n_T_383[27]), .Y(csr_n793)
         );
  AO22X1_LVT csr_U1211 ( .A1(csr_n1128), .A2(csr_wdata_31_), .A3(
        csr_n_T_44[25]), .A4(csr_n494), .Y(csr_N1522) );
  AO22X1_LVT csr_U1210 ( .A1(csr_n1158), .A2(csr_wdata_31_), .A3(
        csr_io_tval[31]), .A4(csr_n1159), .Y(csr_N1413) );
  AO22X1_LVT csr_U1209 ( .A1(csr_n1151), .A2(csr_wdata_31_), .A3(
        csr_io_tval[31]), .A4(csr_n1152), .Y(csr_N1024) );
  AO22X1_LVT csr_U1208 ( .A1(csr_n1149), .A2(csr_wdata_31_), .A3(
        csr_n_T_52[25]), .A4(csr_n496), .Y(csr_N1916) );
  AO22X1_LVT csr_U1207 ( .A1(csr_n493), .A2(csr_n_T_44[17]), .A3(csr_wdata_23_), .A4(csr_n492), .Y(csr_N1514) );
  MUX21X1_LVT csr_U1206 ( .A1(csr_io_pc[23]), .A2(csr_wdata_23_), .S0(csr_n514), .Y(csr_net35013) );
  AO21X1_LVT csr_U1205 ( .A1(csr_n1919), .A2(csr_n504), .A3(csr_n376), .Y(
        csr_N1582) );
  AO22X1_LVT csr_U1204 ( .A1(csr_n1152), .A2(csr_io_tval[23]), .A3(
        csr_wdata_23_), .A4(csr_n1151), .Y(csr_N1016) );
  AO22X1_LVT csr_U1203 ( .A1(csr_n1150), .A2(csr_n_T_52[17]), .A3(
        csr_wdata_23_), .A4(csr_n1149), .Y(csr_N1908) );
  NAND2X0_LVT csr_U1202 ( .A1(csr_n1605), .A2(csr_n789), .Y(
        csr_io_rw_rdata[23]) );
  NOR4X1_LVT csr_U1201 ( .A1(csr_n788), .A2(csr_n787), .A3(csr_n786), .A4(
        csr_n1602), .Y(csr_n789) );
  OR3X1_LVT csr_U1200 ( .A1(csr_n785), .A2(csr_n784), .A3(csr_n783), .Y(
        csr_n786) );
  AO22X1_LVT csr_U1199 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[23]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[23]), .Y(csr_n783) );
  NAND4X0_LVT csr_U1198 ( .A1(csr_n782), .A2(csr_n781), .A3(csr_n780), .A4(
        csr_n779), .Y(csr_n785) );
  NAND2X0_LVT csr_U1197 ( .A1(csr_n1510), .A2(csr_reg_dscratch[23]), .Y(
        csr_n779) );
  NAND2X0_LVT csr_U1196 ( .A1(csr_n1507), .A2(io_ptw_pmp_2_cfg_l), .Y(csr_n780) );
  AOI21X1_LVT csr_U1195 ( .A1(csr_n_T_45_23_), .A2(csr_n1689), .A3(csr_n1604), 
        .Y(csr_n781) );
  NAND2X0_LVT csr_U1194 ( .A1(csr_n1153), .A2(csr_n_T_383[23]), .Y(csr_n782)
         );
  AO22X1_LVT csr_U1193 ( .A1(csr_n1508), .A2(csr_reg_sscratch[23]), .A3(
        csr_n1162), .A4(csr_io_time[23]), .Y(csr_n787) );
  MUX21X1_LVT csr_U1192 ( .A1(csr_io_pc[9]), .A2(csr_wdata_9_), .S0(csr_n515), 
        .Y(csr_net35277) );
  MUX21X1_LVT csr_U1191 ( .A1(io_ptw_pmp_6_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n511), .Y(csr_n_GEN_300[9]) );
  AO22X1_LVT csr_U1190 ( .A1(csr_n1128), .A2(csr_wdata_60_), .A3(
        csr_n_T_44[54]), .A4(csr_n494), .Y(csr_N1551) );
  AO22X1_LVT csr_U1189 ( .A1(csr_n1149), .A2(csr_wdata_60_), .A3(
        csr_n_T_52[54]), .A4(csr_n496), .Y(csr_N1945) );
  OR2X1_LVT csr_U1188 ( .A1(csr_n778), .A2(csr_n1690), .Y(csr_io_rw_rdata[60])
         );
  AOI21X1_LVT csr_U1187 ( .A1(csr_n1507), .A2(io_ptw_pmp_7_cfg_a[1]), .A3(
        csr_n774), .Y(csr_n775) );
  AO22X1_LVT csr_U1186 ( .A1(csr_n1689), .A2(csr_n_T_45_60_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[60]), .Y(csr_n774) );
  AOI22X1_LVT csr_U1185 ( .A1(csr_n1508), .A2(csr_reg_sscratch[60]), .A3(
        csr_n1162), .A4(csr_n1939), .Y(csr_n777) );
  AO22X1_LVT csr_U1184 ( .A1(csr_n1128), .A2(csr_wdata_59_), .A3(
        csr_n_T_44[53]), .A4(csr_n495), .Y(csr_N1550) );
  AO22X1_LVT csr_U1183 ( .A1(csr_n1149), .A2(csr_wdata_59_), .A3(
        csr_n_T_52[53]), .A4(csr_n496), .Y(csr_N1944) );
  OR2X1_LVT csr_U1182 ( .A1(csr_n773), .A2(csr_n1690), .Y(csr_io_rw_rdata[59])
         );
  OR3X1_LVT csr_U1181 ( .A1(csr_n772), .A2(csr_n771), .A3(csr_n770), .Y(
        csr_n773) );
  AO22X1_LVT csr_U1180 ( .A1(csr_n1508), .A2(csr_reg_sscratch[59]), .A3(
        csr_n1162), .A4(csr_n1940), .Y(csr_n770) );
  NAND2X0_LVT csr_U1179 ( .A1(csr_n1507), .A2(io_ptw_pmp_7_cfg_a[0]), .Y(
        csr_n767) );
  NAND2X0_LVT csr_U1178 ( .A1(csr_n1481), .A2(csr_n_T_366_59_), .Y(csr_n768)
         );
  AOI22X1_LVT csr_U1177 ( .A1(csr_n1689), .A2(csr_n_T_45_59_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[59]), .Y(csr_n769) );
  AO21X1_LVT csr_U1176 ( .A1(csr_n_T_3678_63_), .A2(csr_n504), .A3(csr_n376), 
        .Y(csr_N1622) );
  AO22X1_LVT csr_U1175 ( .A1(csr_n1498), .A2(csr_n1201), .A3(csr_wdata_63_), 
        .A4(csr_n955), .Y(csr_N944) );
  AO22X1_LVT csr_U1174 ( .A1(csr_n1501), .A2(csr_n1201), .A3(csr_wdata_63_), 
        .A4(csr_n923), .Y(csr_N1333) );
  AND2X1_LVT csr_U1173 ( .A1(wb_cause[63]), .A2(csr_n1697), .Y(csr_n1201) );
  OR3X1_LVT csr_U1172 ( .A1(csr_n766), .A2(csr_n1672), .A3(csr_n1690), .Y(
        csr_io_rw_rdata[63]) );
  NAND4X0_LVT csr_U1171 ( .A1(csr_n765), .A2(csr_n764), .A3(csr_n763), .A4(
        csr_n762), .Y(csr_n766) );
  NAND2X0_LVT csr_U1170 ( .A1(csr_n1162), .A2(csr_n1936), .Y(csr_n762) );
  NAND2X0_LVT csr_U1169 ( .A1(csr_n1452), .A2(csr_n_T_3678_63_), .Y(csr_n763)
         );
  AND4X1_LVT csr_U1168 ( .A1(csr_n1155), .A2(csr_n761), .A3(csr_n760), .A4(
        csr_n759), .Y(csr_n764) );
  NAND2X0_LVT csr_U1167 ( .A1(csr_n488), .A2(io_ptw_ptbr_mode[3]), .Y(csr_n759) );
  NAND2X0_LVT csr_U1166 ( .A1(csr_n1507), .A2(io_ptw_pmp_7_cfg_l), .Y(csr_n760) );
  AOI22X1_LVT csr_U1165 ( .A1(csr_n1689), .A2(csr_n_T_45_63_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[63]), .Y(csr_n761) );
  AOI22X1_LVT csr_U1164 ( .A1(csr_n1161), .A2(csr_reg_mcause[63]), .A3(
        csr_n1168), .A4(csr_reg_scause[63]), .Y(csr_n765) );
  AO22X1_LVT csr_U1163 ( .A1(csr_n1129), .A2(csr_n_T_44[8]), .A3(csr_wdata_14_), .A4(csr_n491), .Y(csr_N1505) );
  INVX1_LVT csr_U1162 ( .A(csr_wdata_14_), .Y(csr_n51) );
  MUX21X1_LVT csr_U1161 ( .A1(csr_io_pc[14]), .A2(csr_wdata_14_), .S0(csr_n514), .Y(csr_net35040) );
  AO22X1_LVT csr_U1160 ( .A1(csr_n1159), .A2(csr_io_tval[14]), .A3(
        csr_wdata_14_), .A4(csr_n1158), .Y(csr_N1396) );
  AO22X1_LVT csr_U1159 ( .A1(csr_n1152), .A2(csr_io_tval[14]), .A3(
        csr_wdata_14_), .A4(csr_n1151), .Y(csr_N1007) );
  AO22X1_LVT csr_U1158 ( .A1(csr_n1150), .A2(csr_n_T_52[8]), .A3(csr_wdata_14_), .A4(csr_n1149), .Y(csr_N1899) );
  AO22X1_LVT csr_U1157 ( .A1(csr_n493), .A2(csr_n_T_44[7]), .A3(csr_wdata_13_), 
        .A4(csr_n491), .Y(csr_N1504) );
  AO22X1_LVT csr_U1156 ( .A1(csr_n1159), .A2(csr_io_tval[13]), .A3(
        csr_wdata_13_), .A4(csr_n1158), .Y(csr_N1395) );
  AO22X1_LVT csr_U1155 ( .A1(csr_n1152), .A2(csr_io_tval[13]), .A3(
        csr_wdata_13_), .A4(csr_n1151), .Y(csr_N1006) );
  AO22X1_LVT csr_U1154 ( .A1(csr_n1150), .A2(csr_n_T_52[7]), .A3(csr_wdata_13_), .A4(csr_n1149), .Y(csr_N1898) );
  NAND2X0_LVT csr_U1153 ( .A1(csr_n1928), .A2(csr_n1154), .Y(csr_n1155) );
  NAND2X0_LVT csr_U1152 ( .A1(csr_n1510), .A2(csr_reg_dscratch[13]), .Y(
        csr_n758) );
  AO22X1_LVT csr_U1151 ( .A1(csr_n492), .A2(csr_wdata_55_), .A3(csr_n_T_44[49]), .A4(csr_n494), .Y(csr_N1546) );
  AO22X1_LVT csr_U1150 ( .A1(csr_n1149), .A2(csr_wdata_55_), .A3(
        csr_n_T_52[49]), .A4(csr_n496), .Y(csr_N1940) );
  NAND4X0_LVT csr_U1149 ( .A1(csr_n968), .A2(csr_n757), .A3(csr_n473), .A4(
        csr_n756), .Y(csr_io_rw_rdata[55]) );
  AO22X1_LVT csr_U1148 ( .A1(csr_n1689), .A2(csr_n_T_45_55_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[55]), .Y(csr_n755) );
  AOI22X1_LVT csr_U1147 ( .A1(csr_n1508), .A2(csr_reg_sscratch[55]), .A3(
        csr_n1162), .A4(csr_n1944), .Y(csr_n757) );
  AO22X1_LVT csr_U1146 ( .A1(csr_wdata_39_), .A2(csr_n1158), .A3(
        csr_io_tval[39]), .A4(csr_n1159), .Y(csr_N1421) );
  MUX21X1_LVT csr_U1145 ( .A1(csr_io_pc[39]), .A2(csr_wdata_39_), .S0(csr_n515), .Y(csr_net35187) );
  AO22X1_LVT csr_U1144 ( .A1(csr_wdata_39_), .A2(csr_n1151), .A3(
        csr_io_tval[39]), .A4(csr_n1152), .Y(csr_N1032) );
  AO22X1_LVT csr_U1143 ( .A1(csr_n492), .A2(csr_wdata_39_), .A3(csr_n_T_44[33]), .A4(csr_n495), .Y(csr_N1530) );
  AO22X1_LVT csr_U1142 ( .A1(csr_n1149), .A2(csr_wdata_39_), .A3(
        csr_n_T_52[33]), .A4(csr_n496), .Y(csr_N1924) );
  OR2X1_LVT csr_U1141 ( .A1(csr_n754), .A2(csr_n1690), .Y(csr_io_rw_rdata[39])
         );
  AOI21X1_LVT csr_U1140 ( .A1(csr_n1507), .A2(io_ptw_pmp_4_cfg_l), .A3(
        csr_n750), .Y(csr_n751) );
  AO22X1_LVT csr_U1139 ( .A1(csr_n1689), .A2(csr_n_T_45_39_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[39]), .Y(csr_n750) );
  AOI22X1_LVT csr_U1138 ( .A1(csr_n1508), .A2(csr_reg_sscratch[39]), .A3(
        csr_n1162), .A4(csr_n1960), .Y(csr_n753) );
  NAND3X0_LVT csr_U1137 ( .A1(csr_n748), .A2(csr_n747), .A3(csr_n746), .Y(
        csr_n749) );
  NAND2X0_LVT csr_U1136 ( .A1(csr_n_T_383[39]), .A2(csr_n1153), .Y(csr_n746)
         );
  AOI21X1_LVT csr_U1135 ( .A1(csr_n1493), .A2(csr_reg_dpc_39_), .A3(csr_n1649), 
        .Y(csr_n747) );
  NAND2X0_LVT csr_U1134 ( .A1(csr_n_T_444[39]), .A2(csr_n1160), .Y(csr_n748)
         );
  MUX21X1_LVT csr_U1133 ( .A1(csr_io_pc[9]), .A2(csr_wdata_9_), .S0(csr_n513), 
        .Y(csr_net34853) );
  MUX21X1_LVT csr_U1132 ( .A1(io_ptw_pmp_1_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n506), .Y(csr_n_GEN_265[9]) );
  NAND3X0_LVT csr_U1131 ( .A1(csr_n463), .A2(io_ptw_pmp_2_cfg_l), .A3(
        io_ptw_pmp_2_cfg_a[0]), .Y(csr_n744) );
  AO22X1_LVT csr_U1130 ( .A1(csr_n1158), .A2(csr_wdata_9_), .A3(csr_io_tval[9]), .A4(csr_n1159), .Y(csr_N1391) );
  AO22X1_LVT csr_U1129 ( .A1(csr_n1151), .A2(csr_wdata_9_), .A3(csr_io_tval[9]), .A4(csr_n1152), .Y(csr_N1002) );
  AO22X1_LVT csr_U1128 ( .A1(csr_n498), .A2(csr_n_T_52[3]), .A3(csr_wdata_9_), 
        .A4(csr_n1149), .Y(csr_N1894) );
  NAND2X0_LVT csr_U1127 ( .A1(csr_n503), .A2(csr_n743), .Y(csr_n879) );
  NAND3X0_LVT csr_U1126 ( .A1(csr_n741), .A2(csr_n740), .A3(csr_n739), .Y(
        csr_io_rw_rdata[9]) );
  NOR4X1_LVT csr_U1125 ( .A1(csr_n738), .A2(csr_n737), .A3(csr_n736), .A4(
        csr_n735), .Y(csr_n739) );
  AO22X1_LVT csr_U1124 ( .A1(csr_n1508), .A2(csr_reg_sscratch[9]), .A3(
        csr_n1506), .A4(csr_reg_sepc_9_), .Y(csr_n735) );
  AO22X1_LVT csr_U1123 ( .A1(csr_n1160), .A2(csr_n_T_444[9]), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_9_), .Y(csr_n737) );
  AO22X1_LVT csr_U1122 ( .A1(csr_n1485), .A2(csr_reg_mscratch[9]), .A3(
        csr_n1489), .A4(csr_reg_mepc_9_), .Y(csr_n738) );
  AND4X1_LVT csr_U1121 ( .A1(csr_n734), .A2(csr_n733), .A3(csr_n732), .A4(
        csr_n731), .Y(csr_n740) );
  NAND2X0_LVT csr_U1120 ( .A1(io_ptw_pmp_1_addr[9]), .A2(csr_n1496), .Y(
        csr_n731) );
  NAND2X0_LVT csr_U1119 ( .A1(csr_read_mideleg_9_), .A2(csr_n730), .Y(csr_n732) );
  NAND3X0_LVT csr_U1118 ( .A1(csr_n742), .A2(csr_n1553), .A3(csr_n729), .Y(
        csr_n730) );
  NAND2X0_LVT csr_U1117 ( .A1(csr_n1136), .A2(csr_n1475), .Y(csr_n729) );
  NAND2X0_LVT csr_U1116 ( .A1(csr_reg_mie_9_), .A2(csr_n1503), .Y(csr_n742) );
  AND2X1_LVT csr_U1115 ( .A1(csr_n1504), .A2(csr_n1515), .Y(csr_n1503) );
  AOI22X1_LVT csr_U1114 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[9]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[9]), .Y(csr_n734) );
  NOR4X1_LVT csr_U1113 ( .A1(csr_n728), .A2(csr_n727), .A3(csr_n726), .A4(
        csr_n725), .Y(csr_n741) );
  AO22X1_LVT csr_U1112 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[9]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[9]), .Y(csr_n725) );
  NAND4X0_LVT csr_U1111 ( .A1(csr_n724), .A2(csr_n723), .A3(csr_n722), .A4(
        csr_n721), .Y(csr_n726) );
  NAND2X0_LVT csr_U1110 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[9]), .Y(
        csr_n721) );
  NAND2X0_LVT csr_U1109 ( .A1(csr_reg_stvec_9_), .A2(csr_n1487), .Y(csr_n722)
         );
  AND3X1_LVT csr_U1108 ( .A1(csr_n720), .A2(csr_n719), .A3(csr_n718), .Y(
        csr_n723) );
  OA21X1_LVT csr_U1107 ( .A1(csr_n1912), .A2(csr_n866), .A3(csr_n717), .Y(
        csr_n718) );
  AOI22X1_LVT csr_U1106 ( .A1(csr_n1689), .A2(csr_n_T_45_9_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[9]), .Y(csr_n717) );
  NAND3X0_LVT csr_U1105 ( .A1(csr_n716), .A2(csr_n942), .A3(csr_n715), .Y(
        csr_n866) );
  AND4X1_LVT csr_U1104 ( .A1(csr_n1513), .A2(csr_io_rw_addr[7]), .A3(
        csr_io_rw_addr[6]), .A4(csr_n1522), .Y(csr_n715) );
  AND2X1_LVT csr_U1103 ( .A1(csr_io_rw_addr[10]), .A2(csr_io_rw_addr[9]), .Y(
        csr_n942) );
  AOI22X1_LVT csr_U1102 ( .A1(csr_n1493), .A2(csr_reg_dpc_9_), .A3(csr_n1488), 
        .A4(io_ptw_ptbr_ppn[9]), .Y(csr_n719) );
  NAND2X0_LVT csr_U1101 ( .A1(csr_n1507), .A2(io_ptw_pmp_1_cfg_w), .Y(csr_n720) );
  NAND2X0_LVT csr_U1100 ( .A1(io_ptw_pmp_7_addr[9]), .A2(csr_n1479), .Y(
        csr_n724) );
  AO22X1_LVT csr_U1099 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[9]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[9]), .Y(csr_n727) );
  AO22X1_LVT csr_U1098 ( .A1(csr_n1502), .A2(csr_reg_mie_9_), .A3(csr_n1162), 
        .A4(csr_io_time[9]), .Y(csr_n728) );
  AO22X1_LVT csr_U1097 ( .A1(csr_n1474), .A2(csr_n714), .A3(csr_n_T_3694_9_), 
        .A4(csr_n713), .Y(csr_n200) );
  NAND2X0_LVT csr_U1096 ( .A1(csr_n1474), .A2(csr_n1908), .Y(csr_n713) );
  AND2X1_LVT csr_U1095 ( .A1(io_imem_sfence_bits_addr[9]), .A2(csr_n516), .Y(
        csr_n714) );
  INVX1_LVT csr_U1094 ( .A(csr_n1474), .Y(csr_n1899) );
  INVX1_LVT csr_U1093 ( .A(csr_n1475), .Y(csr_n1898) );
  AND2X1_LVT csr_U1092 ( .A1(csr_n1509), .A2(csr_n1505), .Y(csr_n1475) );
  AO22X1_LVT csr_U1091 ( .A1(csr_n712), .A2(csr_n711), .A3(csr_wdata_1_), .A4(
        csr_n491), .Y(csr_N1429) );
  AO21X1_LVT csr_U1090 ( .A1(csr_n_T_45_0_), .A2(csr_io_retire), .A3(
        csr_n_T_45_1_), .Y(csr_n711) );
  OA22X1_LVT csr_U1089 ( .A1(csr_n_T_389_1), .A2(csr_n935), .A3(csr_n934), 
        .A4(csr_n710), .Y(csr_n2155) );
  MUX21X1_LVT csr_U1088 ( .A1(csr_n709), .A2(io_ptw_status_prv[1]), .S0(
        csr_n1449), .Y(csr_n710) );
  AND2X1_LVT csr_U1087 ( .A1(csr_wdata_0_), .A2(csr_wdata_1_), .Y(csr_n709) );
  NAND2X0_LVT csr_U1086 ( .A1(csr_n935), .A2(csr_n590), .Y(csr_n934) );
  OR2X1_LVT csr_U1085 ( .A1(csr_n932), .A2(csr_N467), .Y(csr_n935) );
  INVX1_LVT csr_U1084 ( .A(csr_n1449), .Y(csr_n932) );
  NAND2X0_LVT csr_U1083 ( .A1(csr_n504), .A2(csr_n1495), .Y(csr_n1449) );
  NAND2X0_LVT csr_U1082 ( .A1(csr_n1448), .A2(csr_n590), .Y(csr_N467) );
  NAND3X0_LVT csr_U1081 ( .A1(csr_n1257), .A2(n9516), .A3(csr_n1139), .Y(
        csr_n1448) );
  AND2X1_LVT csr_U1080 ( .A1(csr_n707), .A2(csr_n1226), .Y(csr_n1467) );
  NAND3X0_LVT csr_U1079 ( .A1(csr_n706), .A2(csr_n860), .A3(n9516), .Y(
        csr_n708) );
  NAND2X0_LVT csr_U1078 ( .A1(csr_n1210), .A2(csr_n705), .Y(csr_n706) );
  MUX21X1_LVT csr_U1077 ( .A1(csr_n704), .A2(csr_n703), .S0(
        io_ptw_status_prv[0]), .Y(csr_n705) );
  MUX21X1_LVT csr_U1076 ( .A1(csr_n_T_1155_1_), .A2(csr_n_T_1155_3), .S0(
        io_ptw_status_prv[1]), .Y(csr_n703) );
  AND2X1_LVT csr_U1075 ( .A1(csr_n381), .A2(csr_n_T_1155_0_), .Y(csr_n704) );
  AO22X1_LVT csr_U1074 ( .A1(csr_wdata_1_), .A2(csr_n1158), .A3(csr_io_tval[1]), .A4(csr_n1159), .Y(csr_N1383) );
  AO22X1_LVT csr_U1073 ( .A1(csr_wdata_1_), .A2(csr_n1151), .A3(csr_io_tval[1]), .A4(csr_n1152), .Y(csr_N994) );
  AO22X1_LVT csr_U1072 ( .A1(csr_n1933), .A2(csr_n883), .A3(csr_wdata_1_), 
        .A4(csr_n949), .Y(csr_n1062) );
  INVX1_LVT csr_U1071 ( .A(csr_n917), .Y(csr_n883) );
  INVX1_LVT csr_U1070 ( .A(csr_N290), .Y(csr_n1443) );
  NAND2X0_LVT csr_U1069 ( .A1(csr_n500), .A2(csr_n590), .Y(csr_n917) );
  NAND2X0_LVT csr_U1068 ( .A1(csr_n590), .A2(csr_n702), .Y(csr_N290) );
  NAND2X0_LVT csr_U1067 ( .A1(csr_n503), .A2(csr_n1154), .Y(csr_n702) );
  AO22X1_LVT csr_U1066 ( .A1(csr_n1498), .A2(csr_n1209), .A3(csr_wdata_1_), 
        .A4(csr_n955), .Y(csr_N882) );
  INVX1_LVT csr_U1065 ( .A(csr_n701), .Y(csr_n955) );
  AO222X1_LVT csr_U1064 ( .A1(csr_n700), .A2(csr_n699), .A3(csr_wdata_1_), 
        .A4(csr_n923), .A5(csr_n1500), .A6(wb_cause[1]), .Y(csr_N1271) );
  OR2X1_LVT csr_U1063 ( .A1(io_ptw_status_prv[1]), .A2(csr_io_rw_addr[0]), .Y(
        csr_n700) );
  AO21X1_LVT csr_U1062 ( .A1(csr_n1164), .A2(io_fpu_fcsr_flags_bits[1]), .A3(
        csr_n698), .Y(csr_n_GEN_345[1]) );
  MUX21X1_LVT csr_U1061 ( .A1(csr_wdata_1_), .A2(csr_read_fcsr_1_), .S0(
        csr_n1163), .Y(csr_n698) );
  AND2X1_LVT csr_U1060 ( .A1(csr_n697), .A2(csr_n589), .Y(csr_n1476) );
  NAND4X0_LVT csr_U1059 ( .A1(csr_n1555), .A2(csr_n696), .A3(csr_n695), .A4(
        csr_n694), .Y(csr_io_rw_rdata[1]) );
  NAND2X0_LVT csr_U1058 ( .A1(csr_n693), .A2(csr_io_status_isa[2]), .Y(
        csr_n694) );
  AO222X1_LVT csr_U1057 ( .A1(csr_n1493), .A2(csr_reg_dpc_1_), .A3(csr_n1506), 
        .A4(csr_reg_sepc_1_), .A5(csr_reg_mepc_1_), .A6(csr_n1489), .Y(
        csr_n693) );
  NOR4X1_LVT csr_U1056 ( .A1(csr_n692), .A2(csr_n1546), .A3(csr_n1547), .A4(
        csr_n1545), .Y(csr_n695) );
  NAND4X0_LVT csr_U1055 ( .A1(csr_n691), .A2(csr_n690), .A3(csr_n689), .A4(
        csr_n688), .Y(csr_n692) );
  NAND2X0_LVT csr_U1054 ( .A1(csr_n1508), .A2(csr_reg_sscratch[1]), .Y(
        csr_n688) );
  NAND2X0_LVT csr_U1053 ( .A1(csr_n1168), .A2(csr_reg_scause[1]), .Y(csr_n689)
         );
  NAND2X0_LVT csr_U1052 ( .A1(csr_n1160), .A2(csr_n_T_444[1]), .Y(csr_n690) );
  NAND2X0_LVT csr_U1051 ( .A1(csr_n1162), .A2(csr_io_time[1]), .Y(csr_n691) );
  NOR4X1_LVT csr_U1050 ( .A1(csr_n687), .A2(csr_n686), .A3(csr_n685), .A4(
        csr_n684), .Y(csr_n696) );
  AND2X1_LVT csr_U1049 ( .A1(csr_n683), .A2(csr_read_mideleg_1), .Y(csr_n684)
         );
  NAND3X0_LVT csr_U1048 ( .A1(csr_n1553), .A2(csr_n1552), .A3(csr_n1692), .Y(
        csr_n683) );
  AO22X1_LVT csr_U1047 ( .A1(csr_n1161), .A2(csr_reg_mcause[1]), .A3(csr_n1484), .A4(csr_read_mcounteren_1_), .Y(csr_n685) );
  AO21X1_LVT csr_U1046 ( .A1(csr_n1153), .A2(csr_n_T_383[1]), .A3(csr_n682), 
        .Y(csr_n686) );
  AO22X1_LVT csr_U1045 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[1]), .A3(
        csr_n1167), .A4(csr_read_fcsr_1_), .Y(csr_n682) );
  NAND4X0_LVT csr_U1044 ( .A1(csr_n681), .A2(csr_n680), .A3(csr_n679), .A4(
        csr_n678), .Y(csr_n687) );
  NAND2X0_LVT csr_U1043 ( .A1(csr_n1507), .A2(io_ptw_pmp_0_cfg_w), .Y(csr_n678) );
  NAND2X0_LVT csr_U1042 ( .A1(csr_n1481), .A2(csr_io_bp_0_control_w), .Y(
        csr_n679) );
  AOI21X1_LVT csr_U1041 ( .A1(csr_n1495), .A2(csr_n_T_389_1), .A3(csr_n677), 
        .Y(csr_n680) );
  AO21X1_LVT csr_U1040 ( .A1(csr_n_T_45_1_), .A2(csr_n1689), .A3(csr_n1554), 
        .Y(csr_n677) );
  NAND2X0_LVT csr_U1039 ( .A1(csr_n1935), .A2(csr_n1154), .Y(csr_n681) );
  NAND2X0_LVT csr_U1038 ( .A1(csr_n676), .A2(csr_n858), .Y(csr_n1553) );
  OR2X1_LVT csr_U1037 ( .A1(csr_n675), .A2(csr_n1543), .Y(csr_io_rw_rdata[5])
         );
  NAND3X0_LVT csr_U1036 ( .A1(csr_n1544), .A2(csr_n674), .A3(csr_n380), .Y(
        csr_n675) );
  AND2X1_LVT csr_U1035 ( .A1(csr_n1487), .A2(csr_n658), .Y(csr_n1478) );
  INVX1_LVT csr_U1034 ( .A(csr_n1477), .Y(csr_n1696) );
  AND2X1_LVT csr_U1033 ( .A1(csr_n1167), .A2(csr_io_rw_addr[1]), .Y(csr_n1477)
         );
  AO22X1_LVT csr_U1032 ( .A1(csr_n495), .A2(csr_n_T_44[6]), .A3(csr_wdata_12_), 
        .A4(csr_n491), .Y(csr_N1503) );
  AND2X1_LVT csr_U1031 ( .A1(csr_n957), .A2(csr_n590), .Y(csr_n961) );
  AND2X1_LVT csr_U1030 ( .A1(csr_n960), .A2(csr_n_T_45_4_), .Y(csr_n1459) );
  AND2X1_LVT csr_U1029 ( .A1(csr_n959), .A2(csr_n_T_45_3_), .Y(csr_n960) );
  AND2X1_LVT csr_U1028 ( .A1(csr_n956), .A2(csr_n_T_45_2_), .Y(csr_n959) );
  AND2X1_LVT csr_U1027 ( .A1(csr_io_retire), .A2(csr_n670), .Y(csr_n956) );
  AND2X1_LVT csr_U1026 ( .A1(csr_n_T_45_1_), .A2(csr_n_T_45_0_), .Y(csr_n670)
         );
  AO22X1_LVT csr_U1025 ( .A1(csr_io_tval[12]), .A2(csr_n1159), .A3(
        csr_wdata_12_), .A4(csr_n1158), .Y(csr_N1394) );
  AO22X1_LVT csr_U1024 ( .A1(csr_io_tval[12]), .A2(csr_n1152), .A3(
        csr_wdata_12_), .A4(csr_n1151), .Y(csr_N1005) );
  AO22X1_LVT csr_U1023 ( .A1(csr_n1150), .A2(csr_n_T_52[6]), .A3(csr_wdata_12_), .A4(csr_n1149), .Y(csr_N1897) );
  INVX1_LVT csr_U1022 ( .A(csr_n1670), .Y(csr_n1083) );
  AND2X1_LVT csr_U1021 ( .A1(n9516), .A2(csr_n_T_389_2), .Y(csr_io_singleStep)
         );
  MUX21X1_LVT csr_U1020 ( .A1(csr_io_pc[2]), .A2(csr_wdata_2_), .S0(csr_n515), 
        .Y(csr_net35298) );
  AO22X1_LVT csr_U1019 ( .A1(csr_io_tval[2]), .A2(csr_n1159), .A3(csr_wdata_2_), .A4(csr_n1158), .Y(csr_N1384) );
  AO22X1_LVT csr_U1018 ( .A1(csr_io_tval[2]), .A2(csr_n1152), .A3(csr_wdata_2_), .A4(csr_n1151), .Y(csr_N995) );
  NAND2X0_LVT csr_U1017 ( .A1(csr_n1161), .A2(csr_n503), .Y(csr_n701) );
  AND2X1_LVT csr_U1016 ( .A1(wb_cause[2]), .A2(csr_n1697), .Y(csr_n1220) );
  NAND2X0_LVT csr_U1015 ( .A1(csr_io_rw_rdata[2]), .A2(csr_n589), .Y(csr_n668)
         );
  NAND2X0_LVT csr_U1014 ( .A1(csr_n1671), .A2(csr_n667), .Y(csr_io_rw_rdata[2]) );
  NOR4X1_LVT csr_U1013 ( .A1(csr_n1660), .A2(csr_n1658), .A3(csr_n666), .A4(
        csr_n665), .Y(csr_n667) );
  OR3X1_LVT csr_U1012 ( .A1(csr_n664), .A2(csr_n663), .A3(csr_n1659), .Y(
        csr_n665) );
  AO22X1_LVT csr_U1011 ( .A1(csr_n1485), .A2(csr_reg_mscratch[2]), .A3(
        csr_read_mcounteren_2_), .A4(csr_n1484), .Y(csr_n663) );
  AND2X1_LVT csr_U1010 ( .A1(csr_n858), .A2(csr_n662), .Y(csr_n1484) );
  AO22X1_LVT csr_U1009 ( .A1(csr_n1153), .A2(csr_n_T_383[2]), .A3(csr_n1161), 
        .A4(csr_reg_mcause[2]), .Y(csr_n664) );
  NAND4X0_LVT csr_U1008 ( .A1(csr_n661), .A2(csr_n660), .A3(csr_n657), .A4(
        csr_n656), .Y(csr_n666) );
  NAND2X0_LVT csr_U1007 ( .A1(io_ptw_pmp_2_addr[2]), .A2(csr_n1492), .Y(
        csr_n656) );
  NAND2X0_LVT csr_U1006 ( .A1(csr_io_status_isa[2]), .A2(csr_n1452), .Y(
        csr_n657) );
  AOI22X1_LVT csr_U1005 ( .A1(csr_n1510), .A2(csr_reg_dscratch[2]), .A3(
        csr_n1493), .A4(csr_reg_dpc_2_), .Y(csr_n660) );
  AOI22X1_LVT csr_U1004 ( .A1(csr_n1160), .A2(csr_n_T_444[2]), .A3(csr_n1168), 
        .A4(csr_reg_scause[2]), .Y(csr_n661) );
  NAND2X0_LVT csr_U1003 ( .A1(csr_n654), .A2(csr_n1514), .Y(csr_n655) );
  NAND3X0_LVT csr_U1002 ( .A1(csr_n1517), .A2(csr_n1518), .A3(
        csr_io_rw_addr[8]), .Y(csr_n654) );
  AO21X1_LVT csr_U1001 ( .A1(csr_n1164), .A2(io_fpu_fcsr_flags_bits[0]), .A3(
        csr_n653), .Y(csr_n_GEN_345[0]) );
  MUX21X1_LVT csr_U1000 ( .A1(csr_wdata_0_), .A2(csr_read_fcsr_0_), .S0(
        csr_n1163), .Y(csr_n653) );
  AND2X1_LVT csr_U999 ( .A1(io_fpu_fcsr_flags_valid), .A2(csr_n1163), .Y(
        csr_n1164) );
  NAND2X0_LVT csr_U998 ( .A1(csr_n1167), .A2(csr_n504), .Y(csr_n1163) );
  NAND3X0_LVT csr_U997 ( .A1(csr_n652), .A2(csr_n651), .A3(csr_n650), .Y(
        csr_io_rw_rdata[0]) );
  NOR4X1_LVT csr_U996 ( .A1(csr_n649), .A2(csr_n648), .A3(csr_n1655), .A4(
        csr_n647), .Y(csr_n651) );
  OR3X1_LVT csr_U995 ( .A1(csr_n646), .A2(csr_n645), .A3(csr_n644), .Y(
        csr_n647) );
  NAND3X0_LVT csr_U994 ( .A1(csr_n643), .A2(csr_n642), .A3(csr_n641), .Y(
        csr_n644) );
  AOI22X1_LVT csr_U993 ( .A1(csr_n1167), .A2(csr_read_fcsr_0_), .A3(csr_n1466), 
        .A4(io_fpu_fcsr_rm[0]), .Y(csr_n641) );
  AND2X1_LVT csr_U992 ( .A1(csr_n1486), .A2(csr_n671), .Y(csr_n1466) );
  AND2X1_LVT csr_U991 ( .A1(csr_n1486), .A2(csr_io_rw_addr[0]), .Y(csr_n1167)
         );
  AND3X1_LVT csr_U990 ( .A1(csr_n1511), .A2(csr_n1514), .A3(csr_n1513), .Y(
        csr_n1486) );
  AOI22X1_LVT csr_U989 ( .A1(csr_n1481), .A2(csr_io_bp_0_control_r), .A3(
        csr_n1490), .A4(csr_io_bp_0_address[0]), .Y(csr_n642) );
  NAND2X0_LVT csr_U988 ( .A1(io_ptw_pmp_0_addr[0]), .A2(csr_n1480), .Y(
        csr_n643) );
  AO21X1_LVT csr_U987 ( .A1(csr_n1161), .A2(csr_reg_mcause[0]), .A3(csr_n639), 
        .Y(csr_n645) );
  AO21X1_LVT csr_U986 ( .A1(csr_read_scounteren_0_), .A2(csr_n1465), .A3(
        csr_n638), .Y(csr_n639) );
  NAND4X0_LVT csr_U985 ( .A1(csr_n637), .A2(csr_n636), .A3(csr_n635), .A4(
        csr_n634), .Y(csr_n638) );
  NAND2X0_LVT csr_U984 ( .A1(csr_n1507), .A2(io_ptw_pmp_0_cfg_r), .Y(csr_n634)
         );
  AOI22X1_LVT csr_U983 ( .A1(csr_n1495), .A2(csr_n_T_389_0), .A3(csr_n488), 
        .A4(io_ptw_ptbr_ppn[0]), .Y(csr_n635) );
  AOI22X1_LVT csr_U982 ( .A1(csr_n1689), .A2(csr_n_T_45_0_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[0]), .Y(csr_n636) );
  NAND2X0_LVT csr_U981 ( .A1(csr_n1520), .A2(csr_n1656), .Y(csr_n637) );
  AND3X1_LVT csr_U980 ( .A1(csr_n1527), .A2(csr_n633), .A3(csr_n662), .Y(
        csr_n1465) );
  AO22X1_LVT csr_U979 ( .A1(csr_n1153), .A2(csr_n_T_383[0]), .A3(csr_n1452), 
        .A4(csr_io_status_isa_0_), .Y(csr_n646) );
  AND2X1_LVT csr_U978 ( .A1(csr_n858), .A2(csr_n716), .Y(csr_n1452) );
  AO22X1_LVT csr_U977 ( .A1(csr_n1168), .A2(csr_reg_scause[0]), .A3(csr_n1162), 
        .A4(csr_io_time[0]), .Y(csr_n648) );
  AO22X1_LVT csr_U976 ( .A1(csr_n1160), .A2(csr_n_T_444[0]), .A3(csr_n1497), 
        .A4(csr_n416), .Y(csr_n649) );
  NOR3X0_LVT csr_U975 ( .A1(csr_n1651), .A2(csr_n1654), .A3(csr_n1652), .Y(
        csr_n652) );
  MUX21X1_LVT csr_U974 ( .A1(csr_io_pc[15]), .A2(csr_wdata_15_), .S0(csr_n514), 
        .Y(csr_net35037) );
  MUX21X1_LVT csr_U973 ( .A1(csr_io_pc[15]), .A2(csr_wdata_15_), .S0(csr_n515), 
        .Y(csr_net35259) );
  AO22X1_LVT csr_U972 ( .A1(csr_n1159), .A2(csr_io_tval[15]), .A3(
        csr_wdata_15_), .A4(csr_n1158), .Y(csr_N1397) );
  AO22X1_LVT csr_U971 ( .A1(csr_n1152), .A2(csr_io_tval[15]), .A3(
        csr_wdata_15_), .A4(csr_n1151), .Y(csr_N1008) );
  AO22X1_LVT csr_U970 ( .A1(csr_n1150), .A2(csr_n_T_52[9]), .A3(csr_wdata_15_), 
        .A4(csr_n1149), .Y(csr_N1900) );
  NAND2X0_LVT csr_U969 ( .A1(csr_n1493), .A2(csr_reg_dpc_15_), .Y(csr_n631) );
  NAND2X0_LVT csr_U968 ( .A1(io_ptw_pmp_1_cfg_l), .A2(csr_n1507), .Y(csr_n632)
         );
  AO22X1_LVT csr_U967 ( .A1(csr_n1158), .A2(csr_wdata_11_), .A3(
        csr_io_tval[11]), .A4(csr_n1159), .Y(csr_N1393) );
  AO22X1_LVT csr_U966 ( .A1(csr_n1151), .A2(csr_wdata_11_), .A3(
        csr_io_tval[11]), .A4(csr_n1152), .Y(csr_N1004) );
  AND2X1_LVT csr_U965 ( .A1(csr_n1139), .A2(csr_n590), .Y(csr_n1499) );
  NAND2X0_LVT csr_U964 ( .A1(csr_n504), .A2(csr_n1161), .Y(csr_n1460) );
  AND2X1_LVT csr_U963 ( .A1(csr_n1501), .A2(csr_n1697), .Y(csr_n1500) );
  AND2X1_LVT csr_U962 ( .A1(csr_n1455), .A2(csr_n1139), .Y(csr_n1501) );
  NAND2X0_LVT csr_U961 ( .A1(csr_n504), .A2(csr_n1168), .Y(csr_n1455) );
  AO22X1_LVT csr_U960 ( .A1(csr_n498), .A2(csr_n_T_52[5]), .A3(csr_wdata_11_), 
        .A4(csr_n1149), .Y(csr_N1896) );
  AND2X1_LVT csr_U959 ( .A1(csr_n1142), .A2(csr_io_time[2]), .Y(csr_n1144) );
  NAND3X0_LVT csr_U958 ( .A1(csr_n503), .A2(csr_n672), .A3(csr_n630), .Y(
        csr_n629) );
  INVX1_LVT csr_U957 ( .A(csr_n1674), .Y(csr_n672) );
  NAND3X0_LVT csr_U956 ( .A1(csr_n628), .A2(csr_n627), .A3(csr_n626), .Y(
        csr_io_rw_rdata[11]) );
  NOR4X1_LVT csr_U955 ( .A1(csr_n625), .A2(csr_n624), .A3(csr_n623), .A4(
        csr_n622), .Y(csr_n626) );
  AO22X1_LVT csr_U954 ( .A1(csr_n1506), .A2(csr_reg_sepc_11_), .A3(csr_n1502), 
        .A4(csr_reg_mie_11_), .Y(csr_n622) );
  AND2X1_LVT csr_U953 ( .A1(csr_n1509), .A2(csr_n857), .Y(csr_n1168) );
  AO22X1_LVT csr_U952 ( .A1(csr_n1160), .A2(csr_n_T_444[11]), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_11_), .Y(csr_n624) );
  AO22X1_LVT csr_U951 ( .A1(csr_n1485), .A2(csr_reg_mscratch[11]), .A3(
        csr_n1489), .A4(csr_reg_mepc_11_), .Y(csr_n625) );
  NOR3X0_LVT csr_U950 ( .A1(csr_n619), .A2(csr_n618), .A3(csr_n617), .Y(
        csr_n627) );
  AO22X1_LVT csr_U949 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[11]), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[11]), .Y(csr_n617) );
  AND2X1_LVT csr_U948 ( .A1(csr_n671), .A2(csr_io_rw_addr[2]), .Y(csr_n662) );
  AO22X1_LVT csr_U947 ( .A1(csr_n1474), .A2(io_interrupts_meip), .A3(csr_n1157), .A4(csr_n_1930_), .Y(csr_n618) );
  NAND2X0_LVT csr_U946 ( .A1(csr_n858), .A2(csr_n1512), .Y(csr_n1041) );
  AND2X1_LVT csr_U945 ( .A1(csr_n1527), .A2(csr_n615), .Y(csr_n858) );
  AND2X1_LVT csr_U944 ( .A1(csr_n620), .A2(csr_n857), .Y(csr_n1161) );
  NOR4X1_LVT csr_U943 ( .A1(csr_n614), .A2(csr_n613), .A3(csr_n612), .A4(
        csr_n611), .Y(csr_n628) );
  AO22X1_LVT csr_U942 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[11]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[11]), .Y(csr_n611) );
  AND3X1_LVT csr_U941 ( .A1(csr_n1518), .A2(csr_io_rw_addr[1]), .A3(
        csr_io_rw_addr[0]), .Y(csr_n676) );
  AO22X1_LVT csr_U940 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[11]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[11]), .Y(csr_n612) );
  AND2X1_LVT csr_U939 ( .A1(csr_n610), .A2(csr_io_rw_addr[2]), .Y(csr_n621) );
  AO22X1_LVT csr_U938 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[11]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[11]), .Y(csr_n613) );
  AND2X1_LVT csr_U937 ( .A1(csr_n630), .A2(csr_io_rw_addr[2]), .Y(csr_n1505)
         );
  NAND4X0_LVT csr_U936 ( .A1(csr_n609), .A2(csr_n608), .A3(csr_n607), .A4(
        csr_n606), .Y(csr_n614) );
  NAND2X0_LVT csr_U935 ( .A1(csr_io_bp_0_address[11]), .A2(csr_n1490), .Y(
        csr_n606) );
  AND2X1_LVT csr_U934 ( .A1(csr_n671), .A2(csr_n1518), .Y(csr_n857) );
  AND2X1_LVT csr_U933 ( .A1(csr_n1526), .A2(csr_io_rw_addr[10]), .Y(csr_n640)
         );
  NAND2X0_LVT csr_U932 ( .A1(csr_reg_stvec_11_), .A2(csr_n1487), .Y(csr_n607)
         );
  AND3X1_LVT csr_U931 ( .A1(csr_n604), .A2(csr_n603), .A3(csr_n602), .Y(
        csr_n608) );
  AOI22X1_LVT csr_U930 ( .A1(csr_n1493), .A2(csr_reg_dpc_11_), .A3(csr_n488), 
        .A4(io_ptw_ptbr_ppn[11]), .Y(csr_n602) );
  NAND4X0_LVT csr_U929 ( .A1(csr_n1513), .A2(csr_io_rw_addr[7]), .A3(csr_n1522), .A4(csr_n445), .Y(csr_n601) );
  AOI22X1_LVT csr_U928 ( .A1(csr_n1689), .A2(csr_n_T_45_11_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[11]), .Y(csr_n603) );
  NAND2X0_LVT csr_U927 ( .A1(io_ptw_pmp_1_cfg_a[0]), .A2(csr_n1507), .Y(
        csr_n604) );
  NAND2X0_LVT csr_U926 ( .A1(csr_n1162), .A2(csr_io_time[11]), .Y(csr_n609) );
  OA21X1_LVT csr_U925 ( .A1(csr_n1918), .A2(csr_n599), .A3(csr_n590), .Y(
        csr_N1693) );
  AND3X1_LVT csr_U924 ( .A1(csr_n1134), .A2(csr_io_rw_addr[9]), .A3(csr_n1519), 
        .Y(csr_n599) );
  OR2X1_LVT csr_U923 ( .A1(wb_ctrl_csr[1]), .A2(wb_ctrl_csr[0]), .Y(csr_n597)
         );
  AND2X1_LVT csr_U922 ( .A1(csr_n1519), .A2(csr_io_rw_addr[0]), .Y(csr_n610)
         );
  AND2X1_LVT csr_U921 ( .A1(csr_n1520), .A2(csr_io_rw_addr[1]), .Y(csr_n671)
         );
  AND4X1_LVT csr_U920 ( .A1(csr_n615), .A2(csr_io_rw_addr[11]), .A3(
        csr_io_rw_addr[8]), .A4(csr_n1514), .Y(csr_n596) );
  AND2X1_LVT csr_U919 ( .A1(csr_n1516), .A2(csr_io_rw_addr[9]), .Y(csr_n615)
         );
  AND3X1_LVT csr_U918 ( .A1(csr_n1557), .A2(csr_n1529), .A3(csr_n595), .Y(
        csr_n1511) );
  NOR2X0_LVT csr_U917 ( .A1(csr_io_rw_addr[8]), .A2(csr_n605), .Y(csr_n595) );
  INVX1_LVT csr_U916 ( .A(csr_io_rw_addr[6]), .Y(csr_n1516) );
  INVX1_LVT csr_U915 ( .A(csr_io_rw_addr[5]), .Y(csr_n1517) );
  NAND2X0_LVT csr_U914 ( .A1(csr_read_mideleg_5), .A2(csr_n1539), .Y(csr_n487)
         );
  NAND3X0_LVT csr_U913 ( .A1(csr_n388), .A2(csr_n469), .A3(csr_n486), .Y(
        csr_n1540) );
  NAND2X0_LVT csr_U912 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[5]), .Y(
        csr_n486) );
  NAND3X0_LVT csr_U911 ( .A1(csr_n480), .A2(csr_n484), .A3(csr_n485), .Y(
        csr_n1627) );
  NAND2X0_LVT csr_U910 ( .A1(csr_n1489), .A2(csr_reg_mepc_30_), .Y(csr_n485)
         );
  NAND3X0_LVT csr_U909 ( .A1(csr_n382), .A2(csr_n471), .A3(csr_n483), .Y(
        csr_n1669) );
  NAND2X0_LVT csr_U908 ( .A1(csr_reg_stvec_2_), .A2(csr_n1478), .Y(csr_n483)
         );
  NAND3X0_LVT csr_U907 ( .A1(csr_n479), .A2(csr_n481), .A3(csr_n482), .Y(
        csr_n1679) );
  NAND2X0_LVT csr_U906 ( .A1(csr_n1508), .A2(csr_reg_sscratch[46]), .Y(
        csr_n482) );
  AND3X1_LVT csr_U905 ( .A1(csr_n384), .A2(csr_n379), .A3(csr_n476), .Y(
        csr_n674) );
  AND2X1_LVT csr_U904 ( .A1(csr_n1510), .A2(csr_reg_dscratch[46]), .Y(csr_n998) );
  AND2X1_LVT csr_U903 ( .A1(csr_n1689), .A2(csr_n_T_45_41_), .Y(csr_n1009) );
  AND2X1_LVT csr_U902 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[37]), .Y(
        csr_n1644) );
  NAND2X0_LVT csr_U901 ( .A1(csr_n1507), .A2(io_ptw_pmp_4_cfg_a[1]), .Y(
        csr_n802) );
  AND2X1_LVT csr_U900 ( .A1(csr_n1489), .A2(csr_reg_mepc_34_), .Y(csr_n1634)
         );
  AND2X1_LVT csr_U899 ( .A1(csr_n1489), .A2(csr_reg_mepc_32_), .Y(csr_n1631)
         );
  NAND2X0_LVT csr_U898 ( .A1(csr_n1485), .A2(csr_reg_mscratch[30]), .Y(
        csr_n1040) );
  AND2X1_LVT csr_U897 ( .A1(csr_n1489), .A2(csr_reg_mepc_29_), .Y(csr_n1049)
         );
  AND2X1_LVT csr_U896 ( .A1(csr_n1160), .A2(csr_n_T_444[27]), .Y(csr_n794) );
  NAND2X0_LVT csr_U895 ( .A1(csr_n1497), .A2(csr_reg_mtvec_24_), .Y(csr_n1061)
         );
  AND2X1_LVT csr_U894 ( .A1(csr_n1452), .A2(csr_n1919), .Y(csr_n784) );
  NAND2X0_LVT csr_U893 ( .A1(csr_n1153), .A2(csr_n_T_383[20]), .Y(csr_n1072)
         );
  AND2X1_LVT csr_U892 ( .A1(csr_n1485), .A2(csr_reg_mscratch[19]), .Y(
        csr_n1081) );
  AND2X1_LVT csr_U891 ( .A1(csr_n1497), .A2(csr_reg_mtvec_18_), .Y(csr_n1106)
         );
  AND2X1_LVT csr_U890 ( .A1(csr_n1493), .A2(csr_reg_dpc_17_), .Y(csr_n1578) );
  NAND2X0_LVT csr_U889 ( .A1(csr_n1160), .A2(csr_n_T_444[16]), .Y(csr_n1123)
         );
  AND2X1_LVT csr_U888 ( .A1(csr_n1153), .A2(csr_n_T_383[11]), .Y(csr_n619) );
  NAND2X0_LVT csr_U887 ( .A1(csr_n1153), .A2(csr_n_T_383[9]), .Y(csr_n733) );
  AND2X1_LVT csr_U886 ( .A1(csr_n1477), .A2(io_fpu_fcsr_rm[2]), .Y(csr_n827)
         );
  NAND2X0_LVT csr_U885 ( .A1(csr_n1485), .A2(csr_reg_mscratch[62]), .Y(
        csr_n963) );
  NAND2X0_LVT csr_U884 ( .A1(csr_n1485), .A2(csr_reg_mscratch[61]), .Y(
        csr_n966) );
  NAND2X0_LVT csr_U883 ( .A1(csr_n1485), .A2(csr_reg_mscratch[60]), .Y(
        csr_n776) );
  AND2X1_LVT csr_U882 ( .A1(csr_n1485), .A2(csr_reg_mscratch[59]), .Y(csr_n771) );
  NAND2X0_LVT csr_U881 ( .A1(csr_n1162), .A2(csr_n1941), .Y(csr_n970) );
  NAND2X0_LVT csr_U880 ( .A1(csr_n1162), .A2(csr_n1942), .Y(csr_n972) );
  NAND2X0_LVT csr_U879 ( .A1(csr_n1485), .A2(csr_reg_mscratch[56]), .Y(
        csr_n975) );
  NAND2X0_LVT csr_U878 ( .A1(csr_n1485), .A2(csr_reg_mscratch[55]), .Y(
        csr_n756) );
  NAND2X0_LVT csr_U877 ( .A1(csr_n1485), .A2(csr_reg_mscratch[54]), .Y(
        csr_n978) );
  NAND2X0_LVT csr_U876 ( .A1(csr_n1485), .A2(csr_reg_mscratch[53]), .Y(
        csr_n982) );
  NAND2X0_LVT csr_U875 ( .A1(csr_n1485), .A2(csr_reg_mscratch[52]), .Y(
        csr_n816) );
  NAND2X0_LVT csr_U874 ( .A1(csr_n1508), .A2(csr_reg_sscratch[51]), .Y(
        csr_n812) );
  NAND2X0_LVT csr_U873 ( .A1(csr_n1508), .A2(csr_reg_sscratch[50]), .Y(
        csr_n987) );
  NAND2X0_LVT csr_U872 ( .A1(csr_n1485), .A2(csr_reg_mscratch[49]), .Y(
        csr_n991) );
  NAND2X0_LVT csr_U871 ( .A1(csr_n1508), .A2(csr_reg_sscratch[48]), .Y(
        csr_n995) );
  NAND2X0_LVT csr_U870 ( .A1(csr_n1485), .A2(csr_reg_mscratch[47]), .Y(
        csr_n808) );
  NAND2X0_LVT csr_U869 ( .A1(csr_n1485), .A2(csr_reg_mscratch[45]), .Y(
        csr_n1000) );
  NAND2X0_LVT csr_U868 ( .A1(csr_n1485), .A2(csr_reg_mscratch[44]), .Y(
        csr_n824) );
  NAND2X0_LVT csr_U867 ( .A1(csr_n1508), .A2(csr_reg_sscratch[43]), .Y(
        csr_n820) );
  NAND2X0_LVT csr_U866 ( .A1(csr_n1508), .A2(csr_reg_sscratch[42]), .Y(
        csr_n1005) );
  AND2X1_LVT csr_U865 ( .A1(csr_n1485), .A2(csr_reg_mscratch[41]), .Y(
        csr_n1008) );
  NAND2X0_LVT csr_U864 ( .A1(csr_n1485), .A2(csr_reg_mscratch[40]), .Y(
        csr_n1013) );
  NAND2X0_LVT csr_U863 ( .A1(csr_n1485), .A2(csr_reg_mscratch[39]), .Y(
        csr_n752) );
  AND2X1_LVT csr_U862 ( .A1(csr_n1485), .A2(csr_reg_mscratch[37]), .Y(
        csr_n1645) );
  NAND2X0_LVT csr_U861 ( .A1(csr_n1506), .A2(csr_reg_sepc_36_), .Y(csr_n804)
         );
  AND2X1_LVT csr_U860 ( .A1(csr_n1493), .A2(csr_reg_dpc_34_), .Y(csr_n1636) );
  AND2X1_LVT csr_U859 ( .A1(csr_n1510), .A2(csr_reg_dscratch[32]), .Y(
        csr_n1629) );
  AND2X1_LVT csr_U858 ( .A1(csr_n1160), .A2(csr_n_T_444[29]), .Y(csr_n1045) );
  AND2X1_LVT csr_U857 ( .A1(csr_n1162), .A2(csr_io_time[27]), .Y(csr_n797) );
  NAND2X0_LVT csr_U856 ( .A1(csr_n1160), .A2(csr_n_T_444[24]), .Y(csr_n1060)
         );
  AND2X1_LVT csr_U855 ( .A1(csr_n1489), .A2(csr_reg_mepc_23_), .Y(csr_n788) );
  NAND2X0_LVT csr_U854 ( .A1(csr_n1508), .A2(csr_reg_sscratch[20]), .Y(
        csr_n1073) );
  AND2X1_LVT csr_U853 ( .A1(csr_n1162), .A2(csr_io_time[19]), .Y(csr_n1092) );
  AND2X1_LVT csr_U852 ( .A1(csr_n1160), .A2(csr_n_T_444[18]), .Y(csr_n1105) );
  AND2X1_LVT csr_U851 ( .A1(csr_n1160), .A2(csr_n_T_444[17]), .Y(csr_n1577) );
  NAND2X0_LVT csr_U850 ( .A1(csr_n1162), .A2(csr_io_time[16]), .Y(csr_n1124)
         );
  AND2X1_LVT csr_U849 ( .A1(csr_n1508), .A2(csr_reg_sscratch[11]), .Y(csr_n623) );
  AND2X1_LVT csr_U848 ( .A1(csr_n1474), .A2(csr_n1136), .Y(csr_n736) );
  AND2X1_LVT csr_U847 ( .A1(csr_n1508), .A2(csr_reg_sscratch[7]), .Y(csr_n832)
         );
  AND2X1_LVT csr_U846 ( .A1(csr_wdata_4_), .A2(csr_n923), .Y(csr_N1274) );
  AND3X1_LVT csr_U845 ( .A1(csr_n1220), .A2(csr_n954), .A3(csr_n1209), .Y(
        csr_n707) );
  NAND3X0_LVT csr_U844 ( .A1(csr_n752), .A2(csr_n751), .A3(csr_n753), .Y(
        csr_n754) );
  NAND3X0_LVT csr_U843 ( .A1(csr_n768), .A2(csr_n767), .A3(csr_n769), .Y(
        csr_n772) );
  NAND3X0_LVT csr_U842 ( .A1(csr_n776), .A2(csr_n775), .A3(csr_n777), .Y(
        csr_n778) );
  AND3X1_LVT csr_U841 ( .A1(csr_n807), .A2(csr_n806), .A3(csr_n808), .Y(
        csr_n809) );
  AND3X1_LVT csr_U840 ( .A1(csr_n811), .A2(csr_n810), .A3(csr_n812), .Y(
        csr_n813) );
  AND3X1_LVT csr_U839 ( .A1(csr_n815), .A2(csr_n814), .A3(csr_n816), .Y(
        csr_n817) );
  AND3X1_LVT csr_U838 ( .A1(csr_n819), .A2(csr_n818), .A3(csr_n820), .Y(
        csr_n821) );
  NAND3X0_LVT csr_U837 ( .A1(csr_n824), .A2(csr_n823), .A3(csr_n825), .Y(
        csr_n826) );
  NAND3X0_LVT csr_U836 ( .A1(csr_n963), .A2(csr_n962), .A3(csr_n964), .Y(
        csr_n965) );
  AND3X1_LVT csr_U835 ( .A1(csr_n974), .A2(csr_n973), .A3(csr_n975), .Y(
        csr_n976) );
  NAND3X0_LVT csr_U834 ( .A1(csr_n978), .A2(csr_n977), .A3(csr_n979), .Y(
        csr_n980) );
  NAND3X0_LVT csr_U833 ( .A1(csr_n982), .A2(csr_n981), .A3(csr_n983), .Y(
        csr_n984) );
  AND3X1_LVT csr_U832 ( .A1(csr_n986), .A2(csr_n985), .A3(csr_n987), .Y(
        csr_n988) );
  AND3X1_LVT csr_U831 ( .A1(csr_n990), .A2(csr_n989), .A3(csr_n991), .Y(
        csr_n992) );
  AND3X1_LVT csr_U830 ( .A1(csr_n994), .A2(csr_n993), .A3(csr_n995), .Y(
        csr_n996) );
  NAND3X0_LVT csr_U829 ( .A1(csr_n1000), .A2(csr_n999), .A3(csr_n1001), .Y(
        csr_n1002) );
  AND3X1_LVT csr_U828 ( .A1(csr_n1004), .A2(csr_n1003), .A3(csr_n1005), .Y(
        csr_n1006) );
  AND3X1_LVT csr_U827 ( .A1(csr_n1012), .A2(csr_n1011), .A3(csr_n1013), .Y(
        csr_n1014) );
  NAND3X0_LVT csr_U826 ( .A1(csr_n1234), .A2(csr_n1233), .A3(csr_n1235), .Y(
        csr_io_evec[6]) );
  NAND3X0_LVT csr_U825 ( .A1(csr_n1241), .A2(csr_n1240), .A3(csr_n1242), .Y(
        csr_io_evec[7]) );
  NAND2X0_LVT csr_U824 ( .A1(csr_n1487), .A2(csr_reg_stvec_30_), .Y(csr_n480)
         );
  NAND2X0_LVT csr_U823 ( .A1(csr_n1689), .A2(csr_n_T_45_46_), .Y(csr_n479) );
  AOI21X1_LVT csr_U822 ( .A1(csr_n1493), .A2(csr_reg_dpc_19_), .A3(csr_n1591), 
        .Y(csr_n478) );
  AOI22X1_LVT csr_U821 ( .A1(csr_n1510), .A2(csr_reg_dscratch[5]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[5]), .Y(csr_n476) );
  AOI21X1_LVT csr_U820 ( .A1(csr_n1507), .A2(io_ptw_pmp_7_cfg_w), .A3(csr_n971), .Y(csr_n475) );
  AOI21X1_LVT csr_U819 ( .A1(csr_n1507), .A2(io_ptw_pmp_7_cfg_x), .A3(csr_n969), .Y(csr_n474) );
  AOI21X1_LVT csr_U818 ( .A1(csr_n1507), .A2(io_ptw_pmp_6_cfg_l), .A3(csr_n755), .Y(csr_n473) );
  AOI22X1_LVT csr_U817 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[2]), .A3(
        csr_n1466), .A4(io_fpu_fcsr_rm[2]), .Y(csr_n471) );
  AOI22X1_LVT csr_U816 ( .A1(csr_n1502), .A2(csr_reg_mie_5_), .A3(csr_n1508), 
        .A4(csr_reg_sscratch[5]), .Y(csr_n469) );
  AOI22X1_LVT csr_U815 ( .A1(csr_n1160), .A2(csr_n_T_444[5]), .A3(csr_n1496), 
        .A4(io_ptw_pmp_1_addr[5]), .Y(csr_n468) );
  AOI22X1_LVT csr_U814 ( .A1(csr_n1689), .A2(csr_n_T_45_61_), .A3(csr_n1510), 
        .A4(csr_reg_dscratch[61]), .Y(csr_n467) );
  AOI22X1_LVT csr_U813 ( .A1(csr_n1508), .A2(csr_reg_sscratch[27]), .A3(
        csr_n1506), .A4(csr_reg_sepc_27_), .Y(csr_n466) );
  AND2X1_LVT csr_U812 ( .A1(csr_n1512), .A2(csr_n1514), .Y(csr_n445) );
  AND2X1_LVT csr_U811 ( .A1(wb_ctrl_csr[0]), .A2(csr_n589), .Y(csr_n444) );
  NBUFFX2_LVT csr_U810 ( .A(csr_n1348), .Y(csr_n499) );
  NBUFFX2_LVT csr_U809 ( .A(csr_n1128), .Y(csr_n492) );
  AOI22X1_LVT csr_U808 ( .A1(csr_n1153), .A2(csr_n_T_383[5]), .A3(
        csr_reg_mtvec_5_), .A4(csr_n1470), .Y(csr_n388) );
  AOI22X1_LVT csr_U807 ( .A1(csr_n1452), .A2(csr_n1923), .A3(csr_reg_mepc_5_), 
        .A4(csr_n1489), .Y(csr_n385) );
  AOI22X1_LVT csr_U806 ( .A1(csr_n1689), .A2(csr_n_T_45_5_), .A3(csr_n1477), 
        .A4(io_fpu_fcsr_rm[0]), .Y(csr_n384) );
  AOI22X1_LVT csr_U805 ( .A1(csr_n1162), .A2(csr_io_time[2]), .A3(csr_n1689), 
        .A4(csr_n_T_45_2_), .Y(csr_n382) );
  AND3X1_LVT csr_U804 ( .A1(csr_n468), .A2(csr_n385), .A3(csr_n487), .Y(
        csr_n380) );
  AOI22X1_LVT csr_U803 ( .A1(csr_n1478), .A2(csr_reg_stvec_5_), .A3(csr_n1162), 
        .A4(csr_io_time[5]), .Y(csr_n379) );
  NOR4X1_LVT csr_U802 ( .A1(csr_n1601), .A2(csr_n1600), .A3(csr_n1599), .A4(
        csr_n1598), .Y(csr_n1605) );
  AND2X1_LVT csr_U801 ( .A1(csr_n1504), .A2(csr_io_rw_addr[9]), .Y(csr_n1502)
         );
  NOR4X1_LVT csr_U800 ( .A1(csr_n1670), .A2(csr_n1669), .A3(csr_n1668), .A4(
        csr_n1667), .Y(csr_n1671) );
  NOR4X1_LVT csr_U799 ( .A1(csr_n1578), .A2(csr_n1577), .A3(csr_n1576), .A4(
        csr_n1575), .Y(csr_n1580) );
  NOR4X1_LVT csr_U798 ( .A1(csr_n1574), .A2(csr_n1573), .A3(csr_n1572), .A4(
        csr_n1571), .Y(csr_n1581) );
  NOR4X1_LVT csr_U797 ( .A1(csr_n1551), .A2(csr_n1550), .A3(csr_n1549), .A4(
        csr_n1548), .Y(csr_n1555) );
  NOR4X1_LVT csr_U796 ( .A1(csr_n1537), .A2(csr_n1536), .A3(csr_n1535), .A4(
        csr_n1534), .Y(csr_n1544) );
  NOR4X1_LVT csr_U795 ( .A1(csr_n1611), .A2(csr_n1610), .A3(csr_n1609), .A4(
        csr_n1608), .Y(csr_n1613) );
  NOR4X1_LVT csr_U794 ( .A1(csr_n1567), .A2(csr_n1566), .A3(csr_n1565), .A4(
        csr_n1564), .Y(csr_n1570) );
  NAND2X0_LVT csr_U793 ( .A1(csr_n1134), .A2(csr_n655), .Y(csr_n1903) );
  NBUFFX2_LVT csr_U792 ( .A(csr_net34920), .Y(csr_n571) );
  NBUFFX2_LVT csr_U791 ( .A(csr_net34935), .Y(csr_n558) );
  NBUFFX2_LVT csr_U790 ( .A(csr_net34885), .Y(csr_n580) );
  NBUFFX2_LVT csr_U789 ( .A(csr_net34935), .Y(csr_n557) );
  NBUFFX2_LVT csr_U788 ( .A(csr_net34722), .Y(csr_n587) );
  AND2X1_LVT csr_U787 ( .A1(csr_n1460), .A2(csr_n1499), .Y(csr_n1498) );
  NBUFFX2_LVT csr_U786 ( .A(csr_net35324), .Y(csr_n520) );
  NBUFFX2_LVT csr_U785 ( .A(csr_net35324), .Y(csr_n517) );
  NBUFFX2_LVT csr_U784 ( .A(csr_net35324), .Y(csr_n519) );
  NBUFFX2_LVT csr_U783 ( .A(csr_net35324), .Y(csr_n518) );
  NBUFFX2_LVT csr_U782 ( .A(csr_net35324), .Y(csr_n521) );
  XOR2X1_LVT csr_U781 ( .A1(csr_n1147), .A2(csr_io_time[5]), .Y(csr_n1148) );
  NOR4X1_LVT csr_U780 ( .A1(csr_wdata_62_), .A2(csr_wdata_61_), .A3(
        csr_wdata_60_), .A4(csr_n1673), .Y(csr_N1426) );
  INVX1_LVT csr_U779 ( .A(csr_io_rw_addr[8]), .Y(csr_n600) );
  AND2X1_LVT csr_U778 ( .A1(csr_n610), .A2(csr_n1518), .Y(csr_n716) );
  AND4X1_LVT csr_U777 ( .A1(csr_n1514), .A2(csr_n1528), .A3(csr_n1513), .A4(
        csr_n1522), .Y(csr_n1527) );
  INVX1_LVT csr_U776 ( .A(csr_io_rw_addr[0]), .Y(csr_n1520) );
  NAND3X0_LVT csr_U775 ( .A1(csr_n1557), .A2(csr_n1529), .A3(csr_n596), .Y(
        csr_n1674) );
  AND3X1_LVT csr_U774 ( .A1(csr_io_rw_addr[10]), .A2(csr_n1523), .A3(csr_n1518), .Y(csr_n1532) );
  NAND2X0_LVT csr_U773 ( .A1(csr_n1903), .A2(csr_n1697), .Y(csr_io_eret) );
  NAND2X0_LVT csr_U772 ( .A1(csr_n504), .A2(csr_n1153), .Y(csr_n1457) );
  NAND2X0_LVT csr_U771 ( .A1(csr_n504), .A2(csr_n1160), .Y(csr_n1456) );
  NAND2X0_LVT csr_U770 ( .A1(csr_n1506), .A2(csr_n504), .Y(csr_n448) );
  NAND2X0_LVT csr_U769 ( .A1(csr_n1489), .A2(csr_n504), .Y(csr_n449) );
  AND2X1_LVT csr_U768 ( .A1(csr_n961), .A2(csr_n_T_45_5_), .Y(csr_n673) );
  NBUFFX2_LVT csr_U767 ( .A(csr_n1129), .Y(csr_n493) );
  NBUFFX2_LVT csr_U766 ( .A(csr_n1129), .Y(csr_n494) );
  NBUFFX2_LVT csr_U765 ( .A(csr_n1129), .Y(csr_n495) );
  NAND2X0_LVT csr_U764 ( .A1(csr_n504), .A2(csr_n1493), .Y(csr_n450) );
  NBUFFX2_LVT csr_U763 ( .A(clock), .Y(csr_n591) );
  AND2X1_LVT csr_U762 ( .A1(csr_n1147), .A2(csr_io_time[5]), .Y(csr_n1445) );
  NBUFFX2_LVT csr_U761 ( .A(csr_n1150), .Y(csr_n496) );
  NBUFFX2_LVT csr_U760 ( .A(csr_n1150), .Y(csr_n497) );
  NBUFFX2_LVT csr_U759 ( .A(csr_n1150), .Y(csr_n498) );
  AND2X1_LVT csr_U758 ( .A1(csr_n744), .A2(csr_n440), .Y(csr_n745) );
  AND2X1_LVT csr_U757 ( .A1(csr_n1507), .A2(csr_n504), .Y(csr_n1463) );
  INVX1_LVT csr_U756 ( .A(csr_io_rw_addr[11]), .Y(csr_n1513) );
  INVX1_LVT csr_U755 ( .A(csr_io_rw_addr[10]), .Y(csr_n1514) );
  AND2X1_LVT csr_U754 ( .A1(csr_n1523), .A2(csr_n1514), .Y(csr_n616) );
  AND2X1_LVT csr_U753 ( .A1(csr_n616), .A2(csr_n1505), .Y(csr_n1491) );
  AND2X1_LVT csr_U752 ( .A1(csr_n616), .A2(csr_n716), .Y(csr_n1496) );
  AND2X1_LVT csr_U751 ( .A1(csr_n671), .A2(csr_n1532), .Y(csr_n1510) );
  NOR2X0_LVT csr_U750 ( .A1(csr_n605), .A2(csr_n601), .Y(csr_n1488) );
  AND2X1_LVT csr_U749 ( .A1(csr_n616), .A2(csr_n621), .Y(csr_n1472) );
  AND2X1_LVT csr_U748 ( .A1(csr_n640), .A2(csr_n857), .Y(csr_n1490) );
  AND2X1_LVT csr_U747 ( .A1(csr_n1509), .A2(csr_n716), .Y(csr_n1506) );
  AND2X1_LVT csr_U746 ( .A1(csr_n620), .A2(csr_n716), .Y(csr_n1489) );
  AND2X1_LVT csr_U745 ( .A1(csr_n1509), .A2(csr_n1512), .Y(csr_n1508) );
  AND2X1_LVT csr_U744 ( .A1(csr_n858), .A2(csr_n621), .Y(csr_n1497) );
  AND2X1_LVT csr_U743 ( .A1(csr_n1509), .A2(csr_n676), .Y(csr_n1160) );
  AND2X1_LVT csr_U742 ( .A1(csr_n630), .A2(csr_n1531), .Y(csr_n1162) );
  AND2X1_LVT csr_U741 ( .A1(csr_n616), .A2(csr_n1512), .Y(csr_n1480) );
  AND2X1_LVT csr_U740 ( .A1(csr_n616), .A2(csr_n676), .Y(csr_n1473) );
  AND2X1_LVT csr_U739 ( .A1(csr_n616), .A2(csr_n857), .Y(csr_n1492) );
  AND2X1_LVT csr_U738 ( .A1(csr_n616), .A2(csr_n662), .Y(csr_n1494) );
  AND2X1_LVT csr_U737 ( .A1(csr_n620), .A2(csr_n1512), .Y(csr_n1485) );
  AND2X1_LVT csr_U736 ( .A1(csr_n610), .A2(csr_n1532), .Y(csr_n1493) );
  AND2X1_LVT csr_U735 ( .A1(csr_n630), .A2(csr_n1532), .Y(csr_n1495) );
  AND2X1_LVT csr_U734 ( .A1(csr_n640), .A2(csr_n716), .Y(csr_n1481) );
  OR2X1_LVT csr_U733 ( .A1(csr_n749), .A2(csr_n1650), .Y(csr_n1690) );
  INVX1_LVT csr_U732 ( .A(csr_n1690), .Y(csr_n481) );
  AND2X1_LVT csr_U731 ( .A1(csr_io_rw_cmd_2_), .A2(csr_n598), .Y(csr_n1134) );
  NAND2X0_LVT csr_U730 ( .A1(csr_n1134), .A2(csr_n600), .Y(csr_n1697) );
  OR2X1_LVT csr_U729 ( .A1(csr_n1918), .A2(io_wfi), .Y(csr_io_csr_stall) );
  INVX1_LVT csr_U728 ( .A(csr_n1220), .Y(csr_n899) );
  OR2X1_LVT csr_U727 ( .A1(csr_n882), .A2(csr_n1903), .Y(csr_n451) );
  INVX1_LVT csr_U726 ( .A(csr_n451), .Y(csr_n502) );
  AND2X1_LVT csr_U725 ( .A1(csr_n1134), .A2(csr_n942), .Y(csr_n1356) );
  INVX1_LVT csr_U724 ( .A(csr_n1355), .Y(csr_n501) );
  INVX1_LVT csr_U723 ( .A(csr_n501), .Y(csr_n500) );
  NAND2X0_LVT csr_U722 ( .A1(csr_io_rw_cmd_2_), .A2(csr_n597), .Y(csr_n387) );
  INVX1_LVT csr_U721 ( .A(csr_n387), .Y(csr_n504) );
  NBUFFX2_LVT csr_U720 ( .A(wb_ctrl_csr[1]), .Y(csr_n589) );
  INVX1_LVT csr_U719 ( .A(csr_n444), .Y(csr_n516) );
  INVX1_LVT csr_U718 ( .A(csr_n1457), .Y(csr_n1151) );
  INVX1_LVT csr_U717 ( .A(csr_n1456), .Y(csr_n1158) );
  AO22X1_LVT csr_U716 ( .A1(io_imem_sfence_bits_addr[1]), .A2(csr_n516), .A3(
        csr_io_rw_rdata[1]), .A4(csr_n1476), .Y(csr_wdata_1_) );
  MUX21X1_LVT csr_U715 ( .A1(csr_n668), .A2(csr_n444), .S0(
        io_imem_sfence_bits_addr[2]), .Y(csr_n1483) );
  INVX1_LVT csr_U714 ( .A(csr_n1483), .Y(csr_wdata_2_) );
  INVX1_LVT csr_U713 ( .A(csr_n449), .Y(csr_n514) );
  NAND2X0_LVT csr_U712 ( .A1(csr_n1479), .A2(csr_n442), .Y(csr_n386) );
  INVX1_LVT csr_U711 ( .A(csr_n450), .Y(csr_n515) );
  NAND2X0_LVT csr_U710 ( .A1(csr_n1496), .A2(csr_n745), .Y(csr_n431) );
  INVX1_LVT csr_U709 ( .A(csr_n448), .Y(csr_n513) );
  INVX1_LVT csr_U708 ( .A(csr_n430), .Y(csr_n505) );
  INVX1_LVT csr_U707 ( .A(csr_n386), .Y(csr_n512) );
  INVX1_LVT csr_U706 ( .A(csr_n435), .Y(csr_n511) );
  INVX1_LVT csr_U705 ( .A(csr_n431), .Y(csr_n506) );
  INVX1_LVT csr_U704 ( .A(csr_n434), .Y(csr_n510) );
  INVX1_LVT csr_U703 ( .A(csr_n432), .Y(csr_n507) );
  INVX1_LVT csr_U702 ( .A(csr_n433), .Y(csr_n509) );
  INVX1_LVT csr_U701 ( .A(csr_n436), .Y(csr_n508) );
  MUX21X1_LVT csr_U700 ( .A1(io_ptw_pmp_0_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n505), .Y(csr_n_GEN_258[9]) );
  MUX21X1_LVT csr_U699 ( .A1(io_ptw_pmp_2_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n507), .Y(csr_n_GEN_272[9]) );
  MUX21X1_LVT csr_U698 ( .A1(io_ptw_pmp_7_addr[9]), .A2(csr_wdata_9_), .S0(
        csr_n512), .Y(csr_n_GEN_307[9]) );
  MUX21X1_LVT csr_U697 ( .A1(io_ptw_pmp_1_addr[3]), .A2(csr_wdata_3_), .S0(
        csr_n506), .Y(csr_n_GEN_265[3]) );
  MUX21X1_LVT csr_U696 ( .A1(csr_io_pc[7]), .A2(csr_wdata_7_), .S0(csr_n514), 
        .Y(csr_net35061) );
  MUX21X1_LVT csr_U695 ( .A1(csr_io_pc[7]), .A2(csr_wdata_7_), .S0(csr_n515), 
        .Y(csr_net35283) );
  MUX21X1_LVT csr_U694 ( .A1(csr_io_pc[7]), .A2(csr_wdata_7_), .S0(csr_n513), 
        .Y(csr_net34859) );
  MUX21X1_LVT csr_U693 ( .A1(csr_io_pc[11]), .A2(csr_wdata_11_), .S0(csr_n515), 
        .Y(csr_net35271) );
  MUX21X1_LVT csr_U692 ( .A1(csr_io_pc[11]), .A2(csr_wdata_11_), .S0(csr_n513), 
        .Y(csr_net34847) );
  INVX1_LVT csr_U691 ( .A(ibuf_io_inst_0_bits_raw[21]), .Y(csr_n1407) );
  INVX1_LVT csr_U690 ( .A(ibuf_io_inst_0_bits_raw[27]), .Y(csr_n1386) );
  OR2X1_LVT csr_U689 ( .A1(csr_n1370), .A2(csr_n1369), .Y(csr_n1419) );
  MUX21X1_LVT csr_U688 ( .A1(csr_n1411), .A2(csr_n1410), .S0(
        ibuf_io_inst_0_bits_raw[20]), .Y(csr_n1415) );
  MUX21X1_LVT csr_U687 ( .A1(csr_n905), .A2(csr_n904), .S0(csr_n1201), .Y(
        csr_n906) );
  NAND2X0_LVT csr_U686 ( .A1(csr_n906), .A2(csr_n381), .Y(csr_n1255) );
  MUX21X1_LVT csr_U685 ( .A1(csr_n927), .A2(csr_n926), .S0(csr_n387), .Y(
        csr_n928) );
  NAND4X0_LVT csr_U684 ( .A1(csr_n915), .A2(csr_n590), .A3(csr_n387), .A4(
        csr_n501), .Y(csr_n921) );
  NBUFFX2_LVT csr_U683 ( .A(n3785), .Y(csr_n592) );
  NBUFFX2_LVT csr_U682 ( .A(csr_n531), .Y(csr_n543) );
  NBUFFX2_LVT csr_U681 ( .A(csr_n531), .Y(csr_n541) );
  NBUFFX2_LVT csr_U680 ( .A(csr_n531), .Y(csr_n542) );
  NBUFFX2_LVT csr_U679 ( .A(csr_n531), .Y(csr_n544) );
  NAND3X0_LVT csr_U678 ( .A1(csr_n1462), .A2(csr_n1443), .A3(csr_n501), .Y(
        csr_n1917) );
  NAND4X0_LVT csr_U677 ( .A1(csr_n940), .A2(csr_n590), .A3(csr_n939), .A4(
        csr_n938), .Y(csr_n2160) );
  NBUFFX2_LVT csr_U676 ( .A(csr_net35092), .Y(csr_n532) );
  NBUFFX2_LVT csr_U675 ( .A(csr_net35092), .Y(csr_n533) );
  NBUFFX2_LVT csr_U674 ( .A(csr_net35092), .Y(csr_n534) );
  NBUFFX2_LVT csr_U673 ( .A(csr_net35092), .Y(csr_n535) );
  NBUFFX2_LVT csr_U672 ( .A(csr_net35092), .Y(csr_n536) );
  NBUFFX2_LVT csr_U671 ( .A(csr_net35092), .Y(csr_n537) );
  NBUFFX2_LVT csr_U670 ( .A(csr_net35092), .Y(csr_n539) );
  NBUFFX2_LVT csr_U669 ( .A(csr_net35092), .Y(csr_n540) );
  NBUFFX2_LVT csr_U668 ( .A(csr_net35092), .Y(csr_n538) );
  NBUFFX2_LVT csr_U667 ( .A(csr_n1128), .Y(csr_n491) );
  NBUFFX2_LVT csr_U666 ( .A(csr_net34895), .Y(csr_n572) );
  NBUFFX2_LVT csr_U665 ( .A(csr_net34930), .Y(csr_n559) );
  NBUFFX2_LVT csr_U664 ( .A(csr_net34895), .Y(csr_n574) );
  NBUFFX2_LVT csr_U663 ( .A(csr_net34895), .Y(csr_n573) );
  NBUFFX2_LVT csr_U662 ( .A(n3785), .Y(csr_n593) );
  NBUFFX2_LVT csr_U661 ( .A(csr_net34930), .Y(csr_n561) );
  NBUFFX2_LVT csr_U660 ( .A(csr_net34930), .Y(csr_n560) );
  NBUFFX2_LVT csr_U659 ( .A(csr_net34925), .Y(csr_n564) );
  NBUFFX2_LVT csr_U658 ( .A(csr_net34925), .Y(csr_n562) );
  NBUFFX2_LVT csr_U657 ( .A(csr_net34955), .Y(csr_n550) );
  NBUFFX2_LVT csr_U656 ( .A(csr_net34955), .Y(csr_n552) );
  NBUFFX2_LVT csr_U655 ( .A(csr_net34955), .Y(csr_n548) );
  NBUFFX2_LVT csr_U654 ( .A(csr_net34925), .Y(csr_n566) );
  NBUFFX2_LVT csr_U653 ( .A(csr_net35309), .Y(csr_n526) );
  NBUFFX2_LVT csr_U652 ( .A(csr_net35309), .Y(csr_n524) );
  NBUFFX2_LVT csr_U651 ( .A(csr_net35309), .Y(csr_n523) );
  NBUFFX2_LVT csr_U650 ( .A(csr_net35309), .Y(csr_n522) );
  NBUFFX2_LVT csr_U649 ( .A(csr_net34955), .Y(csr_n549) );
  NBUFFX2_LVT csr_U648 ( .A(csr_net34925), .Y(csr_n563) );
  NBUFFX2_LVT csr_U647 ( .A(csr_net35309), .Y(csr_n525) );
  NBUFFX2_LVT csr_U646 ( .A(csr_net34925), .Y(csr_n565) );
  NBUFFX2_LVT csr_U645 ( .A(csr_net34955), .Y(csr_n551) );
  NBUFFX2_LVT csr_U644 ( .A(csr_net34880), .Y(csr_n583) );
  NBUFFX2_LVT csr_U643 ( .A(csr_net35304), .Y(csr_n528) );
  NBUFFX2_LVT csr_U642 ( .A(csr_net35082), .Y(csr_n547) );
  NBUFFX2_LVT csr_U641 ( .A(csr_net34880), .Y(csr_n582) );
  NBUFFX2_LVT csr_U640 ( .A(csr_net35082), .Y(csr_n545) );
  NBUFFX2_LVT csr_U639 ( .A(csr_net35082), .Y(csr_n546) );
  NBUFFX2_LVT csr_U638 ( .A(csr_net35304), .Y(csr_n530) );
  NBUFFX2_LVT csr_U637 ( .A(csr_net34880), .Y(csr_n581) );
  NBUFFX2_LVT csr_U636 ( .A(csr_net35304), .Y(csr_n529) );
  NBUFFX2_LVT csr_U635 ( .A(csr_net34890), .Y(csr_n578) );
  NBUFFX2_LVT csr_U634 ( .A(csr_net34890), .Y(csr_n575) );
  NBUFFX2_LVT csr_U633 ( .A(csr_net34890), .Y(csr_n577) );
  NBUFFX2_LVT csr_U632 ( .A(csr_net34890), .Y(csr_n576) );
  NBUFFX2_LVT csr_U631 ( .A(csr_net34920), .Y(csr_n568) );
  NBUFFX2_LVT csr_U630 ( .A(csr_net34920), .Y(csr_n570) );
  NBUFFX2_LVT csr_U629 ( .A(csr_net34920), .Y(csr_n569) );
  NBUFFX2_LVT csr_U628 ( .A(csr_net34890), .Y(csr_n579) );
  NBUFFX2_LVT csr_U627 ( .A(csr_net34950), .Y(csr_n555) );
  NBUFFX2_LVT csr_U626 ( .A(csr_net34950), .Y(csr_n554) );
  NBUFFX2_LVT csr_U625 ( .A(csr_net35309), .Y(csr_n527) );
  NBUFFX2_LVT csr_U624 ( .A(csr_net34955), .Y(csr_n553) );
  NBUFFX2_LVT csr_U623 ( .A(csr_net34925), .Y(csr_n567) );
  NBUFFX2_LVT csr_U622 ( .A(csr_net34950), .Y(csr_n556) );
  NBUFFX2_LVT csr_U621 ( .A(csr_net34722), .Y(csr_n584) );
  NBUFFX2_LVT csr_U620 ( .A(csr_net34722), .Y(csr_n585) );
  NBUFFX2_LVT csr_U619 ( .A(csr_net34722), .Y(csr_n586) );
  NBUFFX2_LVT csr_U618 ( .A(n3785), .Y(csr_n594) );
  OAI21X1_LVT csr_U617 ( .A1(csr_n_T_45_2_), .A2(csr_n956), .A3(csr_n961), .Y(
        csr_n958) );
  MUX21X1_LVT csr_U616 ( .A1(csr_io_pc[9]), .A2(csr_wdata_9_), .S0(csr_n514), 
        .Y(csr_net35055) );
  MUX21X1_LVT csr_U615 ( .A1(csr_io_pc[3]), .A2(csr_wdata_3_), .S0(csr_n515), 
        .Y(csr_net35295) );
  MUX21X1_LVT csr_U614 ( .A1(csr_n588), .A2(csr_n880), .S0(csr_n879), .Y(
        csr_n1909) );
  IBUFFX4_LVT csr_U613 ( .A(reset), .Y(csr_n590) );
  NBUFFX2_LVT csr_U612 ( .A(csr_net35092), .Y(csr_n531) );
  OR2X1_LVT csr_U611 ( .A1(csr_io_rw_addr[6]), .A2(csr_io_rw_addr[9]), .Y(
        csr_n605) );
  NOR2X1_LVT csr_U610 ( .A1(io_ptw_status_prv[0]), .A2(csr_io_rw_addr[0]), .Y(
        csr_n953) );
  INVX0_LVT csr_U609 ( .A(csr_n597), .Y(csr_n598) );
  INVX0_LVT csr_U608 ( .A(ibuf_io_inst_0_bits_raw[28]), .Y(csr_n1371) );
  INVX0_LVT csr_U607 ( .A(csr_n605), .Y(csr_n633) );
  INVX1_LVT csr_U606 ( .A(ibuf_io_inst_0_bits_raw[30]), .Y(csr_n489) );
  OR2X1_LVT csr_U605 ( .A1(ibuf_io_inst_0_bits_raw[24]), .A2(
        ibuf_io_inst_0_bits_raw[23]), .Y(csr_n1392) );
  AND2X1_LVT csr_U604 ( .A1(csr_n630), .A2(csr_n1518), .Y(csr_n1512) );
  NOR4X0_LVT csr_U603 ( .A1(csr_io_rw_addr[4]), .A2(csr_io_rw_addr[3]), .A3(
        csr_n1525), .A4(csr_n1524), .Y(csr_n1526) );
  INVX0_LVT csr_U602 ( .A(csr_n1172), .Y(csr_n1173) );
  INVX0_LVT csr_U601 ( .A(csr_n1176), .Y(csr_n1187) );
  NOR2X1_LVT csr_U600 ( .A1(ibuf_io_inst_0_bits_inst_rs3_2_), .A2(
        ibuf_io_inst_0_bits_raw[26]), .Y(csr_n1379) );
  INVX1_LVT csr_U599 ( .A(csr_n489), .Y(csr_n490) );
  NOR2X1_LVT csr_U598 ( .A1(ibuf_io_inst_0_bits_raw[21]), .A2(
        ibuf_io_inst_0_bits_raw[20]), .Y(csr_n1390) );
  INVX0_LVT csr_U597 ( .A(csr_n1178), .Y(csr_n1177) );
  OR2X1_LVT csr_U596 ( .A1(io_interrupts_seip), .A2(csr_n_T_3694_9_), .Y(
        csr_n1136) );
  INVX0_LVT csr_U595 ( .A(csr_n1134), .Y(csr_n941) );
  NAND2X0_LVT csr_U594 ( .A1(csr_n504), .A2(csr_n590), .Y(csr_n389) );
  NOR2X1_LVT csr_U593 ( .A1(csr_n427), .A2(wb_cause[3]), .Y(csr_n901) );
  AND2X1_LVT csr_U592 ( .A1(csr_n858), .A2(csr_n857), .Y(csr_n1469) );
  INVX0_LVT csr_U591 ( .A(csr_n1192), .Y(csr_n1184) );
  NOR2X1_LVT csr_U590 ( .A1(csr_n605), .A2(csr_n601), .Y(csr_n488) );
  AND2X1_LVT csr_U589 ( .A1(csr_n620), .A2(csr_n676), .Y(csr_n1153) );
  INVX0_LVT csr_U588 ( .A(csr_n1144), .Y(csr_n1141) );
  AND2X1_LVT csr_U587 ( .A1(csr_n620), .A2(csr_n1505), .Y(csr_n1474) );
  INVX0_LVT csr_U586 ( .A(csr_n1179), .Y(csr_n1169) );
  INVX0_LVT csr_U585 ( .A(csr_n866), .Y(csr_n743) );
  NOR2X1_LVT csr_U584 ( .A1(csr_n1520), .A2(csr_n1697), .Y(csr_n1210) );
  INVX0_LVT csr_U583 ( .A(csr_n1368), .Y(csr_n1369) );
  INVX0_LVT csr_U582 ( .A(csr_n1697), .Y(csr_n699) );
  MUX21X1_LVT csr_U581 ( .A1(csr_n953), .A2(csr_n954), .S0(csr_n1697), .Y(
        csr_n891) );
  NOR2X1_LVT csr_U580 ( .A1(csr_io_rw_addr[9]), .A2(csr_n1903), .Y(csr_n1355)
         );
  MUX21X1_LVT csr_U579 ( .A1(csr_n1520), .A2(wb_cause[3]), .S0(csr_n1697), .Y(
        csr_n1226) );
  MUX21X1_LVT csr_U578 ( .A1(csr_n700), .A2(wb_cause[1]), .S0(csr_n1697), .Y(
        csr_n1209) );
  INVX0_LVT csr_U577 ( .A(csr_n1903), .Y(csr_n1199) );
  INVX0_LVT csr_U576 ( .A(csr_n1154), .Y(csr_n1026) );
  INVX0_LVT csr_U575 ( .A(csr_n1210), .Y(csr_n1211) );
  AND3X1_LVT csr_U574 ( .A1(csr_io_rw_addr[1]), .A2(csr_n1520), .A3(csr_n1531), 
        .Y(csr_n1689) );
  INVX0_LVT csr_U573 ( .A(csr_n1155), .Y(csr_n1156) );
  INVX0_LVT csr_U572 ( .A(csr_n1384), .Y(csr_n1385) );
  INVX0_LVT csr_U571 ( .A(csr_n1378), .Y(csr_n1380) );
  OR2X1_LVT csr_U570 ( .A1(csr_n699), .A2(csr_io_exception), .Y(csr_n1139) );
  INVX1_LVT csr_U569 ( .A(csr_n1041), .Y(csr_n1157) );
  INVX1_LVT csr_U568 ( .A(csr_n891), .Y(csr_n1202) );
  INVX0_LVT csr_U567 ( .A(csr_n1226), .Y(csr_n895) );
  INVX0_LVT csr_U566 ( .A(csr_n1209), .Y(csr_n888) );
  NAND3X0_LVT csr_U565 ( .A1(csr_n503), .A2(csr_n672), .A3(csr_n671), .Y(
        csr_n957) );
  INVX0_LVT csr_U564 ( .A(csr_n1171), .Y(csr_n1170) );
  INVX0_LVT csr_U563 ( .A(csr_n1139), .Y(csr_n1442) );
  INVX0_LVT csr_U562 ( .A(csr_n1455), .Y(csr_n923) );
  NOR2X1_LVT csr_U561 ( .A1(csr_n1180), .A2(csr_n1189), .Y(csr_n1185) );
  INVX0_LVT csr_U560 ( .A(csr_n1445), .Y(csr_n1447) );
  INVX0_LVT csr_U559 ( .A(csr_n702), .Y(csr_n949) );
  NOR2X1_LVT csr_U558 ( .A1(csr_n1584), .A2(csr_n1583), .Y(csr_n1109) );
  AND2X1_LVT csr_U557 ( .A1(csr_n629), .A2(csr_n590), .Y(csr_n1446) );
  INVX0_LVT csr_U556 ( .A(csr_n1375), .Y(csr_n1377) );
  INVX0_LVT csr_U555 ( .A(csr_n1419), .Y(csr_n1420) );
  OA22X1_LVT csr_U554 ( .A1(csr_n490), .A2(csr_n1419), .A3(
        ibuf_io_inst_0_bits_raw[27]), .A4(csr_n1398), .Y(csr_n1404) );
  INVX0_LVT csr_U553 ( .A(csr_n1381), .Y(csr_n1367) );
  INVX0_LVT csr_U552 ( .A(csr_n1495), .Y(csr_n484) );
  INVX0_LVT csr_U551 ( .A(csr_n961), .Y(csr_n1458) );
  OR2X1_LVT csr_U550 ( .A1(csr_n708), .A2(csr_n1467), .Y(csr_n1257) );
  NOR2X1_LVT csr_U549 ( .A1(csr_n1621), .A2(csr_n1624), .Y(csr_n1052) );
  INVX0_LVT csr_U548 ( .A(csr_n1432), .Y(csr_n1433) );
  NOR2X1_LVT csr_U547 ( .A1(csr_n1585), .A2(csr_n1586), .Y(csr_n1107) );
  NOR2X1_LVT csr_U546 ( .A1(csr_n1590), .A2(csr_n1589), .Y(csr_n1094) );
  NOR2X1_LVT csr_U545 ( .A1(csr_n1140), .A2(csr_n1139), .Y(csr_N1821) );
  NOR2X1_LVT csr_U544 ( .A1(csr_n1653), .A2(csr_n1657), .Y(csr_n650) );
  INVX0_LVT csr_U543 ( .A(csr_n1427), .Y(csr_n1418) );
  NOR2X1_LVT csr_U542 ( .A1(csr_n1458), .A2(csr_n956), .Y(csr_n712) );
  NOR2X1_LVT csr_U541 ( .A1(csr_n1481), .A2(csr_n1690), .Y(csr_n968) );
  INVX0_LVT csr_U540 ( .A(csr_n1374), .Y(csr_n1373) );
  INVX0_LVT csr_U539 ( .A(csr_n1416), .Y(csr_n1436) );
  INVX0_LVT csr_U538 ( .A(csr_n908), .Y(csr_n911) );
  OR2X1_LVT csr_U537 ( .A1(csr_n1199), .A2(csr_n1441), .Y(csr_n1352) );
  INVX1_LVT csr_U536 ( .A(csr_n925), .Y(csr_n1461) );
  OR2X1_LVT csr_U535 ( .A1(csr_n1442), .A2(csr_n1441), .Y(csr_n1462) );
  INVX1_LVT csr_U534 ( .A(csr_n1352), .Y(csr_n1348) );
  INVX0_LVT csr_U533 ( .A(csr_n1468), .Y(csr_n1346) );
  IBUFFX2_LVT csr_U532 ( .A(csr_n590), .Y(csr_n376) );
  INVX1_LVT csr_U531 ( .A(io_interrupts_debug), .Y(csr_n1186) );
  INVX1_LVT csr_U530 ( .A(csr_n590), .Y(csr_n378) );
  INVX1_LVT csr_U529 ( .A(csr_io_rw_addr[4]), .Y(csr_n1521) );
  NOR2X1_LVT csr_U528 ( .A1(csr_io_rw_addr[0]), .A2(csr_io_rw_addr[1]), .Y(
        csr_n630) );
  INVX0_LVT csr_U527 ( .A(csr_io_rw_addr[9]), .Y(csr_n1515) );
  INVX1_LVT csr_U526 ( .A(io_imem_sfence_bits_addr[1]), .Y(csr_n697) );
  INVX1_LVT csr_U525 ( .A(csr_io_rw_addr[1]), .Y(csr_n1519) );
  NOR2X1_LVT csr_U524 ( .A1(csr_io_rw_addr[4]), .A2(csr_io_rw_addr[3]), .Y(
        csr_n1529) );
  INVX0_LVT csr_U523 ( .A(csr_io_rw_addr[7]), .Y(csr_n1528) );
  INVX0_LVT csr_U522 ( .A(csr_io_rw_addr[2]), .Y(csr_n1518) );
  INVX1_LVT csr_U521 ( .A(io_imem_sfence_bits_addr[5]), .Y(csr_n1904) );
  INVX1_LVT csr_U520 ( .A(io_imem_sfence_bits_addr[9]), .Y(csr_n1907) );
  INVX1_LVT csr_U519 ( .A(ibuf_io_inst_0_bits_raw[23]), .Y(csr_n1430) );
  INVX1_LVT csr_U518 ( .A(ibuf_io_inst_0_bits_raw[22]), .Y(csr_n1417) );
  INVX1_LVT csr_U517 ( .A(n2576), .Y(csr_n1405) );
  INVX1_LVT csr_U516 ( .A(ibuf_io_inst_0_bits_raw[26]), .Y(csr_n1376) );
  INVX0_LVT csr_U515 ( .A(ibuf_io_inst_0_bits_raw[25]), .Y(csr_n1406) );
  INVX1_LVT csr_U514 ( .A(wb_cause[1]), .Y(csr_n902) );
  INVX1_LVT csr_U513 ( .A(wb_cause[0]), .Y(csr_n954) );
  INVX2_LVT csr_U512 ( .A(csr_n389), .Y(csr_n375) );
  INVX1_LVT csr_U511 ( .A(csr_n389), .Y(csr_n503) );
  IBUFFX2_LVT csr_U510 ( .A(csr_n957), .Y(csr_n1128) );
  AND2X1_LVT csr_U509 ( .A1(csr_n1446), .A2(csr_n1445), .Y(csr_n1150) );
  AND2X1_LVT csr_U508 ( .A1(csr_n1459), .A2(csr_n673), .Y(csr_n1129) );
  AND2X1_LVT csr_U507 ( .A1(csr_n375), .A2(csr_wdata_55_), .Y(csr_n374) );
  OR2X1_LVT csr_U506 ( .A1(csr_n860), .A2(csr_n372), .Y(csr_n373) );
  AND2X1_LVT csr_U505 ( .A1(csr_n590), .A2(csr_wdata_0_), .Y(csr_n371) );
  AND2X1_LVT csr_U504 ( .A1(csr_wdata_48_), .A2(csr_wdata_49_), .Y(csr_n369)
         );
  AND2X4_LVT csr_U503 ( .A1(csr_n1139), .A2(csr_n1457), .Y(csr_n1152) );
  IBUFFX8_LVT csr_U502 ( .A(csr_n629), .Y(csr_n1149) );
  AND2X4_LVT csr_U501 ( .A1(csr_n1139), .A2(csr_n1456), .Y(csr_n1159) );
  IBUFFX2_LVT csr_U500 ( .A(csr_wdata_3_), .Y(csr_n588) );
  AO22X1_LVT csr_U498 ( .A1(csr_n1149), .A2(csr_wdata_0_), .A3(csr_n361), .A4(
        csr_n1446), .Y(csr_N1822) );
  HADDX1_LVT csr_U497 ( .A0(csr_io_csr_stall), .B0(csr_n417), .SO(csr_n361) );
  OA222X1_LVT csr_U496 ( .A1(io_imem_sfence_bits_addr[12]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[12]), .A4(csr_io_rw_rdata[12]), .A5(
        csr_n516), .A6(csr_n360), .Y(csr_wdata_12_) );
  INVX0_LVT csr_U495 ( .A(io_imem_sfence_bits_addr[12]), .Y(csr_n360) );
  OA222X1_LVT csr_U494 ( .A1(io_imem_sfence_bits_addr[8]), .A2(csr_n589), .A3(
        io_imem_sfence_bits_addr[8]), .A4(csr_io_rw_rdata[8]), .A5(csr_n516), 
        .A6(csr_n359), .Y(csr_wdata_8_) );
  INVX0_LVT csr_U493 ( .A(io_imem_sfence_bits_addr[8]), .Y(csr_n359) );
  OAI22X1_LVT csr_U492 ( .A1(csr_n1455), .A2(csr_n1483), .A3(csr_n899), .A4(
        csr_n358), .Y(csr_N1272) );
  INVX0_LVT csr_U491 ( .A(csr_n1501), .Y(csr_n358) );
  OA222X1_LVT csr_U490 ( .A1(io_imem_sfence_bits_addr[38]), .A2(
        csr_io_rw_rdata[38]), .A3(io_imem_sfence_bits_addr[38]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n357), .Y(csr_wdata_38_) );
  INVX0_LVT csr_U489 ( .A(io_imem_sfence_bits_addr[38]), .Y(csr_n357) );
  OA222X1_LVT csr_U488 ( .A1(n_T_1165[54]), .A2(csr_io_rw_rdata[54]), .A3(
        n_T_1165[54]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n356), .Y(
        csr_wdata_54_) );
  INVX0_LVT csr_U487 ( .A(n_T_1165[54]), .Y(csr_n356) );
  OA222X1_LVT csr_U486 ( .A1(n_T_1165[47]), .A2(csr_io_rw_rdata[47]), .A3(
        n_T_1165[47]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n355), .Y(
        csr_wdata_47_) );
  INVX0_LVT csr_U485 ( .A(n_T_1165[47]), .Y(csr_n355) );
  OA222X1_LVT csr_U484 ( .A1(n_T_1165[46]), .A2(csr_io_rw_rdata[46]), .A3(
        n_T_1165[46]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n354), .Y(
        csr_wdata_46_) );
  INVX0_LVT csr_U483 ( .A(n_T_1165[46]), .Y(csr_n354) );
  OA222X1_LVT csr_U482 ( .A1(n_T_1165[61]), .A2(csr_io_rw_rdata[61]), .A3(
        n_T_1165[61]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n353), .Y(
        csr_wdata_61_) );
  INVX0_LVT csr_U481 ( .A(n_T_1165[61]), .Y(csr_n353) );
  OA222X1_LVT csr_U480 ( .A1(io_imem_sfence_bits_addr[35]), .A2(
        csr_io_rw_rdata[35]), .A3(io_imem_sfence_bits_addr[35]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n352), .Y(csr_wdata_35_) );
  INVX0_LVT csr_U479 ( .A(io_imem_sfence_bits_addr[35]), .Y(csr_n352) );
  OA222X1_LVT csr_U478 ( .A1(io_imem_sfence_bits_addr[34]), .A2(
        csr_io_rw_rdata[34]), .A3(io_imem_sfence_bits_addr[34]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n351), .Y(csr_wdata_34_) );
  INVX0_LVT csr_U477 ( .A(io_imem_sfence_bits_addr[34]), .Y(csr_n351) );
  OA222X1_LVT csr_U476 ( .A1(io_imem_sfence_bits_addr[32]), .A2(
        csr_io_rw_rdata[32]), .A3(io_imem_sfence_bits_addr[32]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n350), .Y(csr_wdata_32_) );
  INVX0_LVT csr_U475 ( .A(io_imem_sfence_bits_addr[32]), .Y(csr_n350) );
  OA222X1_LVT csr_U474 ( .A1(io_imem_sfence_bits_addr[31]), .A2(
        csr_io_rw_rdata[31]), .A3(io_imem_sfence_bits_addr[31]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n349), .Y(csr_wdata_31_) );
  INVX0_LVT csr_U473 ( .A(io_imem_sfence_bits_addr[31]), .Y(csr_n349) );
  OA222X1_LVT csr_U472 ( .A1(io_imem_sfence_bits_addr[13]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[13]), .A4(csr_io_rw_rdata[13]), .A5(
        csr_n516), .A6(csr_n348), .Y(csr_wdata_13_) );
  INVX0_LVT csr_U471 ( .A(io_imem_sfence_bits_addr[13]), .Y(csr_n348) );
  OA222X1_LVT csr_U470 ( .A1(io_imem_sfence_bits_addr[23]), .A2(
        csr_io_rw_rdata[23]), .A3(io_imem_sfence_bits_addr[23]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n347), .Y(csr_wdata_23_) );
  INVX0_LVT csr_U469 ( .A(io_imem_sfence_bits_addr[23]), .Y(csr_n347) );
  OA222X1_LVT csr_U468 ( .A1(io_imem_sfence_bits_addr[19]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[19]), .A4(csr_io_rw_rdata[19]), .A5(
        csr_n516), .A6(csr_n346), .Y(csr_wdata_19_) );
  INVX0_LVT csr_U467 ( .A(io_imem_sfence_bits_addr[19]), .Y(csr_n346) );
  OA222X1_LVT csr_U466 ( .A1(io_imem_sfence_bits_addr[15]), .A2(
        csr_io_rw_rdata[15]), .A3(io_imem_sfence_bits_addr[15]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n345), .Y(csr_wdata_15_) );
  INVX0_LVT csr_U465 ( .A(io_imem_sfence_bits_addr[15]), .Y(csr_n345) );
  OA222X1_LVT csr_U464 ( .A1(io_imem_sfence_bits_addr[16]), .A2(
        csr_io_rw_rdata[16]), .A3(io_imem_sfence_bits_addr[16]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n344), .Y(csr_wdata_16_) );
  INVX0_LVT csr_U463 ( .A(io_imem_sfence_bits_addr[16]), .Y(csr_n344) );
  OA222X1_LVT csr_U462 ( .A1(io_imem_sfence_bits_addr[27]), .A2(
        csr_io_rw_rdata[27]), .A3(io_imem_sfence_bits_addr[27]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n343), .Y(csr_wdata_27_) );
  INVX0_LVT csr_U461 ( .A(io_imem_sfence_bits_addr[27]), .Y(csr_n343) );
  OA222X1_LVT csr_U460 ( .A1(io_imem_sfence_bits_addr[29]), .A2(
        csr_io_rw_rdata[29]), .A3(io_imem_sfence_bits_addr[29]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n342), .Y(csr_wdata_29_) );
  INVX0_LVT csr_U459 ( .A(io_imem_sfence_bits_addr[29]), .Y(csr_n342) );
  OA222X1_LVT csr_U458 ( .A1(io_imem_sfence_bits_addr[14]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[14]), .A4(csr_io_rw_rdata[14]), .A5(
        csr_n516), .A6(csr_n341), .Y(csr_wdata_14_) );
  INVX0_LVT csr_U457 ( .A(io_imem_sfence_bits_addr[14]), .Y(csr_n341) );
  OA222X1_LVT csr_U456 ( .A1(io_imem_sfence_bits_addr[4]), .A2(csr_n589), .A3(
        io_imem_sfence_bits_addr[4]), .A4(csr_io_rw_rdata[4]), .A5(csr_n516), 
        .A6(csr_n340), .Y(csr_wdata_4_) );
  INVX0_LVT csr_U455 ( .A(io_imem_sfence_bits_addr[4]), .Y(csr_n340) );
  OA222X1_LVT csr_U454 ( .A1(io_imem_sfence_bits_addr[6]), .A2(
        csr_io_rw_rdata[6]), .A3(io_imem_sfence_bits_addr[6]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n339), .Y(csr_wdata_6_) );
  INVX0_LVT csr_U453 ( .A(io_imem_sfence_bits_addr[6]), .Y(csr_n339) );
  AND2X1_LVT csr_U452 ( .A1(csr_n1527), .A2(csr_n338), .Y(csr_n1487) );
  AND4X1_LVT csr_U451 ( .A1(csr_io_rw_addr[0]), .A2(csr_io_rw_addr[2]), .A3(
        csr_n1519), .A4(csr_n633), .Y(csr_n338) );
  NAND3X0_LVT csr_U450 ( .A1(csr_n328), .A2(csr_n329), .A3(csr_n337), .Y(
        csr_io_rw_rdata[21]) );
  NOR4X0_LVT csr_U449 ( .A1(csr_n330), .A2(csr_n331), .A3(csr_n332), .A4(
        csr_n336), .Y(csr_n337) );
  AO22X1_LVT csr_U447 ( .A1(csr_n1508), .A2(csr_reg_sscratch[21]), .A3(
        csr_n1157), .A4(csr_n1925), .Y(csr_n334) );
  AO222X1_LVT csr_U446 ( .A1(csr_n1689), .A2(csr_n_T_45_21_), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_21_), .A5(csr_n1487), .A6(csr_reg_stvec_21_), .Y(
        csr_n333) );
  AO22X1_LVT csr_U445 ( .A1(csr_n1160), .A2(csr_n_T_444[21]), .A3(csr_n1489), 
        .A4(csr_reg_mepc_21_), .Y(csr_n332) );
  AO22X1_LVT csr_U444 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[21]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[21]), .Y(csr_n331) );
  AO22X1_LVT csr_U443 ( .A1(csr_n1485), .A2(csr_reg_mscratch[21]), .A3(
        csr_n1493), .A4(csr_reg_dpc_21_), .Y(csr_n330) );
  AOI22X1_LVT csr_U442 ( .A1(csr_n1506), .A2(csr_reg_sepc_21_), .A3(csr_n1490), 
        .A4(csr_io_bp_0_address[21]), .Y(csr_n329) );
  NOR4X0_LVT csr_U441 ( .A1(csr_n324), .A2(csr_n325), .A3(csr_n326), .A4(
        csr_n327), .Y(csr_n328) );
  AO22X1_LVT csr_U440 ( .A1(csr_n1510), .A2(csr_reg_dscratch[21]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[21]), .Y(csr_n327) );
  AO22X1_LVT csr_U439 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[21]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[21]), .Y(csr_n326) );
  AO22X1_LVT csr_U438 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[21]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[21]), .Y(csr_n325) );
  AO22X1_LVT csr_U437 ( .A1(csr_n1162), .A2(csr_io_time[21]), .A3(csr_n1472), 
        .A4(io_ptw_pmp_5_addr[21]), .Y(csr_n324) );
  OR3X1_LVT csr_U436 ( .A1(csr_n1392), .A2(csr_n490), .A3(
        ibuf_io_inst_0_bits_raw[25]), .Y(csr_n1378) );
  AO21X1_LVT csr_U435 ( .A1(csr_n1190), .A2(csr_n322), .A3(csr_n1182), .Y(
        csr_n323) );
  INVX0_LVT csr_U434 ( .A(csr_n1181), .Y(csr_n322) );
  OA222X1_LVT csr_U433 ( .A1(io_imem_sfence_bits_addr[0]), .A2(csr_n589), .A3(
        io_imem_sfence_bits_addr[0]), .A4(csr_io_rw_rdata[0]), .A5(csr_n516), 
        .A6(csr_n321), .Y(csr_wdata_0_) );
  INVX0_LVT csr_U432 ( .A(io_imem_sfence_bits_addr[0]), .Y(csr_n321) );
  OA222X1_LVT csr_U431 ( .A1(io_imem_sfence_bits_addr[7]), .A2(csr_n589), .A3(
        io_imem_sfence_bits_addr[7]), .A4(csr_io_rw_rdata[7]), .A5(csr_n516), 
        .A6(csr_n320), .Y(csr_wdata_7_) );
  INVX0_LVT csr_U430 ( .A(io_imem_sfence_bits_addr[7]), .Y(csr_n320) );
  AND3X1_LVT csr_U429 ( .A1(csr_n503), .A2(csr_n319), .A3(csr_io_status_debug), 
        .Y(csr_n1482) );
  OA222X1_LVT csr_U428 ( .A1(n_T_1165[59]), .A2(csr_n_T_366_59_), .A3(
        n_T_1165[59]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n318), .Y(
        csr_n319) );
  INVX0_LVT csr_U427 ( .A(n_T_1165[59]), .Y(csr_n318) );
  AO22X1_LVT csr_U426 ( .A1(csr_n497), .A2(csr_n_T_52[48]), .A3(csr_wdata_54_), 
        .A4(csr_n1149), .Y(csr_N1939) );
  OA222X1_LVT csr_U425 ( .A1(n_T_1165[43]), .A2(csr_io_rw_rdata[43]), .A3(
        n_T_1165[43]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n317), .Y(
        csr_wdata_43_) );
  INVX0_LVT csr_U424 ( .A(n_T_1165[43]), .Y(csr_n317) );
  OA222X1_LVT csr_U423 ( .A1(io_imem_sfence_bits_addr[37]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[37]), .A4(csr_io_rw_rdata[37]), .A5(
        csr_n516), .A6(csr_n316), .Y(csr_wdata_37_) );
  INVX0_LVT csr_U422 ( .A(io_imem_sfence_bits_addr[37]), .Y(csr_n316) );
  OA222X1_LVT csr_U421 ( .A1(io_imem_sfence_bits_addr[36]), .A2(
        csr_io_rw_rdata[36]), .A3(io_imem_sfence_bits_addr[36]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n315), .Y(csr_wdata_36_) );
  INVX0_LVT csr_U420 ( .A(io_imem_sfence_bits_addr[36]), .Y(csr_n315) );
  OA222X1_LVT csr_U419 ( .A1(io_imem_sfence_bits_addr[33]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[33]), .A4(csr_io_rw_rdata[33]), .A5(
        csr_n516), .A6(csr_n314), .Y(csr_wdata_33_) );
  INVX0_LVT csr_U418 ( .A(io_imem_sfence_bits_addr[33]), .Y(csr_n314) );
  OA222X1_LVT csr_U417 ( .A1(io_imem_sfence_bits_addr[30]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[30]), .A4(csr_io_rw_rdata[30]), .A5(
        csr_n516), .A6(csr_n313), .Y(csr_wdata_30_) );
  INVX0_LVT csr_U416 ( .A(io_imem_sfence_bits_addr[30]), .Y(csr_n313) );
  OA222X1_LVT csr_U415 ( .A1(io_imem_sfence_bits_addr[28]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[28]), .A4(csr_io_rw_rdata[28]), .A5(
        csr_n516), .A6(csr_n312), .Y(csr_wdata_28_) );
  INVX0_LVT csr_U414 ( .A(io_imem_sfence_bits_addr[28]), .Y(csr_n312) );
  OA222X1_LVT csr_U413 ( .A1(io_imem_sfence_bits_addr[18]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[18]), .A4(csr_io_rw_rdata[18]), .A5(
        csr_n516), .A6(csr_n311), .Y(csr_wdata_18_) );
  INVX0_LVT csr_U412 ( .A(io_imem_sfence_bits_addr[18]), .Y(csr_n311) );
  OA222X1_LVT csr_U411 ( .A1(io_imem_sfence_bits_addr[20]), .A2(
        csr_io_rw_rdata[20]), .A3(io_imem_sfence_bits_addr[20]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n310), .Y(csr_wdata_20_) );
  INVX0_LVT csr_U410 ( .A(io_imem_sfence_bits_addr[20]), .Y(csr_n310) );
  OA222X1_LVT csr_U409 ( .A1(io_imem_sfence_bits_addr[21]), .A2(
        csr_io_rw_rdata[21]), .A3(io_imem_sfence_bits_addr[21]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n309), .Y(csr_wdata_21_) );
  INVX0_LVT csr_U408 ( .A(io_imem_sfence_bits_addr[21]), .Y(csr_n309) );
  OA222X1_LVT csr_U407 ( .A1(io_imem_sfence_bits_addr[22]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[22]), .A4(csr_io_rw_rdata[22]), .A5(
        csr_n516), .A6(csr_n308), .Y(csr_wdata_22_) );
  INVX0_LVT csr_U406 ( .A(io_imem_sfence_bits_addr[22]), .Y(csr_n308) );
  OA222X1_LVT csr_U405 ( .A1(io_imem_sfence_bits_addr[24]), .A2(
        csr_io_rw_rdata[24]), .A3(io_imem_sfence_bits_addr[24]), .A4(csr_n589), 
        .A5(csr_n516), .A6(csr_n307), .Y(csr_wdata_24_) );
  INVX0_LVT csr_U404 ( .A(io_imem_sfence_bits_addr[24]), .Y(csr_n307) );
  OA222X1_LVT csr_U403 ( .A1(io_imem_sfence_bits_addr[26]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[26]), .A4(csr_io_rw_rdata[26]), .A5(
        csr_n516), .A6(csr_n306), .Y(csr_wdata_26_) );
  INVX0_LVT csr_U402 ( .A(io_imem_sfence_bits_addr[26]), .Y(csr_n306) );
  OA222X1_LVT csr_U401 ( .A1(io_imem_sfence_bits_addr[10]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[10]), .A4(csr_io_rw_rdata[10]), .A5(
        csr_n516), .A6(csr_n305), .Y(csr_wdata_10_) );
  INVX0_LVT csr_U400 ( .A(io_imem_sfence_bits_addr[10]), .Y(csr_n305) );
  NAND2X0_LVT csr_U399 ( .A1(csr_wdata_31_), .A2(csr_n304), .Y(csr_n370) );
  INVX0_LVT csr_U398 ( .A(csr_n376), .Y(csr_n304) );
  OA21X1_LVT csr_U397 ( .A1(csr_n1201), .A2(csr_n303), .A3(csr_n1471), .Y(
        csr_n366) );
  INVX0_LVT csr_U396 ( .A(csr_n1467), .Y(csr_n303) );
  AND3X1_LVT csr_U395 ( .A1(csr_n1514), .A2(csr_n1512), .A3(csr_n1526), .Y(
        csr_n1507) );
  AND3X1_LVT csr_U394 ( .A1(csr_io_time[0]), .A2(csr_io_time[1]), .A3(csr_n302), .Y(csr_n1142) );
  INVX0_LVT csr_U393 ( .A(csr_io_csr_stall), .Y(csr_n302) );
  NAND4X0_LVT csr_U392 ( .A1(csr_n284), .A2(csr_n292), .A3(csr_n296), .A4(
        csr_n301), .Y(csr_io_rw_rdata[8]) );
  NOR4X0_LVT csr_U391 ( .A1(csr_n297), .A2(csr_n298), .A3(csr_n299), .A4(
        csr_n300), .Y(csr_n301) );
  AO22X1_LVT csr_U390 ( .A1(csr_n1507), .A2(io_ptw_pmp_1_cfg_r), .A3(csr_n1506), .A4(csr_reg_sepc_8_), .Y(csr_n300) );
  AO22X1_LVT csr_U389 ( .A1(csr_n1508), .A2(csr_reg_sscratch[8]), .A3(
        csr_n1510), .A4(csr_reg_dscratch[8]), .Y(csr_n299) );
  AO22X1_LVT csr_U388 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[8]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[8]), .Y(csr_n298) );
  AO22X1_LVT csr_U387 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[8]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[8]), .Y(csr_n297) );
  NOR3X0_LVT csr_U386 ( .A1(csr_n293), .A2(csr_n294), .A3(csr_n295), .Y(
        csr_n296) );
  AO22X1_LVT csr_U385 ( .A1(csr_n1485), .A2(csr_reg_mscratch[8]), .A3(
        csr_n1489), .A4(csr_reg_mepc_8_), .Y(csr_n295) );
  AO22X1_LVT csr_U384 ( .A1(csr_n1162), .A2(csr_io_time[8]), .A3(csr_n1494), 
        .A4(io_ptw_pmp_6_addr[8]), .Y(csr_n294) );
  AO22X1_LVT csr_U383 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[8]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[8]), .Y(csr_n293) );
  NOR4X0_LVT csr_U382 ( .A1(csr_n288), .A2(csr_n289), .A3(csr_n290), .A4(
        csr_n291), .Y(csr_n292) );
  AO22X1_LVT csr_U381 ( .A1(csr_n1160), .A2(csr_n_T_444[8]), .A3(csr_n1469), 
        .A4(csr_read_medeleg_8), .Y(csr_n291) );
  AO22X1_LVT csr_U380 ( .A1(csr_n1153), .A2(csr_n_T_383[8]), .A3(csr_n1452), 
        .A4(csr_n1922), .Y(csr_n290) );
  AO22X1_LVT csr_U379 ( .A1(csr_n1487), .A2(csr_reg_stvec_8_), .A3(csr_n1154), 
        .A4(csr_n1931), .Y(csr_n289) );
  NAND3X0_LVT csr_U377 ( .A1(csr_n285), .A2(csr_n948), .A3(csr_n947), .Y(
        csr_n286) );
  NAND2X0_LVT csr_U376 ( .A1(io_ptw_ptbr_ppn[8]), .A2(csr_n1488), .Y(csr_n285)
         );
  AOI22X1_LVT csr_U375 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[8]), .A3(
        csr_n1481), .A4(csr_io_bp_0_control_tmatch[1]), .Y(csr_n284) );
  OR3X1_LVT csr_U374 ( .A1(csr_n280), .A2(csr_n281), .A3(csr_n283), .Y(
        csr_io_rw_rdata[38]) );
  AO22X1_LVT csr_U373 ( .A1(csr_n1160), .A2(csr_n_T_444[38]), .A3(csr_n1489), 
        .A4(csr_reg_mepc_38_), .Y(csr_n282) );
  AO22X1_LVT csr_U372 ( .A1(csr_n1510), .A2(csr_reg_dscratch[38]), .A3(
        csr_n1508), .A4(csr_reg_sscratch[38]), .Y(csr_n281) );
  AO22X1_LVT csr_U370 ( .A1(csr_n1506), .A2(csr_reg_sepc_38_), .A3(csr_n1153), 
        .A4(csr_n_T_383[38]), .Y(csr_n278) );
  AO22X1_LVT csr_U369 ( .A1(csr_n1689), .A2(csr_n_T_45_38_), .A3(csr_n1493), 
        .A4(csr_reg_dpc_38_), .Y(csr_n277) );
  OA222X1_LVT csr_U368 ( .A1(n_T_1165[53]), .A2(csr_io_rw_rdata[53]), .A3(
        n_T_1165[53]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n276), .Y(
        csr_wdata_53_) );
  INVX0_LVT csr_U367 ( .A(n_T_1165[53]), .Y(csr_n276) );
  OA222X1_LVT csr_U366 ( .A1(n_T_1165[42]), .A2(csr_io_rw_rdata[42]), .A3(
        n_T_1165[42]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n275), .Y(
        csr_wdata_42_) );
  INVX0_LVT csr_U365 ( .A(n_T_1165[42]), .Y(csr_n275) );
  OA222X1_LVT csr_U364 ( .A1(n_T_1165[55]), .A2(csr_io_rw_rdata[55]), .A3(
        n_T_1165[55]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n274), .Y(
        csr_wdata_55_) );
  INVX0_LVT csr_U363 ( .A(n_T_1165[55]), .Y(csr_n274) );
  AO22X1_LVT csr_U362 ( .A1(csr_n497), .A2(csr_n_T_52[52]), .A3(csr_wdata_58_), 
        .A4(csr_n1149), .Y(csr_N1943) );
  OA222X1_LVT csr_U361 ( .A1(io_imem_sfence_bits_addr[17]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[17]), .A4(csr_io_rw_rdata[17]), .A5(
        csr_n516), .A6(csr_n273), .Y(csr_wdata_17_) );
  INVX0_LVT csr_U360 ( .A(io_imem_sfence_bits_addr[17]), .Y(csr_n273) );
  NAND3X0_LVT csr_U359 ( .A1(csr_n271), .A2(csr_n917), .A3(csr_n272), .Y(
        csr_n1914) );
  NAND2X0_LVT csr_U358 ( .A1(csr_n1935), .A2(csr_n1443), .Y(csr_n272) );
  NAND2X0_LVT csr_U357 ( .A1(csr_wdata_5_), .A2(csr_n949), .Y(csr_n271) );
  AND4X1_LVT csr_U356 ( .A1(csr_io_rw_addr[0]), .A2(csr_io_rw_addr[1]), .A3(
        csr_n616), .A4(csr_io_rw_addr[2]), .Y(csr_n1479) );
  AO22X1_LVT csr_U355 ( .A1(csr_n1508), .A2(csr_reg_sscratch[31]), .A3(
        csr_n1162), .A4(csr_io_time[31]), .Y(csr_n268) );
  AO22X1_LVT csr_U353 ( .A1(csr_n1493), .A2(csr_reg_dpc_31_), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_31_), .Y(csr_n265) );
  AO22X1_LVT csr_U352 ( .A1(csr_n1489), .A2(csr_reg_mepc_31_), .A3(csr_n1506), 
        .A4(csr_reg_sepc_31_), .Y(csr_n264) );
  AO22X1_LVT csr_U351 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[31]), .A3(
        csr_n1487), .A4(csr_reg_stvec_31_), .Y(csr_n263) );
  AO22X1_LVT csr_U350 ( .A1(csr_n1160), .A2(csr_n_T_444[31]), .A3(csr_n1153), 
        .A4(csr_n_T_383[31]), .Y(csr_n262) );
  NAND4X0_LVT csr_U349 ( .A1(csr_n248), .A2(csr_n249), .A3(csr_n250), .A4(
        csr_n261), .Y(csr_io_rw_rdata[28]) );
  NOR4X0_LVT csr_U348 ( .A1(csr_n251), .A2(csr_n252), .A3(csr_n253), .A4(
        csr_n260), .Y(csr_n261) );
  AO22X1_LVT csr_U347 ( .A1(csr_n1162), .A2(csr_io_time[28]), .A3(csr_n1160), 
        .A4(csr_n_T_444[28]), .Y(csr_n259) );
  AO22X1_LVT csr_U345 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[28]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[28]), .Y(csr_n256) );
  AO21X1_LVT csr_U344 ( .A1(csr_n1493), .A2(csr_reg_dpc_28_), .A3(csr_n254), 
        .Y(csr_n255) );
  AO222X1_LVT csr_U343 ( .A1(csr_n1689), .A2(csr_n_T_45_28_), .A3(csr_n1506), 
        .A4(csr_reg_sepc_28_), .A5(csr_n1489), .A6(csr_reg_mepc_28_), .Y(
        csr_n254) );
  AO22X1_LVT csr_U342 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[28]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[28]), .Y(csr_n253) );
  AO22X1_LVT csr_U341 ( .A1(csr_n1510), .A2(csr_reg_dscratch[28]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[28]), .Y(csr_n252) );
  AO22X1_LVT csr_U340 ( .A1(csr_n1508), .A2(csr_reg_sscratch[28]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[28]), .Y(csr_n251) );
  AOI22X1_LVT csr_U339 ( .A1(csr_n1485), .A2(csr_reg_mscratch[28]), .A3(
        csr_n1487), .A4(csr_reg_stvec_28_), .Y(csr_n250) );
  AOI22X1_LVT csr_U338 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[28]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[28]), .Y(csr_n249) );
  AOI22X1_LVT csr_U337 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[28]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_28_), .Y(csr_n248) );
  NAND2X0_LVT csr_U336 ( .A1(csr_n239), .A2(csr_n247), .Y(csr_io_rw_rdata[26])
         );
  NOR4X0_LVT csr_U335 ( .A1(csr_n240), .A2(csr_n244), .A3(csr_n245), .A4(
        csr_n246), .Y(csr_n247) );
  AO22X1_LVT csr_U334 ( .A1(csr_n1506), .A2(csr_reg_sepc_26_), .A3(csr_n1490), 
        .A4(csr_io_bp_0_address[26]), .Y(csr_n246) );
  AO22X1_LVT csr_U333 ( .A1(csr_n1162), .A2(csr_io_time[26]), .A3(csr_n1496), 
        .A4(io_ptw_pmp_1_addr[26]), .Y(csr_n245) );
  AO22X1_LVT csr_U331 ( .A1(csr_n1153), .A2(csr_n_T_383[26]), .A3(csr_n1479), 
        .A4(io_ptw_pmp_7_addr[26]), .Y(csr_n242) );
  AO222X1_LVT csr_U330 ( .A1(csr_n1689), .A2(csr_n_T_45_26_), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_26_), .A5(csr_reg_dpc_26_), .A6(csr_n1493), .Y(
        csr_n241) );
  AO222X1_LVT csr_U329 ( .A1(csr_n1489), .A2(csr_reg_mepc_26_), .A3(csr_n1492), 
        .A4(io_ptw_pmp_2_addr[26]), .A5(csr_n1487), .A6(csr_reg_stvec_26_), 
        .Y(csr_n240) );
  NOR4X0_LVT csr_U328 ( .A1(csr_n235), .A2(csr_n236), .A3(csr_n237), .A4(
        csr_n238), .Y(csr_n239) );
  AO22X1_LVT csr_U327 ( .A1(csr_n1507), .A2(io_ptw_pmp_3_cfg_x), .A3(csr_n1472), .A4(io_ptw_pmp_5_addr[26]), .Y(csr_n238) );
  AO22X1_LVT csr_U326 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[26]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[26]), .Y(csr_n237) );
  AO22X1_LVT csr_U325 ( .A1(csr_n1485), .A2(csr_reg_mscratch[26]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[26]), .Y(csr_n236) );
  AO222X1_LVT csr_U324 ( .A1(csr_n1508), .A2(csr_reg_sscratch[26]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[26]), .A5(csr_n1160), .A6(
        csr_n_T_444[26]), .Y(csr_n235) );
  OA222X1_LVT csr_U323 ( .A1(n_T_1165[45]), .A2(csr_io_rw_rdata[45]), .A3(
        n_T_1165[45]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n234), .Y(
        csr_wdata_45_) );
  INVX0_LVT csr_U322 ( .A(n_T_1165[45]), .Y(csr_n234) );
  OA222X1_LVT csr_U321 ( .A1(n_T_1165[40]), .A2(csr_io_rw_rdata[40]), .A3(
        n_T_1165[40]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n233), .Y(
        csr_wdata_40_) );
  INVX0_LVT csr_U320 ( .A(n_T_1165[40]), .Y(csr_n233) );
  OA222X1_LVT csr_U319 ( .A1(csr_n232), .A2(wb_ctrl_csr[1]), .A3(csr_n232), 
        .A4(csr_io_rw_rdata[5]), .A5(csr_n516), .A6(csr_n1904), .Y(
        csr_wdata_5_) );
  INVX0_LVT csr_U318 ( .A(csr_n1904), .Y(csr_n232) );
  OR3X1_LVT csr_U317 ( .A1(csr_n223), .A2(csr_n230), .A3(csr_n231), .Y(
        csr_io_rw_rdata[33]) );
  AO22X1_LVT csr_U316 ( .A1(csr_n1508), .A2(csr_reg_sscratch[33]), .A3(
        csr_n1507), .A4(io_ptw_pmp_4_cfg_w), .Y(csr_n231) );
  NAND4X0_LVT csr_U314 ( .A1(csr_n1026), .A2(csr_n225), .A3(csr_n226), .A4(
        csr_n227), .Y(csr_n228) );
  AOI22X1_LVT csr_U313 ( .A1(csr_n1153), .A2(csr_n_T_383[33]), .A3(csr_n1487), 
        .A4(csr_reg_stvec_33_), .Y(csr_n227) );
  AOI22X1_LVT csr_U312 ( .A1(csr_n1493), .A2(csr_reg_dpc_33_), .A3(csr_n1490), 
        .A4(csr_io_bp_0_address[33]), .Y(csr_n226) );
  AOI22X1_LVT csr_U311 ( .A1(csr_n1510), .A2(csr_reg_dscratch[33]), .A3(
        csr_n1689), .A4(csr_n_T_45_33_), .Y(csr_n225) );
  AO22X1_LVT csr_U310 ( .A1(csr_n1162), .A2(csr_n1966), .A3(csr_n1506), .A4(
        csr_reg_sepc_33_), .Y(csr_n224) );
  AO22X1_LVT csr_U309 ( .A1(csr_n1485), .A2(csr_reg_mscratch[33]), .A3(
        csr_n1489), .A4(csr_reg_mepc_33_), .Y(csr_n223) );
  NAND4X0_LVT csr_U308 ( .A1(csr_n214), .A2(csr_n219), .A3(csr_n220), .A4(
        csr_n222), .Y(csr_io_rw_rdata[10]) );
  AOI21X1_LVT csr_U307 ( .A1(csr_n1487), .A2(csr_reg_stvec_10_), .A3(csr_n221), 
        .Y(csr_n222) );
  AO22X1_LVT csr_U306 ( .A1(csr_n1508), .A2(csr_reg_sscratch[10]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_10_), .Y(csr_n221) );
  AOI22X1_LVT csr_U305 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[10]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[10]), .Y(csr_n220) );
  NOR4X0_LVT csr_U304 ( .A1(csr_n215), .A2(csr_n216), .A3(csr_n217), .A4(
        csr_n218), .Y(csr_n219) );
  AO222X1_LVT csr_U303 ( .A1(csr_n1485), .A2(csr_reg_mscratch[10]), .A3(
        csr_n488), .A4(io_ptw_ptbr_ppn[10]), .A5(csr_n1160), .A6(
        csr_n_T_444[10]), .Y(csr_n218) );
  AO22X1_LVT csr_U302 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[10]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[10]), .Y(csr_n217) );
  AO222X1_LVT csr_U301 ( .A1(csr_n1489), .A2(csr_reg_mepc_10_), .A3(csr_n1473), 
        .A4(io_ptw_pmp_3_addr[10]), .A5(io_ptw_pmp_1_addr[10]), .A6(csr_n1496), 
        .Y(csr_n216) );
  AO22X1_LVT csr_U300 ( .A1(csr_n1689), .A2(csr_n_T_45_10_), .A3(csr_n1153), 
        .A4(csr_n_T_383[10]), .Y(csr_n215) );
  NOR4X0_LVT csr_U299 ( .A1(csr_n210), .A2(csr_n211), .A3(csr_n212), .A4(
        csr_n213), .Y(csr_n214) );
  AO22X1_LVT csr_U298 ( .A1(csr_n1510), .A2(csr_reg_dscratch[10]), .A3(
        csr_n1493), .A4(csr_reg_dpc_10_), .Y(csr_n213) );
  AO22X1_LVT csr_U297 ( .A1(csr_n1162), .A2(csr_io_time[10]), .A3(csr_n1472), 
        .A4(io_ptw_pmp_5_addr[10]), .Y(csr_n212) );
  AO22X1_LVT csr_U296 ( .A1(csr_n1507), .A2(io_ptw_pmp_1_cfg_x), .A3(csr_n1506), .A4(csr_reg_sepc_10_), .Y(csr_n211) );
  AO22X1_LVT csr_U295 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[10]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[10]), .Y(csr_n210) );
  NAND3X0_LVT csr_U294 ( .A1(csr_n209), .A2(csr_n208), .A3(csr_n1186), .Y(
        csr_io_interrupt_cause[3]) );
  OR2X1_LVT csr_U293 ( .A1(csr_n1187), .A2(csr_n1188), .Y(csr_n209) );
  NAND3X0_LVT csr_U292 ( .A1(csr_n1192), .A2(csr_n1193), .A3(csr_n207), .Y(
        csr_n208) );
  AO21X1_LVT csr_U291 ( .A1(csr_n1191), .A2(csr_n1190), .A3(csr_n1189), .Y(
        csr_n207) );
  OAI22X1_LVT csr_U290 ( .A1(csr_n701), .A2(csr_n1483), .A3(csr_n899), .A4(
        csr_n206), .Y(csr_N883) );
  INVX0_LVT csr_U289 ( .A(csr_n1498), .Y(csr_n206) );
  OA222X1_LVT csr_U288 ( .A1(n_T_1165[44]), .A2(csr_io_rw_rdata[44]), .A3(
        n_T_1165[44]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n205), .Y(
        csr_wdata_44_) );
  INVX0_LVT csr_U287 ( .A(n_T_1165[44]), .Y(csr_n205) );
  OA222X1_LVT csr_U286 ( .A1(n_T_1165[41]), .A2(csr_io_rw_rdata[41]), .A3(
        n_T_1165[41]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n204), .Y(
        csr_wdata_41_) );
  INVX0_LVT csr_U285 ( .A(n_T_1165[41]), .Y(csr_n204) );
  AO22X1_LVT csr_U284 ( .A1(csr_n497), .A2(csr_n_T_52[44]), .A3(csr_wdata_50_), 
        .A4(csr_n1149), .Y(csr_N1935) );
  OA222X1_LVT csr_U283 ( .A1(io_imem_sfence_bits_addr[25]), .A2(
        csr_io_rw_rdata[25]), .A3(io_imem_sfence_bits_addr[25]), .A4(
        wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n203), .Y(csr_wdata_25_) );
  INVX0_LVT csr_U282 ( .A(io_imem_sfence_bits_addr[25]), .Y(csr_n203) );
  AND3X1_LVT csr_U281 ( .A1(csr_io_rw_addr[6]), .A2(csr_n1515), .A3(csr_n1527), 
        .Y(csr_n1509) );
  OR3X1_LVT csr_U280 ( .A1(csr_n190), .A2(csr_n201), .A3(csr_n202), .Y(
        csr_io_rw_rdata[35]) );
  AO22X1_LVT csr_U279 ( .A1(csr_n1508), .A2(csr_reg_sscratch[35]), .A3(
        csr_n1506), .A4(csr_reg_sepc_35_), .Y(csr_n202) );
  NAND4X0_LVT csr_U277 ( .A1(csr_n192), .A2(csr_n1041), .A3(csr_n193), .A4(
        csr_n195), .Y(csr_n196) );
  NAND2X0_LVT csr_U276 ( .A1(csr_n1493), .A2(csr_reg_dpc_35_), .Y(csr_n195) );
  AOI22X1_LVT csr_U275 ( .A1(csr_n1507), .A2(io_ptw_pmp_4_cfg_a[0]), .A3(
        csr_n1490), .A4(csr_io_bp_0_address[35]), .Y(csr_n193) );
  AOI22X1_LVT csr_U274 ( .A1(csr_n1510), .A2(csr_reg_dscratch[35]), .A3(
        csr_n1689), .A4(csr_n_T_45_35_), .Y(csr_n192) );
  AO22X1_LVT csr_U273 ( .A1(csr_n1162), .A2(csr_n1964), .A3(csr_n1153), .A4(
        csr_n_T_383[35]), .Y(csr_n191) );
  AO222X1_LVT csr_U272 ( .A1(csr_n1485), .A2(csr_reg_mscratch[35]), .A3(
        csr_n1489), .A4(csr_reg_mepc_35_), .A5(csr_n_T_444[35]), .A6(csr_n1160), .Y(csr_n190) );
  NAND2X0_LVT csr_U271 ( .A1(csr_n184), .A2(csr_n189), .Y(csr_io_rw_rdata[15])
         );
  NOR4X0_LVT csr_U270 ( .A1(csr_n185), .A2(csr_n186), .A3(csr_n187), .A4(
        csr_n188), .Y(csr_n189) );
  AO22X1_LVT csr_U269 ( .A1(csr_n1510), .A2(csr_reg_dscratch[15]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[15]), .Y(csr_n188) );
  AO22X1_LVT csr_U268 ( .A1(csr_n1508), .A2(csr_reg_sscratch[15]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[15]), .Y(csr_n187) );
  AO22X1_LVT csr_U267 ( .A1(csr_n1489), .A2(csr_reg_mepc_15_), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_15_), .Y(csr_n186) );
  AO22X1_LVT csr_U266 ( .A1(csr_n1153), .A2(csr_n_T_383[15]), .A3(csr_n1494), 
        .A4(io_ptw_pmp_6_addr[15]), .Y(csr_n185) );
  NOR4X0_LVT csr_U265 ( .A1(csr_n175), .A2(csr_n176), .A3(csr_n182), .A4(
        csr_n183), .Y(csr_n184) );
  AO22X1_LVT csr_U264 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[15]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[15]), .Y(csr_n183) );
  AO22X1_LVT csr_U263 ( .A1(csr_n1162), .A2(csr_io_time[15]), .A3(csr_n1490), 
        .A4(csr_io_bp_0_address[15]), .Y(csr_n181) );
  NAND3X0_LVT csr_U261 ( .A1(csr_n177), .A2(csr_n631), .A3(csr_n632), .Y(
        csr_n178) );
  AOI22X1_LVT csr_U260 ( .A1(csr_n1495), .A2(csr_n_T_1155_3), .A3(csr_n1488), 
        .A4(io_ptw_ptbr_ppn[15]), .Y(csr_n177) );
  AO22X1_LVT csr_U259 ( .A1(csr_n1491), .A2(io_ptw_pmp_4_addr[15]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[15]), .Y(csr_n176) );
  AO222X1_LVT csr_U258 ( .A1(csr_n1160), .A2(csr_n_T_444[15]), .A3(csr_n1480), 
        .A4(io_ptw_pmp_0_addr[15]), .A5(io_ptw_pmp_5_addr[15]), .A6(csr_n1472), 
        .Y(csr_n175) );
  NAND3X0_LVT csr_U257 ( .A1(csr_n174), .A2(csr_n590), .A3(csr_n173), .Y(
        csr_N334) );
  OR2X1_LVT csr_U256 ( .A1(csr_n931), .A2(csr_n367), .Y(csr_n174) );
  AOI22X1_LVT csr_U255 ( .A1(csr_n_1929_), .A2(csr_n930), .A3(
        io_ptw_status_prv[1]), .A4(csr_n929), .Y(csr_n173) );
  OA222X1_LVT csr_U254 ( .A1(n_T_1165[62]), .A2(csr_n589), .A3(n_T_1165[62]), 
        .A4(csr_io_rw_rdata[62]), .A5(csr_n516), .A6(csr_n172), .Y(
        csr_wdata_62_) );
  INVX0_LVT csr_U253 ( .A(n_T_1165[62]), .Y(csr_n172) );
  OA222X1_LVT csr_U252 ( .A1(n_T_1165[48]), .A2(csr_io_rw_rdata[48]), .A3(
        n_T_1165[48]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n171), .Y(
        csr_wdata_48_) );
  INVX0_LVT csr_U251 ( .A(n_T_1165[48]), .Y(csr_n171) );
  AO22X1_LVT csr_U250 ( .A1(csr_n494), .A2(csr_n_T_44[32]), .A3(csr_wdata_38_), 
        .A4(csr_n1128), .Y(csr_N1529) );
  AO22X1_LVT csr_U249 ( .A1(csr_n1446), .A2(csr_n170), .A3(csr_wdata_1_), .A4(
        csr_n1149), .Y(csr_N1823) );
  OA221X1_LVT csr_U248 ( .A1(csr_io_time[1]), .A2(csr_io_time[0]), .A3(
        csr_io_time[1]), .A4(csr_n168), .A5(csr_n169), .Y(csr_n170) );
  INVX0_LVT csr_U247 ( .A(csr_n1142), .Y(csr_n169) );
  INVX0_LVT csr_U246 ( .A(csr_io_csr_stall), .Y(csr_n168) );
  NAND4X0_LVT csr_U245 ( .A1(csr_n155), .A2(csr_n156), .A3(csr_n157), .A4(
        csr_n167), .Y(csr_io_rw_rdata[25]) );
  NOR4X0_LVT csr_U244 ( .A1(csr_n158), .A2(csr_n159), .A3(csr_n160), .A4(
        csr_n166), .Y(csr_n167) );
  AO22X1_LVT csr_U242 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[25]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[25]), .Y(csr_n164) );
  AO21X1_LVT csr_U241 ( .A1(csr_n1487), .A2(csr_reg_stvec_25_), .A3(csr_n162), 
        .Y(csr_n163) );
  AO21X1_LVT csr_U240 ( .A1(csr_n1510), .A2(csr_reg_dscratch[25]), .A3(
        csr_n161), .Y(csr_n162) );
  AO222X1_LVT csr_U239 ( .A1(csr_n1689), .A2(csr_n_T_45_25_), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_25_), .A5(csr_reg_dpc_25_), .A6(csr_n1493), .Y(
        csr_n161) );
  AO222X1_LVT csr_U238 ( .A1(csr_n1507), .A2(io_ptw_pmp_3_cfg_w), .A3(
        csr_n1496), .A4(io_ptw_pmp_1_addr[25]), .A5(csr_n1160), .A6(
        csr_n_T_444[25]), .Y(csr_n160) );
  AO22X1_LVT csr_U237 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[25]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[25]), .Y(csr_n159) );
  AO22X1_LVT csr_U236 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[25]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[25]), .Y(csr_n158) );
  AOI22X1_LVT csr_U235 ( .A1(csr_n1508), .A2(csr_reg_sscratch[25]), .A3(
        csr_n1485), .A4(csr_reg_mscratch[25]), .Y(csr_n157) );
  AOI22X1_LVT csr_U234 ( .A1(csr_n1162), .A2(csr_io_time[25]), .A3(csr_n1494), 
        .A4(io_ptw_pmp_6_addr[25]), .Y(csr_n156) );
  AOI222X1_LVT csr_U233 ( .A1(csr_n1489), .A2(csr_reg_mepc_25_), .A3(csr_n1506), .A4(csr_reg_sepc_25_), .A5(csr_n1491), .A6(io_ptw_pmp_4_addr[25]), .Y(
        csr_n155) );
  AO22X1_LVT csr_U232 ( .A1(csr_n1443), .A2(csr_n154), .A3(csr_n949), .A4(
        csr_wdata_8_), .Y(csr_n1913) );
  AND2X1_LVT csr_U231 ( .A1(io_ptw_status_prv[0]), .A2(csr_n501), .Y(csr_n154)
         );
  OA222X1_LVT csr_U230 ( .A1(n_T_1165[39]), .A2(csr_io_rw_rdata[39]), .A3(
        n_T_1165[39]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n153), .Y(
        csr_wdata_39_) );
  INVX0_LVT csr_U229 ( .A(n_T_1165[39]), .Y(csr_n153) );
  OA222X1_LVT csr_U228 ( .A1(n_T_1165[49]), .A2(csr_io_rw_rdata[49]), .A3(
        n_T_1165[49]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n152), .Y(
        csr_wdata_49_) );
  INVX0_LVT csr_U227 ( .A(n_T_1165[49]), .Y(csr_n152) );
  AO22X1_LVT csr_U226 ( .A1(csr_wdata_9_), .A2(csr_n150), .A3(csr_n446), .A4(
        csr_n151), .Y(csr_N615) );
  INVX0_LVT csr_U225 ( .A(csr_n742), .Y(csr_n151) );
  AO21X1_LVT csr_U224 ( .A1(csr_read_mideleg_9_), .A2(csr_n1504), .A3(
        csr_n1502), .Y(csr_n150) );
  AND2X1_LVT csr_U223 ( .A1(csr_n149), .A2(csr_n1176), .Y(csr_n1180) );
  INVX0_LVT csr_U222 ( .A(csr_n1183), .Y(csr_n149) );
  NAND4X0_LVT csr_U221 ( .A1(csr_n131), .A2(csr_n136), .A3(csr_n147), .A4(
        csr_n148), .Y(csr_io_rw_rdata[4]) );
  NAND2X0_LVT csr_U220 ( .A1(csr_n1470), .A2(csr_reg_mtvec_4_), .Y(csr_n148)
         );
  NOR4X0_LVT csr_U219 ( .A1(csr_n137), .A2(csr_n138), .A3(csr_n139), .A4(
        csr_n146), .Y(csr_n147) );
  OR3X1_LVT csr_U218 ( .A1(csr_n140), .A2(csr_n141), .A3(csr_n145), .Y(
        csr_n146) );
  AO22X1_LVT csr_U216 ( .A1(csr_n1506), .A2(csr_reg_sepc_4_), .A3(csr_n1481), 
        .A4(csr_io_bp_0_control_s), .Y(csr_n143) );
  AO222X1_LVT csr_U215 ( .A1(csr_n1510), .A2(csr_reg_dscratch[4]), .A3(
        csr_n1507), .A4(io_ptw_pmp_0_cfg_a[1]), .A5(csr_n_T_45_4_), .A6(
        csr_n1689), .Y(csr_n142) );
  AO22X1_LVT csr_U214 ( .A1(csr_n1489), .A2(csr_reg_mepc_4_), .A3(csr_n1496), 
        .A4(io_ptw_pmp_1_addr[4]), .Y(csr_n141) );
  AO22X1_LVT csr_U213 ( .A1(csr_n1160), .A2(csr_n_T_444[4]), .A3(csr_n1153), 
        .A4(csr_n_T_383[4]), .Y(csr_n140) );
  AO22X1_LVT csr_U212 ( .A1(csr_n1508), .A2(csr_reg_sscratch[4]), .A3(
        csr_n1472), .A4(io_ptw_pmp_5_addr[4]), .Y(csr_n139) );
  AO22X1_LVT csr_U211 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[4]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[4]), .Y(csr_n138) );
  AO22X1_LVT csr_U210 ( .A1(csr_n1473), .A2(io_ptw_pmp_3_addr[4]), .A3(
        csr_n1488), .A4(io_ptw_ptbr_ppn[4]), .Y(csr_n137) );
  NOR4X0_LVT csr_U209 ( .A1(csr_n132), .A2(csr_n133), .A3(csr_n134), .A4(
        csr_n135), .Y(csr_n136) );
  AO22X1_LVT csr_U208 ( .A1(csr_n1485), .A2(csr_reg_mscratch[4]), .A3(
        csr_n1469), .A4(csr_read_medeleg_4_), .Y(csr_n135) );
  AO22X1_LVT csr_U207 ( .A1(csr_n1493), .A2(csr_reg_dpc_4_), .A3(csr_n1480), 
        .A4(io_ptw_pmp_0_addr[4]), .Y(csr_n134) );
  AO22X1_LVT csr_U206 ( .A1(csr_n1162), .A2(csr_io_time[4]), .A3(csr_n1491), 
        .A4(io_ptw_pmp_4_addr[4]), .Y(csr_n133) );
  AO22X1_LVT csr_U205 ( .A1(csr_n1168), .A2(csr_reg_scause[4]), .A3(csr_n1478), 
        .A4(csr_reg_stvec_4_), .Y(csr_n132) );
  AOI22X1_LVT csr_U204 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[4]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[4]), .Y(csr_n131) );
  OA222X1_LVT csr_U203 ( .A1(csr_n130), .A2(csr_io_rw_rdata[9]), .A3(csr_n130), 
        .A4(csr_n589), .A5(csr_n516), .A6(csr_n1907), .Y(csr_wdata_9_) );
  INVX0_LVT csr_U202 ( .A(csr_n1907), .Y(csr_n130) );
  OAI222X1_LVT csr_U201 ( .A1(csr_n128), .A2(csr_n954), .A3(csr_n129), .A4(
        csr_n1455), .A5(csr_n953), .A6(csr_n1697), .Y(csr_N1270) );
  INVX0_LVT csr_U200 ( .A(csr_wdata_0_), .Y(csr_n129) );
  INVX0_LVT csr_U199 ( .A(csr_n1500), .Y(csr_n128) );
  OA222X1_LVT csr_U198 ( .A1(n_T_1165[50]), .A2(csr_io_rw_rdata[50]), .A3(
        n_T_1165[50]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n127), .Y(
        csr_wdata_50_) );
  INVX0_LVT csr_U197 ( .A(n_T_1165[50]), .Y(csr_n127) );
  OA222X1_LVT csr_U196 ( .A1(n_T_1165[63]), .A2(csr_io_rw_rdata[63]), .A3(
        n_T_1165[63]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n126), .Y(
        csr_wdata_63_) );
  INVX0_LVT csr_U195 ( .A(n_T_1165[63]), .Y(csr_n126) );
  AO22X1_LVT csr_U194 ( .A1(csr_n492), .A2(csr_wdata_3_), .A3(csr_n124), .A4(
        csr_n125), .Y(csr_N1431) );
  INVX0_LVT csr_U193 ( .A(csr_n960), .Y(csr_n125) );
  OA21X1_LVT csr_U192 ( .A1(csr_n959), .A2(csr_n_T_45_3_), .A3(csr_n961), .Y(
        csr_n124) );
  AND3X1_LVT csr_U191 ( .A1(csr_n1516), .A2(csr_n1512), .A3(csr_n1527), .Y(
        csr_n1154) );
  AND3X1_LVT csr_U190 ( .A1(csr_io_time[3]), .A2(csr_io_time[4]), .A3(
        csr_n1144), .Y(csr_n1147) );
  OA221X1_LVT csr_U189 ( .A1(io_imem_sfence_bits_addr[12]), .A2(csr_n122), 
        .A3(csr_n123), .A4(csr_n516), .A5(csr_n1482), .Y(csr_N485) );
  INVX0_LVT csr_U188 ( .A(io_imem_sfence_bits_addr[12]), .Y(csr_n123) );
  AND2X1_LVT csr_U187 ( .A1(csr_io_bp_0_control_action), .A2(csr_n589), .Y(
        csr_n122) );
  AO22X1_LVT csr_U186 ( .A1(csr_n494), .A2(csr_n_T_44[44]), .A3(csr_wdata_50_), 
        .A4(csr_n1128), .Y(csr_N1541) );
  AO22X1_LVT csr_U185 ( .A1(csr_n497), .A2(csr_n_T_52[32]), .A3(csr_wdata_38_), 
        .A4(csr_n1149), .Y(csr_N1923) );
  AND3X1_LVT csr_U184 ( .A1(csr_n1516), .A2(csr_n1505), .A3(csr_n1527), .Y(
        csr_n1504) );
  AO21X1_LVT csr_U183 ( .A1(csr_n502), .A2(csr_reg_mepc_36_), .A3(csr_n121), 
        .Y(csr_io_evec[36]) );
  AO222X1_LVT csr_U182 ( .A1(csr_n500), .A2(csr_reg_sepc_36_), .A3(csr_n499), 
        .A4(csr_reg_stvec_36_), .A5(csr_n1356), .A6(csr_reg_dpc_36_), .Y(
        csr_n121) );
  NAND3X0_LVT csr_U181 ( .A1(csr_n1480), .A2(csr_n453), .A3(csr_n120), .Y(
        csr_n430) );
  NAND3X0_LVT csr_U180 ( .A1(io_ptw_pmp_1_cfg_a[0]), .A2(csr_n462), .A3(
        io_ptw_pmp_1_cfg_l), .Y(csr_n120) );
  NAND3X0_LVT csr_U179 ( .A1(csr_n1491), .A2(csr_n438), .A3(csr_n119), .Y(
        csr_n433) );
  NAND3X0_LVT csr_U178 ( .A1(io_ptw_pmp_5_cfg_a[0]), .A2(csr_n461), .A3(
        io_ptw_pmp_5_cfg_l), .Y(csr_n119) );
  NAND3X0_LVT csr_U177 ( .A1(csr_n1494), .A2(csr_n439), .A3(csr_n118), .Y(
        csr_n435) );
  NAND3X0_LVT csr_U176 ( .A1(io_ptw_pmp_7_cfg_l), .A2(csr_n459), .A3(
        io_ptw_pmp_7_cfg_a[0]), .Y(csr_n118) );
  NAND3X0_LVT csr_U175 ( .A1(csr_n1492), .A2(csr_n441), .A3(csr_n117), .Y(
        csr_n432) );
  NAND3X0_LVT csr_U174 ( .A1(io_ptw_pmp_3_cfg_a[0]), .A2(csr_n460), .A3(
        io_ptw_pmp_3_cfg_l), .Y(csr_n117) );
  NAND3X0_LVT csr_U173 ( .A1(ibuf_io_inst_0_bits_raw[26]), .A2(csr_n1386), 
        .A3(csr_n116), .Y(csr_n1426) );
  INVX0_LVT csr_U172 ( .A(csr_n1375), .Y(csr_n116) );
  AO22X1_LVT csr_U171 ( .A1(csr_n492), .A2(csr_wdata_0_), .A3(csr_n115), .A4(
        csr_n961), .Y(csr_N1428) );
  HADDX1_LVT csr_U170 ( .A0(csr_io_retire), .B0(csr_n_T_45_0_), .SO(csr_n115)
         );
  OA222X1_LVT csr_U169 ( .A1(n_T_1165[52]), .A2(csr_io_rw_rdata[52]), .A3(
        n_T_1165[52]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n114), .Y(
        csr_wdata_52_) );
  INVX0_LVT csr_U168 ( .A(n_T_1165[52]), .Y(csr_n114) );
  OA222X1_LVT csr_U167 ( .A1(n_T_1165[60]), .A2(csr_n589), .A3(n_T_1165[60]), 
        .A4(csr_io_rw_rdata[60]), .A5(csr_n516), .A6(csr_n113), .Y(
        csr_wdata_60_) );
  INVX0_LVT csr_U166 ( .A(n_T_1165[60]), .Y(csr_n113) );
  OA222X1_LVT csr_U165 ( .A1(io_imem_sfence_bits_addr[11]), .A2(csr_n589), 
        .A3(io_imem_sfence_bits_addr[11]), .A4(csr_io_rw_rdata[11]), .A5(
        csr_n516), .A6(csr_n112), .Y(csr_wdata_11_) );
  INVX0_LVT csr_U164 ( .A(io_imem_sfence_bits_addr[11]), .Y(csr_n112) );
  OR2X1_LVT csr_U163 ( .A1(csr_n1191), .A2(csr_n111), .Y(csr_n1194) );
  NAND4X0_LVT csr_U162 ( .A1(csr_n1185), .A2(csr_n1192), .A3(csr_n1174), .A4(
        csr_n110), .Y(csr_n111) );
  AO22X1_LVT csr_U161 ( .A1(csr_n1179), .A2(csr_n1178), .A3(csr_n1190), .A4(
        csr_n109), .Y(csr_n110) );
  INVX0_LVT csr_U160 ( .A(csr_n1175), .Y(csr_n109) );
  NAND3X0_LVT csr_U159 ( .A1(csr_n1473), .A2(csr_n443), .A3(csr_n108), .Y(
        csr_n436) );
  NAND3X0_LVT csr_U158 ( .A1(io_ptw_pmp_4_cfg_l), .A2(csr_n464), .A3(
        io_ptw_pmp_4_cfg_a[0]), .Y(csr_n108) );
  NAND3X0_LVT csr_U157 ( .A1(csr_n1083), .A2(csr_n106), .A3(csr_n107), .Y(
        csr_n669) );
  AOI22X1_LVT csr_U156 ( .A1(csr_n1689), .A2(csr_n_T_45_12_), .A3(csr_n1495), 
        .A4(csr_n_T_1155_0_), .Y(csr_n107) );
  AOI22X1_LVT csr_U155 ( .A1(csr_n1487), .A2(csr_reg_stvec_12_), .A3(csr_n1469), .A4(csr_read_medeleg_12), .Y(csr_n106) );
  NAND3X0_LVT csr_U154 ( .A1(csr_n1405), .A2(ibuf_io_inst_0_bits_raw[28]), 
        .A3(csr_n105), .Y(csr_n1375) );
  INVX0_LVT csr_U153 ( .A(csr_n1378), .Y(csr_n105) );
  OA21X1_LVT csr_U152 ( .A1(csr_io_retire), .A2(csr_n104), .A3(
        csr_io_singleStep), .Y(csr_N435) );
  NAND2X0_LVT csr_U151 ( .A1(csr_n860), .A2(csr_n1442), .Y(csr_n104) );
  OA222X1_LVT csr_U150 ( .A1(n_T_1165[51]), .A2(csr_io_rw_rdata[51]), .A3(
        n_T_1165[51]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n103), .Y(
        csr_wdata_51_) );
  INVX0_LVT csr_U149 ( .A(n_T_1165[51]), .Y(csr_n103) );
  OA222X1_LVT csr_U148 ( .A1(n_T_1165[59]), .A2(csr_io_rw_rdata[59]), .A3(
        n_T_1165[59]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n102), .Y(
        csr_wdata_59_) );
  INVX0_LVT csr_U147 ( .A(n_T_1165[59]), .Y(csr_n102) );
  OA222X1_LVT csr_U146 ( .A1(io_imem_sfence_bits_addr[3]), .A2(csr_n589), .A3(
        io_imem_sfence_bits_addr[3]), .A4(csr_io_rw_rdata[3]), .A5(csr_n516), 
        .A6(csr_n101), .Y(csr_wdata_3_) );
  INVX0_LVT csr_U145 ( .A(io_imem_sfence_bits_addr[3]), .Y(csr_n101) );
  OA222X1_LVT csr_U144 ( .A1(csr_n99), .A2(csr_n1912), .A3(csr_n99), .A4(
        csr_n590), .A5(csr_n879), .A6(csr_n100), .Y(csr_n1911) );
  INVX0_LVT csr_U143 ( .A(csr_wdata_9_), .Y(csr_n100) );
  INVX0_LVT csr_U142 ( .A(csr_n879), .Y(csr_n99) );
  OR3X1_LVT csr_U141 ( .A1(csr_n82), .A2(csr_n83), .A3(csr_n98), .Y(
        csr_io_rw_rdata[12]) );
  OR3X1_LVT csr_U140 ( .A1(csr_n84), .A2(csr_n85), .A3(csr_n97), .Y(csr_n98)
         );
  OR3X1_LVT csr_U139 ( .A1(csr_n86), .A2(csr_n90), .A3(csr_n96), .Y(csr_n97)
         );
  AO22X1_LVT csr_U138 ( .A1(csr_n1485), .A2(csr_reg_mscratch[12]), .A3(
        csr_n1157), .A4(csr_n_1929_), .Y(csr_n94) );
  AO22X1_LVT csr_U137 ( .A1(csr_n1481), .A2(csr_io_bp_0_control_action), .A3(
        csr_n1452), .A4(csr_io_status_isa_12_), .Y(csr_n92) );
  AO22X1_LVT csr_U136 ( .A1(csr_n1506), .A2(csr_reg_sepc_12_), .A3(csr_n1473), 
        .A4(io_ptw_pmp_3_addr[12]), .Y(csr_n91) );
  AO22X1_LVT csr_U134 ( .A1(csr_n1510), .A2(csr_reg_dscratch[12]), .A3(
        csr_n1488), .A4(io_ptw_ptbr_ppn[12]), .Y(csr_n88) );
  AO22X1_LVT csr_U133 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[12]), .A3(
        csr_n1491), .A4(io_ptw_pmp_4_addr[12]), .Y(csr_n87) );
  AO22X1_LVT csr_U132 ( .A1(csr_n1160), .A2(csr_n_T_444[12]), .A3(csr_n1497), 
        .A4(csr_reg_mtvec_12_), .Y(csr_n86) );
  AO22X1_LVT csr_U131 ( .A1(csr_n1493), .A2(csr_reg_dpc_12_), .A3(csr_n1472), 
        .A4(io_ptw_pmp_5_addr[12]), .Y(csr_n85) );
  AO22X1_LVT csr_U130 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[12]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[12]), .Y(csr_n84) );
  AO22X1_LVT csr_U129 ( .A1(csr_n1162), .A2(csr_io_time[12]), .A3(csr_n1479), 
        .A4(io_ptw_pmp_7_addr[12]), .Y(csr_n83) );
  AO22X1_LVT csr_U128 ( .A1(csr_n1489), .A2(csr_reg_mepc_12_), .A3(csr_n1494), 
        .A4(io_ptw_pmp_6_addr[12]), .Y(csr_n82) );
  AND3X1_LVT csr_U127 ( .A1(csr_io_rw_addr[6]), .A2(csr_io_rw_addr[9]), .A3(
        csr_n1527), .Y(csr_n620) );
  AND3X1_LVT csr_U126 ( .A1(csr_n1405), .A2(ibuf_io_inst_0_bits_raw[25]), .A3(
        csr_n1368), .Y(csr_n1384) );
  OA222X1_LVT csr_U125 ( .A1(n_T_1165[56]), .A2(csr_io_rw_rdata[56]), .A3(
        n_T_1165[56]), .A4(wb_ctrl_csr[1]), .A5(csr_n516), .A6(csr_n81), .Y(
        csr_wdata_56_) );
  INVX0_LVT csr_U124 ( .A(n_T_1165[56]), .Y(csr_n81) );
  NAND3X0_LVT csr_U123 ( .A1(csr_n931), .A2(csr_n590), .A3(csr_n80), .Y(
        csr_N333) );
  AOI22X1_LVT csr_U122 ( .A1(csr_n_1930_), .A2(csr_n930), .A3(
        io_ptw_status_prv[0]), .A4(csr_n929), .Y(csr_n80) );
  AO22X1_LVT csr_U121 ( .A1(csr_n1149), .A2(csr_wdata_3_), .A3(csr_n79), .A4(
        csr_n1446), .Y(csr_N1825) );
  HADDX1_LVT csr_U120 ( .A0(csr_n1144), .B0(csr_io_time[3]), .SO(csr_n79) );
  NAND4X0_LVT csr_U119 ( .A1(csr_n64), .A2(csr_n65), .A3(csr_n66), .A4(csr_n78), .Y(csr_io_rw_rdata[14]) );
  NOR4X0_LVT csr_U118 ( .A1(csr_n67), .A2(csr_n68), .A3(csr_n69), .A4(csr_n77), 
        .Y(csr_n78) );
  AO22X1_LVT csr_U117 ( .A1(csr_n1506), .A2(csr_reg_sepc_14_), .A3(csr_n1472), 
        .A4(io_ptw_pmp_5_addr[14]), .Y(csr_n76) );
  AO21X1_LVT csr_U116 ( .A1(csr_n1510), .A2(csr_reg_dscratch[14]), .A3(csr_n74), .Y(csr_n75) );
  AO22X1_LVT csr_U114 ( .A1(csr_n1153), .A2(csr_n_T_383[14]), .A3(csr_n1488), 
        .A4(io_ptw_ptbr_ppn[14]), .Y(csr_n72) );
  AO21X1_LVT csr_U113 ( .A1(csr_n1487), .A2(csr_reg_stvec_14_), .A3(csr_n70), 
        .Y(csr_n71) );
  AO21X1_LVT csr_U112 ( .A1(io_ptw_pmp_4_addr[14]), .A2(csr_n1491), .A3(
        csr_n1156), .Y(csr_n70) );
  AO222X1_LVT csr_U111 ( .A1(csr_n1162), .A2(csr_io_time[14]), .A3(csr_n1492), 
        .A4(io_ptw_pmp_2_addr[14]), .A5(csr_n1489), .A6(csr_reg_mepc_14_), .Y(
        csr_n69) );
  AO22X1_LVT csr_U110 ( .A1(csr_n1496), .A2(io_ptw_pmp_1_addr[14]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[14]), .Y(csr_n68) );
  AO22X1_LVT csr_U109 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[14]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[14]), .Y(csr_n67) );
  AOI22X1_LVT csr_U108 ( .A1(csr_n1508), .A2(csr_reg_sscratch[14]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_14_), .Y(csr_n66) );
  AOI22X1_LVT csr_U107 ( .A1(csr_n1485), .A2(csr_reg_mscratch[14]), .A3(
        csr_n1493), .A4(csr_reg_dpc_14_), .Y(csr_n65) );
  AOI22X1_LVT csr_U106 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[14]), .A3(
        csr_n1494), .A4(io_ptw_pmp_6_addr[14]), .Y(csr_n64) );
  OA222X1_LVT csr_U105 ( .A1(n_T_1165[57]), .A2(csr_io_rw_rdata[57]), .A3(
        n_T_1165[57]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n63), .Y(
        csr_wdata_57_) );
  INVX0_LVT csr_U104 ( .A(n_T_1165[57]), .Y(csr_n63) );
  AO22X1_LVT csr_U103 ( .A1(csr_n492), .A2(csr_wdata_4_), .A3(csr_n61), .A4(
        csr_n62), .Y(csr_N1432) );
  INVX0_LVT csr_U102 ( .A(csr_n1459), .Y(csr_n62) );
  OA21X1_LVT csr_U101 ( .A1(csr_n960), .A2(csr_n_T_45_4_), .A3(csr_n961), .Y(
        csr_n61) );
  AO221X1_LVT csr_U100 ( .A1(csr_n951), .A2(csr_io_rw_addr[9]), .A3(csr_n951), 
        .A4(csr_n1931), .A5(csr_n60), .Y(csr_n2157) );
  OR3X1_LVT csr_U99 ( .A1(csr_n952), .A2(csr_n950), .A3(csr_n376), .Y(csr_n60)
         );
  NAND4X0_LVT csr_U98 ( .A1(csr_n52), .A2(csr_n53), .A3(csr_n54), .A4(csr_n59), 
        .Y(csr_io_rw_rdata[13]) );
  NOR4X0_LVT csr_U97 ( .A1(csr_n55), .A2(csr_n56), .A3(csr_n57), .A4(csr_n58), 
        .Y(csr_n59) );
  AO22X1_LVT csr_U96 ( .A1(csr_n1508), .A2(csr_reg_sscratch[13]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[13]), .Y(csr_n58) );
  AO22X1_LVT csr_U95 ( .A1(csr_n1160), .A2(csr_n_T_444[13]), .A3(csr_n1153), 
        .A4(csr_n_T_383[13]), .Y(csr_n57) );
  AO22X1_LVT csr_U94 ( .A1(csr_n1162), .A2(csr_io_time[13]), .A3(csr_n1491), 
        .A4(io_ptw_pmp_4_addr[13]), .Y(csr_n56) );
  AO22X1_LVT csr_U93 ( .A1(csr_n1485), .A2(csr_reg_mscratch[13]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_13_), .Y(csr_n55) );
  AOI22X1_LVT csr_U92 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[13]), .A3(
        csr_n1469), .A4(csr_read_medeleg_13), .Y(csr_n54) );
  AOI22X1_LVT csr_U91 ( .A1(csr_n1489), .A2(csr_reg_mepc_13_), .A3(csr_n1494), 
        .A4(io_ptw_pmp_6_addr[13]), .Y(csr_n53) );
  NOR4X0_LVT csr_U90 ( .A1(csr_n45), .A2(csr_n48), .A3(csr_n49), .A4(csr_n50), 
        .Y(csr_n52) );
  AO22X1_LVT csr_U89 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[13]), .A3(
        csr_n1488), .A4(io_ptw_ptbr_ppn[13]), .Y(csr_n50) );
  AO22X1_LVT csr_U88 ( .A1(csr_n1479), .A2(io_ptw_pmp_7_addr[13]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[13]), .Y(csr_n49) );
  NAND4X0_LVT csr_U87 ( .A1(csr_n1155), .A2(csr_n46), .A3(csr_n758), .A4(
        csr_n47), .Y(csr_n48) );
  AOI22X1_LVT csr_U86 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[13]), .A3(
        csr_n1495), .A4(csr_n_T_1155_1_), .Y(csr_n47) );
  AOI21X1_LVT csr_U85 ( .A1(csr_n_T_45_13_), .A2(csr_n1689), .A3(csr_n1559), 
        .Y(csr_n46) );
  AO22X1_LVT csr_U84 ( .A1(csr_n1487), .A2(csr_reg_stvec_13_), .A3(csr_n1496), 
        .A4(io_ptw_pmp_1_addr[13]), .Y(csr_n45) );
  OR3X1_LVT csr_U83 ( .A1(csr_n31), .A2(csr_n35), .A3(csr_n44), .Y(
        csr_io_rw_rdata[22]) );
  OR4X1_LVT csr_U82 ( .A1(csr_n40), .A2(csr_n41), .A3(csr_n42), .A4(csr_n43), 
        .Y(csr_n44) );
  AO22X1_LVT csr_U81 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[22]), .A3(
        csr_n1480), .A4(io_ptw_pmp_0_addr[22]), .Y(csr_n43) );
  AO22X1_LVT csr_U80 ( .A1(csr_n1510), .A2(csr_reg_dscratch[22]), .A3(
        csr_n1506), .A4(csr_reg_sepc_22_), .Y(csr_n42) );
  AO22X1_LVT csr_U79 ( .A1(csr_n1490), .A2(csr_io_bp_0_address[22]), .A3(
        csr_n1497), .A4(csr_reg_mtvec_22_), .Y(csr_n41) );
  AO22X1_LVT csr_U78 ( .A1(csr_n1485), .A2(csr_reg_mscratch[22]), .A3(
        csr_n1492), .A4(io_ptw_pmp_2_addr[22]), .Y(csr_n38) );
  AO22X1_LVT csr_U77 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[22]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[22]), .Y(csr_n37) );
  AO222X1_LVT csr_U76 ( .A1(csr_n1689), .A2(csr_n_T_45_22_), .A3(csr_n1487), 
        .A4(csr_reg_stvec_22_), .A5(csr_n1493), .A6(csr_reg_dpc_22_), .Y(
        csr_n36) );
  AO22X1_LVT csr_U74 ( .A1(csr_n1162), .A2(csr_io_time[22]), .A3(csr_n1491), 
        .A4(io_ptw_pmp_4_addr[22]), .Y(csr_n33) );
  AO22X1_LVT csr_U73 ( .A1(csr_n1508), .A2(csr_reg_sscratch[22]), .A3(
        csr_n1473), .A4(io_ptw_pmp_3_addr[22]), .Y(csr_n32) );
  AO22X1_LVT csr_U72 ( .A1(csr_n1489), .A2(csr_reg_mepc_22_), .A3(csr_n1496), 
        .A4(io_ptw_pmp_1_addr[22]), .Y(csr_n31) );
  AND2X1_LVT csr_U71 ( .A1(csr_n1194), .A2(csr_n1186), .Y(
        csr_io_interrupt_cause[0]) );
  OA222X1_LVT csr_U70 ( .A1(n_T_1165[58]), .A2(csr_io_rw_rdata[58]), .A3(
        n_T_1165[58]), .A4(csr_n589), .A5(csr_n516), .A6(csr_n30), .Y(
        csr_wdata_58_) );
  INVX0_LVT csr_U69 ( .A(n_T_1165[58]), .Y(csr_n30) );
  AO21X1_LVT csr_U68 ( .A1(csr_reg_mepc_34_), .A2(csr_n502), .A3(csr_n29), .Y(
        csr_io_evec[34]) );
  AO222X1_LVT csr_U67 ( .A1(csr_reg_sepc_34_), .A2(csr_n500), .A3(
        csr_reg_dpc_34_), .A4(csr_n1356), .A5(csr_reg_stvec_34_), .A6(csr_n499), .Y(csr_n29) );
  NAND3X0_LVT csr_U66 ( .A1(csr_n1472), .A2(csr_n437), .A3(csr_n28), .Y(
        csr_n434) );
  NAND3X0_LVT csr_U65 ( .A1(io_ptw_pmp_6_cfg_l), .A2(csr_n458), .A3(
        io_ptw_pmp_6_cfg_a[0]), .Y(csr_n28) );
  OR2X1_LVT csr_U64 ( .A1(csr_n1375), .A2(csr_n27), .Y(csr_n1396) );
  NAND4X0_LVT csr_U63 ( .A1(csr_n1390), .A2(csr_n1379), .A3(csr_n1417), .A4(
        ibuf_io_inst_0_bits_raw[27]), .Y(csr_n27) );
  AO22X1_LVT csr_U62 ( .A1(csr_n1129), .A2(csr_n_T_44[52]), .A3(csr_wdata_58_), 
        .A4(csr_n1128), .Y(csr_N1549) );
  INVX0_LVT csr_U60 ( .A(csr_n1357), .Y(csr_n25) );
  AO22X1_LVT csr_U59 ( .A1(csr_reg_sepc_39_), .A2(csr_n1355), .A3(csr_n1356), 
        .A4(csr_reg_dpc_39_), .Y(csr_n24) );
  NAND2X0_LVT csr_U58 ( .A1(csr_n13), .A2(csr_n23), .Y(csr_io_rw_rdata[6]) );
  NOR4X0_LVT csr_U57 ( .A1(csr_n17), .A2(csr_n18), .A3(csr_n19), .A4(csr_n22), 
        .Y(csr_n23) );
  AO22X1_LVT csr_U56 ( .A1(csr_n1472), .A2(io_ptw_pmp_5_addr[6]), .A3(
        csr_n1477), .A4(io_fpu_fcsr_rm[1]), .Y(csr_n21) );
  AO22X1_LVT csr_U55 ( .A1(csr_n1489), .A2(csr_reg_mepc_6_), .A3(csr_n1490), 
        .A4(csr_io_bp_0_address[6]), .Y(csr_n20) );
  AO22X1_LVT csr_U54 ( .A1(csr_n1485), .A2(csr_reg_mscratch[6]), .A3(csr_n1473), .A4(io_ptw_pmp_3_addr[6]), .Y(csr_n19) );
  AO22X1_LVT csr_U53 ( .A1(csr_n1492), .A2(io_ptw_pmp_2_addr[6]), .A3(
        csr_n1469), .A4(csr_read_medeleg_6), .Y(csr_n18) );
  AO22X1_LVT csr_U51 ( .A1(csr_n1494), .A2(io_ptw_pmp_6_addr[6]), .A3(
        csr_n1470), .A4(csr_reg_mtvec_6_), .Y(csr_n15) );
  AO22X1_LVT csr_U50 ( .A1(csr_n1162), .A2(csr_io_time[6]), .A3(csr_n1496), 
        .A4(io_ptw_pmp_1_addr[6]), .Y(csr_n14) );
  NOR4X0_LVT csr_U49 ( .A1(csr_n9), .A2(csr_n10), .A3(csr_n11), .A4(csr_n12), 
        .Y(csr_n13) );
  AO22X1_LVT csr_U48 ( .A1(csr_n1480), .A2(io_ptw_pmp_0_addr[6]), .A3(
        csr_n1479), .A4(io_ptw_pmp_7_addr[6]), .Y(csr_n12) );
  AO22X1_LVT csr_U47 ( .A1(csr_n1508), .A2(csr_reg_sscratch[6]), .A3(csr_n1160), .A4(csr_n_T_444[6]), .Y(csr_n11) );
  AO22X1_LVT csr_U46 ( .A1(csr_n1506), .A2(csr_reg_sepc_6_), .A3(csr_n1478), 
        .A4(csr_reg_stvec_6_), .Y(csr_n10) );
  NAND4X0_LVT csr_U45 ( .A1(csr_n6), .A2(csr_n7), .A3(csr_n924), .A4(csr_n8), 
        .Y(csr_n9) );
  NAND2X0_LVT csr_U44 ( .A1(csr_n1481), .A2(csr_io_bp_0_control_m), .Y(csr_n8)
         );
  AOI22X1_LVT csr_U43 ( .A1(csr_n1510), .A2(csr_reg_dscratch[6]), .A3(
        csr_n1689), .A4(csr_n_T_45_6_), .Y(csr_n7) );
  AOI22X1_LVT csr_U42 ( .A1(csr_n1495), .A2(csr_n_T_389[6]), .A3(csr_n1488), 
        .A4(io_ptw_ptbr_ppn[6]), .Y(csr_n6) );
  AO22X1_LVT csr_U41 ( .A1(csr_n492), .A2(csr_wdata_5_), .A3(csr_n5), .A4(
        csr_n961), .Y(csr_N1433) );
  HADDX1_LVT csr_U40 ( .A0(csr_n1459), .B0(csr_n_T_45_5_), .SO(csr_n5) );
  AO22X1_LVT csr_U38 ( .A1(csr_reg_mepc_30_), .A2(csr_n502), .A3(
        csr_reg_mtvec_30_), .A4(csr_n1333), .Y(csr_n3) );
  AO22X1_LVT csr_U37 ( .A1(csr_reg_sepc_30_), .A2(csr_n500), .A3(
        csr_reg_dpc_30_), .A4(csr_n1356), .Y(csr_n2) );
  NAND2X0_LVT csr_U36 ( .A1(csr_n1374), .A2(csr_n1), .Y(csr_n1416) );
  NAND3X0_LVT csr_U35 ( .A1(csr_n1384), .A2(csr_n489), .A3(csr_n1386), .Y(
        csr_n1) );
  IBUFFX2_LVT csr_U34 ( .A(csr_n1204), .Y(csr_n1333) );
  AO221X1_LVT csr_U33 ( .A1(1'b1), .A2(csr_n2), .A3(csr_n499), .A4(
        csr_reg_stvec_30_), .A5(csr_n3), .Y(csr_io_evec[30]) );
  AO221X1_LVT csr_U32 ( .A1(1'b1), .A2(csr_n20), .A3(csr_n1491), .A4(
        io_ptw_pmp_4_addr[6]), .A5(csr_n21), .Y(csr_n22) );
  AO221X1_LVT csr_U31 ( .A1(1'b1), .A2(csr_n14), .A3(csr_n1493), .A4(
        csr_reg_dpc_6_), .A5(csr_n15), .Y(csr_n17) );
  AO221X1_LVT csr_U30 ( .A1(1'b1), .A2(csr_n24), .A3(csr_reg_mepc_39_), .A4(
        csr_n502), .A5(csr_n25), .Y(csr_io_evec[39]) );
  AO221X1_LVT csr_U29 ( .A1(1'b1), .A2(csr_n36), .A3(csr_n1153), .A4(
        csr_n_T_383[22]), .A5(csr_n39), .Y(csr_n40) );
  AO221X1_LVT csr_U28 ( .A1(1'b1), .A2(csr_n37), .A3(csr_n1157), .A4(csr_n1924), .A5(csr_n38), .Y(csr_n39) );
  AO221X1_LVT csr_U27 ( .A1(1'b1), .A2(csr_n32), .A3(csr_n1160), .A4(
        csr_n_T_444[22]), .A5(csr_n33), .Y(csr_n35) );
  AO221X1_LVT csr_U26 ( .A1(1'b1), .A2(csr_n75), .A3(csr_n1160), .A4(
        csr_n_T_444[14]), .A5(csr_n76), .Y(csr_n77) );
  AO221X1_LVT csr_U25 ( .A1(1'b1), .A2(csr_n71), .A3(csr_n1689), .A4(
        csr_n_T_45_14_), .A5(csr_n72), .Y(csr_n74) );
  AO221X1_LVT csr_U24 ( .A1(1'b1), .A2(csr_n91), .A3(csr_n1153), .A4(
        csr_n_T_383[12]), .A5(csr_n95), .Y(csr_n96) );
  AO221X1_LVT csr_U23 ( .A1(1'b1), .A2(csr_n93), .A3(csr_n1496), .A4(
        io_ptw_pmp_1_addr[12]), .A5(csr_n94), .Y(csr_n95) );
  AO221X1_LVT csr_U22 ( .A1(1'b1), .A2(csr_n669), .A3(io_ptw_pmp_1_cfg_a[1]), 
        .A4(csr_n1507), .A5(csr_n92), .Y(csr_n93) );
  AO221X1_LVT csr_U21 ( .A1(1'b1), .A2(csr_n87), .A3(csr_n1508), .A4(
        csr_reg_sscratch[12]), .A5(csr_n88), .Y(csr_n90) );
  AO221X1_LVT csr_U20 ( .A1(1'b1), .A2(csr_n142), .A3(csr_n1167), .A4(
        csr_read_fcsr_4_), .A5(csr_n143), .Y(csr_n145) );
  AO221X1_LVT csr_U19 ( .A1(1'b1), .A2(csr_n163), .A3(csr_n1153), .A4(
        csr_n_T_383[25]), .A5(csr_n164), .Y(csr_n166) );
  AO221X1_LVT csr_U18 ( .A1(1'b1), .A2(csr_n180), .A3(csr_n1487), .A4(
        csr_reg_stvec_15_), .A5(csr_n181), .Y(csr_n182) );
  AO221X1_LVT csr_U17 ( .A1(1'b1), .A2(csr_n1560), .A3(csr_n_T_45_15_), .A4(
        csr_n1689), .A5(csr_n178), .Y(csr_n180) );
  AO221X1_LVT csr_U16 ( .A1(1'b1), .A2(csr_n191), .A3(csr_n1487), .A4(
        csr_reg_stvec_35_), .A5(csr_n196), .Y(csr_n201) );
  AO221X1_LVT csr_U15 ( .A1(1'b1), .A2(csr_n224), .A3(csr_n1160), .A4(
        csr_n_T_444[33]), .A5(csr_n228), .Y(csr_n230) );
  AO221X1_LVT csr_U14 ( .A1(1'b1), .A2(csr_n241), .A3(csr_n1510), .A4(
        csr_reg_dscratch[26]), .A5(csr_n242), .Y(csr_n244) );
  AO221X1_LVT csr_U13 ( .A1(1'b1), .A2(csr_n258), .A3(csr_n1153), .A4(
        csr_n_T_383[28]), .A5(csr_n259), .Y(csr_n260) );
  AO221X1_LVT csr_U12 ( .A1(1'b1), .A2(csr_n255), .A3(csr_n1507), .A4(
        io_ptw_pmp_3_cfg_a[1]), .A5(csr_n256), .Y(csr_n258) );
  AO221X1_LVT csr_U11 ( .A1(1'b1), .A2(csr_n262), .A3(csr_n1485), .A4(
        csr_reg_mscratch[31]), .A5(csr_n270), .Y(csr_io_rw_rdata[31]) );
  AO221X1_LVT csr_U10 ( .A1(1'b1), .A2(csr_n263), .A3(csr_n1510), .A4(
        csr_reg_dscratch[31]), .A5(csr_n269), .Y(csr_n270) );
  AO221X1_LVT csr_U9 ( .A1(1'b1), .A2(csr_n267), .A3(csr_n1507), .A4(
        io_ptw_pmp_3_cfg_l), .A5(csr_n268), .Y(csr_n269) );
  AO221X1_LVT csr_U8 ( .A1(1'b1), .A2(csr_n264), .A3(csr_n1689), .A4(
        csr_n_T_45_31_), .A5(csr_n265), .Y(csr_n267) );
  AO221X1_LVT csr_U7 ( .A1(1'b1), .A2(csr_n1650), .A3(csr_n1485), .A4(
        csr_reg_mscratch[38]), .A5(csr_n282), .Y(csr_n283) );
  AO221X1_LVT csr_U6 ( .A1(1'b1), .A2(csr_n277), .A3(csr_n1162), .A4(csr_n1961), .A5(csr_n278), .Y(csr_n280) );
  AO221X1_LVT csr_U5 ( .A1(1'b1), .A2(csr_n1533), .A3(csr_n_T_45_8_), .A4(
        csr_n1689), .A5(csr_n286), .Y(csr_n288) );
  AO221X1_LVT csr_U4 ( .A1(1'b1), .A2(csr_n333), .A3(csr_n1153), .A4(
        csr_n_T_383[21]), .A5(csr_n334), .Y(csr_n336) );
  AO222X1_LVT csr_U3 ( .A1(csr_n323), .A2(csr_n1185), .A3(io_interrupts_debug), 
        .A4(1'b1), .A5(csr_n1183), .A6(csr_n1184), .Y(
        csr_io_interrupt_cause[2]) );
  DFFX1_LVT csr_reg_mstatus_mie_reg ( .D(csr_n365), .CLK(csr_net35147), .Q(
        csr_n383), .QN(csr_n1934) );
  OA21X1_LVT csr_reg_mstatus_mie_reg_U2 ( .A1(csr_n1346), .A2(csr_n1041), .A3(
        csr_n194), .Y(csr_n365) );
  DFFX1_LVT csr_reg_dcsr_cause_reg_0_ ( .D(csr_n366), .CLK(csr_net35177), .Q(
        csr_n_T_389[6]) );
  DFFX1_LVT csr_reg_dscratch_reg_2_ ( .D(csr_n1483), .CLK(csr_n527), .QN(
        csr_reg_dscratch[2]) );
  DFFX1_LVT csr_reg_dscratch_reg_12_ ( .D(csr_n367), .CLK(csr_n527), .QN(
        csr_reg_dscratch[12]) );
  DFFX1_LVT csr_reg_mscratch_reg_2_ ( .D(csr_n1483), .CLK(csr_n553), .QN(
        csr_reg_mscratch[2]) );
  DFFX1_LVT csr_reg_mscratch_reg_12_ ( .D(csr_n367), .CLK(csr_n553), .QN(
        csr_reg_mscratch[12]) );
  DFFX1_LVT csr_reg_sscratch_reg_2_ ( .D(csr_n1483), .CLK(csr_n567), .QN(
        csr_reg_sscratch[2]) );
  DFFX1_LVT csr_reg_sscratch_reg_12_ ( .D(csr_n367), .CLK(csr_n567), .QN(
        csr_reg_sscratch[12]) );
  DFFX1_LVT csr_reg_medeleg_reg_2_ ( .D(csr_n1483), .CLK(csr_net35172), .QN(
        csr_read_medeleg_2_) );
  DFFX1_LVT csr_reg_medeleg_reg_12_ ( .D(csr_n367), .CLK(csr_net35172), .QN(
        csr_read_medeleg_12) );
  DFFX1_LVT csr_reg_mcounteren_reg_2_ ( .D(csr_n1483), .CLK(csr_net34945), 
        .QN(csr_read_mcounteren_2_) );
  DFFX1_LVT csr_reg_scounteren_reg_2_ ( .D(csr_n1483), .CLK(csr_net34940), 
        .QN(csr_read_scounteren_2_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_2_ ( .D(csr_n1483), .CLK(csr_n586), .QN(
        csr_io_bp_0_address[2]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_12_ ( .D(csr_n367), .CLK(csr_n586), .QN(
        csr_io_bp_0_address[12]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_14_ ( .D(csr_n51), .CLK(csr_n586), .QN(
        csr_io_bp_0_address[14]) );
  DFFX1_LVT csr_reg_pmp_0_cfg_x_reg ( .D(csr_n1483), .CLK(csr_net34733), .QN(
        io_ptw_pmp_0_cfg_x) );
  DFFX1_LVT csr_reg_misa_reg_12_ ( .D(csr_n368), .CLK(csr_net35137), .Q(
        csr_io_status_isa[12]), .QN(csr_io_status_isa_12_) );
  OA21X1_LVT csr_reg_misa_reg_12__U2 ( .A1(csr_n367), .A2(csr_n387), .A3(
        csr_n590), .Y(csr_n368) );
  INVX0_LVT csr_reg_misa_reg_12__U4 ( .A(csr_wdata_12_), .Y(csr_n367) );
  DFFX1_LVT csr_reg_pmp_6_cfg_w_reg ( .D(csr_n369), .CLK(csr_net35107), .Q(
        io_ptw_pmp_6_cfg_w) );
  DFFX1_LVT csr_reg_mtvec_reg_31_ ( .D(csr_n370), .CLK(csr_net34950), .QN(
        csr_reg_mtvec_31_) );
  DFFX1_LVT csr_reg_mtvec_reg_0_ ( .D(csr_n371), .CLK(csr_net34950), .Q(
        csr_n416), .QN(csr_n659) );
  DFFX1_LVT csr_u_T_41_reg_48_ ( .D(csr_N1545), .CLK(csr_net34890), .Q(
        csr_n_T_45_54_) );
  DFFX1_LVT csr_reg_dcsr_cause_reg_2_ ( .D(csr_n373), .CLK(csr_net35177), .QN(
        csr_n_T_389[8]) );
  INVX0_LVT csr_reg_dcsr_cause_reg_2__U4 ( .A(csr_n1499), .Y(csr_n372) );
  DFFX1_LVT csr_reg_pmp_6_cfg_l_reg ( .D(csr_n374), .CLK(csr_net35102), .Q(
        io_ptw_pmp_6_cfg_l), .QN(csr_n439) );
  DFFX1_LVT csr_reg_mstatus_prv_reg_1_ ( .D(csr_n2160), .CLK(csr_n594), .Q(
        io_ptw_status_prv[1]), .QN(csr_n381) );
  DFFX1_LVT csr_reg_mstatus_prv_reg_0_ ( .D(csr_n2157), .CLK(csr_n594), .Q(
        io_ptw_status_prv[0]), .QN(csr_n429) );
  DFFX1_LVT csr_reg_custom_0_reg_3_ ( .D(csr_n1909), .CLK(csr_n594), .Q(
        csr_n1910), .QN(io_ptw_customCSRs_csrs_0_value[3]) );
  DFFX1_LVT csr_reg_custom_0_reg_9_ ( .D(csr_n1911), .CLK(csr_n594), .Q(
        csr_n1912), .QN(io_ptw_customCSRs_csrs_0_value[9]) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_0_5 csr_clk_gate_reg_mstatus_spie_reg ( .CLK(
        csr_n593), .EN(csr_n1917), .ENCLK(csr_n1915), .TE(1'b0) );
  DFFX1_LVT csr_u_T_1196_reg_1_ ( .D(csr_N1692), .CLK(csr_n593), .Q(
        io_dmem_req_bits_dprv[1]) );
  DFFX1_LVT csr_reg_dpc_reg_12_ ( .D(csr_net35268), .CLK(csr_net35304), .Q(
        csr_reg_dpc_12_) );
  DFFX1_LVT csr_reg_mepc_reg_12_ ( .D(csr_net35046), .CLK(csr_net35082), .Q(
        csr_reg_mepc_12_) );
  DFFX1_LVT csr_reg_sepc_reg_12_ ( .D(csr_net34844), .CLK(csr_net34880), .Q(
        csr_reg_sepc_12_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_12_ ( .D(csr_n_GEN_307[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_7_addr[12]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_12_ ( .D(csr_n_GEN_300[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_6_addr[12]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_12_ ( .D(csr_n_GEN_293[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_5_addr[12]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_12_ ( .D(csr_n_GEN_286[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_4_addr[12]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_12_ ( .D(csr_n_GEN_279[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_3_addr[12]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_12_ ( .D(csr_n_GEN_272[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_2_addr[12]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_12_ ( .D(csr_n_GEN_265[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_1_addr[12]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_12_ ( .D(csr_n_GEN_258[12]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_0_addr[12]) );
  DFFX1_LVT csr_reg_dpc_reg_9_ ( .D(csr_net35277), .CLK(csr_net35304), .Q(
        csr_reg_dpc_9_) );
  DFFX1_LVT csr_reg_mepc_reg_9_ ( .D(csr_net35055), .CLK(csr_net35082), .Q(
        csr_reg_mepc_9_) );
  DFFX1_LVT csr_reg_sepc_reg_9_ ( .D(csr_net34853), .CLK(csr_net34880), .Q(
        csr_reg_sepc_9_) );
  DFFSSRX1_LVT csr_reg_pmp_1_cfg_w_reg ( .D(csr_wdata_8_), .SETB(1'b1), .RSTB(
        csr_wdata_9_), .CLK(csr_net35087), .Q(io_ptw_pmp_1_cfg_w) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_9_ ( .D(csr_n_GEN_307[9]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_7_addr[9]), .QN(csr_n424) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_9_ ( .D(csr_n_GEN_300[9]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_6_addr[9]), .QN(csr_n420) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_9_ ( .D(csr_n_GEN_293[9]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_5_addr[9]), .QN(csr_n422) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_9_ ( .D(csr_n_GEN_286[9]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_4_addr[9]), .QN(csr_n423) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_9_ ( .D(csr_n_GEN_279[9]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_3_addr[9]), .QN(csr_n418) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_9_ ( .D(csr_n_GEN_272[9]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_2_addr[9]), .QN(csr_n421) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_9_ ( .D(csr_n_GEN_265[9]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_1_addr[9]), .QN(csr_n425) );
  DFFX1_LVT csr_reg_wfi_reg ( .D(csr_N1821), .CLK(csr_n591), .Q(io_wfi), .QN(
        csr_n472) );
  DFFX1_LVT csr_reg_mie_reg_9_ ( .D(csr_N615), .CLK(csr_net34728), .Q(
        csr_reg_mie_9_) );
  DFFX1_LVT csr_u_T_49_reg_3_ ( .D(csr_N1894), .CLK(csr_n517), .Q(
        csr_io_time[9]) );
  DFFX1_LVT csr_u_T_41_reg_3_ ( .D(csr_N1500), .CLK(csr_n575), .Q(
        csr_n_T_45_9_) );
  DFFX1_LVT csr_reg_stval_reg_9_ ( .D(csr_N1391), .CLK(csr_net34930), .Q(
        csr_n_T_444[9]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_9_ ( .D(csr_n376), .SETB(csr_wdata_9_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_9_) );
  DFFX1_LVT csr_reg_mtval_reg_9_ ( .D(csr_N1002), .CLK(csr_net34895), .Q(
        csr_n_T_383[9]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[9]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_n587), 
        .Q(csr_io_bp_0_address[9]) );
  DFFX1_LVT csr_reg_sscratch_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[9]) );
  DFFX1_LVT csr_reg_mscratch_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[9]) );
  DFFX1_LVT csr_reg_dscratch_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[9]) );
  DFFX1_LVT csr_reg_dpc_reg_7_ ( .D(csr_net35283), .CLK(csr_net35304), .Q(
        csr_reg_dpc_7_) );
  DFFX1_LVT csr_reg_mepc_reg_7_ ( .D(csr_net35061), .CLK(csr_net35082), .Q(
        csr_reg_mepc_7_) );
  DFFX1_LVT csr_reg_sepc_reg_7_ ( .D(csr_net34859), .CLK(csr_net34880), .Q(
        csr_reg_sepc_7_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_7_ ( .D(csr_n_GEN_307[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_7_addr[7]), .QN(csr_n394) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_7_ ( .D(csr_n_GEN_300[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_6_addr[7]), .QN(csr_n391) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_7_ ( .D(csr_n_GEN_293[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_5_addr[7]), .QN(csr_n392) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_7_ ( .D(csr_n_GEN_286[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_4_addr[7]), .QN(csr_n395) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_7_ ( .D(csr_n_GEN_279[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_3_addr[7]), .QN(csr_n396) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_7_ ( .D(csr_n_GEN_272[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_2_addr[7]), .QN(csr_n393) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_7_ ( .D(csr_n_GEN_265[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_1_addr[7]), .QN(csr_n397) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_7_ ( .D(csr_n_GEN_258[7]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_0_addr[7]), .QN(csr_n398) );
  DFFSSRX1_LVT csr_reg_misa_reg_0_ ( .D(csr_n387), .SETB(csr_wdata_0_), .RSTB(
        csr_n590), .CLK(csr_net35137), .Q(csr_io_status_isa[0]), .QN(
        csr_io_status_isa_0_) );
  DFFX1_LVT csr_reg_mip_ssip_reg ( .D(csr_n2162), .CLK(csr_n533), .Q(
        csr_n_T_61_1) );
  DFFX1_LVT csr_reg_dpc_reg_1_ ( .D(csr_net35301), .CLK(csr_n530), .Q(
        csr_reg_dpc_1_) );
  DFFX1_LVT csr_reg_mepc_reg_1_ ( .D(csr_net35079), .CLK(csr_n547), .Q(
        csr_reg_mepc_1_) );
  DFFX1_LVT csr_reg_sepc_reg_1_ ( .D(csr_net34877), .CLK(csr_n583), .Q(
        csr_reg_sepc_1_) );
  DFFX1_LVT csr_reg_dcsr_prv_reg_1_ ( .D(csr_n2155), .CLK(csr_n593), .Q(
        csr_n_T_389_1) );
  DFFSSRX1_LVT csr_reg_pmp_0_cfg_w_reg ( .D(csr_wdata_1_), .SETB(1'b1), .RSTB(
        csr_wdata_0_), .CLK(csr_net34733), .Q(io_ptw_pmp_0_cfg_w) );
  DFFX1_LVT csr_reg_fflags_reg_1_ ( .D(csr_n_GEN_345[1]), .CLK(csr_n594), .Q(
        csr_read_fcsr_1_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_1_ ( .D(csr_n_GEN_307[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_7_addr[1]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_1_ ( .D(csr_n_GEN_300[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_6_addr[1]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_1_ ( .D(csr_n_GEN_293[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_5_addr[1]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_1_ ( .D(csr_n_GEN_286[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_4_addr[1]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_1_ ( .D(csr_n_GEN_279[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_3_addr[1]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_1_ ( .D(csr_n_GEN_272[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_2_addr[1]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_1_ ( .D(csr_n_GEN_265[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_1_addr[1]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_1_ ( .D(csr_n_GEN_258[1]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_0_addr[1]) );
  DFFX1_LVT csr_reg_dpc_reg_6_ ( .D(csr_net35286), .CLK(csr_n530), .Q(
        csr_reg_dpc_6_) );
  DFFX1_LVT csr_reg_mepc_reg_6_ ( .D(csr_net35064), .CLK(csr_n547), .Q(
        csr_reg_mepc_6_) );
  DFFX1_LVT csr_reg_sepc_reg_6_ ( .D(csr_net34862), .CLK(csr_n583), .Q(
        csr_reg_sepc_6_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_6_ ( .D(csr_n_GEN_307[6]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_7_addr[6]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_6_ ( .D(csr_n_GEN_300[6]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_6_addr[6]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_6_ ( .D(csr_n_GEN_293[6]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_5_addr[6]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_6_ ( .D(csr_n_GEN_286[6]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_4_addr[6]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_6_ ( .D(csr_n_GEN_279[6]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_3_addr[6]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_6_ ( .D(csr_n_GEN_272[6]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_2_addr[6]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_6_ ( .D(csr_n_GEN_265[6]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_1_addr[6]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_6_ ( .D(csr_n_GEN_258[6]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_0_addr[6]) );
  DFFX1_LVT csr_reg_mtval_reg_6_ ( .D(csr_N999), .CLK(csr_net34895), .Q(
        csr_n_T_383[6]) );
  DFFX1_LVT csr_u_T_49_reg_0_ ( .D(csr_N1891), .CLK(csr_n517), .Q(
        csr_io_time[6]), .QN(csr_n456) );
  DFFX1_LVT csr_u_T_41_reg_0_ ( .D(csr_N1497), .CLK(csr_n575), .Q(
        csr_n_T_45_6_), .QN(csr_n455) );
  DFFX1_LVT csr_reg_stval_reg_6_ ( .D(csr_N1388), .CLK(csr_net34930), .Q(
        csr_n_T_444[6]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_6_ ( .D(csr_n378), .SETB(csr_wdata_6_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_6_) );
  DFFX1_LVT csr_reg_satp_ppn_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[6]) );
  DFFX1_LVT csr_reg_bp_0_control_m_reg ( .D(csr_wdata_6_), .CLK(csr_net35319), 
        .Q(csr_io_bp_0_control_m) );
  DFFX1_LVT csr_reg_bp_0_address_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_n587), 
        .Q(csr_io_bp_0_address[6]) );
  DFFX1_LVT csr_reg_sscratch_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[6]) );
  DFFX1_LVT csr_reg_mscratch_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[6]) );
  DFFX1_LVT csr_reg_dscratch_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[6]) );
  DFFX1_LVT csr_reg_medeleg_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_net35172), .Q(
        csr_read_medeleg_6) );
  DFFX1_LVT csr_reg_stvec_reg_6_ ( .D(csr_wdata_6_), .CLK(csr_n571), .Q(
        csr_reg_stvec_6_) );
  DFFX1_LVT csr_reg_frm_reg_1_ ( .D(csr_n_GEN_155[1]), .CLK(csr_net34900), .Q(
        io_fpu_fcsr_rm[1]) );
  DFFX1_LVT csr_reg_mtval_reg_1_ ( .D(csr_N994), .CLK(csr_net34895), .Q(
        csr_n_T_383[1]) );
  DFFX1_LVT csr_reg_mie_reg_1_ ( .D(csr_N607), .CLK(csr_net34728), .Q(
        csr_reg_mie_1_) );
  DFFX1_LVT csr_reg_dpc_reg_5_ ( .D(csr_net35289), .CLK(csr_n530), .Q(
        csr_reg_dpc_5_) );
  DFFX1_LVT csr_reg_mepc_reg_5_ ( .D(csr_net35067), .CLK(csr_n547), .Q(
        csr_reg_mepc_5_) );
  DFFX1_LVT csr_reg_sepc_reg_5_ ( .D(csr_net34865), .CLK(csr_n583), .Q(
        csr_reg_sepc_5_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_5_ ( .D(csr_n_GEN_307[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_7_addr[5]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_5_ ( .D(csr_n_GEN_300[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_6_addr[5]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_5_ ( .D(csr_n_GEN_293[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_5_addr[5]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_5_ ( .D(csr_n_GEN_286[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_4_addr[5]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_5_ ( .D(csr_n_GEN_279[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_3_addr[5]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_5_ ( .D(csr_n_GEN_272[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_2_addr[5]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_5_ ( .D(csr_n_GEN_265[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_1_addr[5]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_5_ ( .D(csr_n_GEN_258[5]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_0_addr[5]) );
  DFFX1_LVT csr_reg_frm_reg_0_ ( .D(csr_n_GEN_155[0]), .CLK(csr_net34900), .Q(
        io_fpu_fcsr_rm[0]) );
  DFFX1_LVT csr_reg_mtval_reg_5_ ( .D(csr_N998), .CLK(csr_net34895), .Q(
        csr_n_T_383[5]) );
  DFFX1_LVT csr_reg_mie_reg_5_ ( .D(csr_N611), .CLK(csr_net34728), .Q(
        csr_reg_mie_5_) );
  DFFX1_LVT csr_u_T_47_reg_5_ ( .D(csr_N1827), .CLK(csr_n591), .Q(
        csr_io_time[5]) );
  DFFSSRX1_LVT csr_reg_misa_reg_5_ ( .D(csr_n387), .SETB(csr_wdata_5_), .RSTB(
        csr_n590), .CLK(csr_net35137), .QN(csr_n1923) );
  DFFX1_LVT csr_reg_dpc_reg_3_ ( .D(csr_net35295), .CLK(csr_n530), .Q(
        csr_reg_dpc_3_) );
  DFFX1_LVT csr_reg_mepc_reg_3_ ( .D(csr_net35073), .CLK(csr_n547), .Q(
        csr_reg_mepc_3_) );
  DFFX1_LVT csr_reg_sepc_reg_3_ ( .D(csr_net34871), .CLK(csr_n583), .Q(
        csr_reg_sepc_3_) );
  DFFX1_LVT csr_reg_fflags_reg_3_ ( .D(csr_n_GEN_345[3]), .CLK(csr_n593), .Q(
        csr_read_fcsr_3_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_3_ ( .D(csr_n_GEN_307[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_7_addr[3]), .QN(csr_n412) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_3_ ( .D(csr_n_GEN_300[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_6_addr[3]), .QN(csr_n413) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_3_ ( .D(csr_n_GEN_293[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_5_addr[3]), .QN(csr_n414) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_3_ ( .D(csr_n_GEN_286[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_4_addr[3]), .QN(csr_n408) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_3_ ( .D(csr_n_GEN_279[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_3_addr[3]), .QN(csr_n409) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_3_ ( .D(csr_n_GEN_272[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_2_addr[3]), .QN(csr_n410) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_3_ ( .D(csr_n_GEN_265[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_1_addr[3]), .QN(csr_n411) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_3_ ( .D(csr_n_GEN_258[3]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_0_addr[3]), .QN(csr_n415) );
  DFFX1_LVT csr_reg_mtval_reg_3_ ( .D(csr_N996), .CLK(csr_n574), .Q(
        csr_n_T_383[3]) );
  DFFX1_LVT csr_reg_mie_reg_3_ ( .D(csr_N609), .CLK(csr_net34728), .Q(
        csr_reg_mie_3_) );
  DFFSSRX1_LVT csr_reg_pmp_0_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_3_), .CLK(csr_net34905), .Q(io_ptw_pmp_0_cfg_a[0]) );
  DFFX1_LVT csr_u_T_39_reg_3_ ( .D(csr_N1431), .CLK(csr_n593), .Q(
        csr_n_T_45_3_) );
  DFFX1_LVT csr_u_T_47_reg_3_ ( .D(csr_N1825), .CLK(csr_n591), .Q(
        csr_io_time[3]) );
  DFFX1_LVT csr_reg_mcause_reg_3_ ( .D(csr_N884), .CLK(csr_n580), .Q(
        csr_reg_mcause[3]) );
  DFFX1_LVT csr_reg_stval_reg_3_ ( .D(csr_N1385), .CLK(csr_net34930), .Q(
        csr_n_T_444[3]) );
  DFFX1_LVT csr_reg_scause_reg_3_ ( .D(csr_N1273), .CLK(csr_n558), .Q(
        csr_reg_scause[3]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_3_ ( .D(csr_n378), .SETB(csr_wdata_3_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_3_) );
  DFFX1_LVT csr_reg_satp_ppn_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[3]) );
  DFFX1_LVT csr_reg_bp_0_control_u_reg ( .D(csr_wdata_3_), .CLK(csr_net35319), 
        .Q(csr_io_bp_0_control_u) );
  DFFX1_LVT csr_reg_bp_0_address_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_n587), 
        .Q(csr_io_bp_0_address[3]) );
  DFFX1_LVT csr_reg_sscratch_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[3]) );
  DFFX1_LVT csr_reg_mscratch_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[3]) );
  DFFX1_LVT csr_reg_dscratch_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[3]) );
  DFFX1_LVT csr_reg_medeleg_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_net35172), .Q(
        csr_read_medeleg_3_) );
  DFFX1_LVT csr_reg_stvec_reg_3_ ( .D(csr_wdata_3_), .CLK(csr_n571), .Q(
        csr_reg_stvec_3_) );
  DFFSSRX1_LVT csr_reg_misa_reg_3_ ( .D(csr_n1346), .SETB(csr_wdata_5_), 
        .RSTB(csr_n590), .CLK(csr_net35137), .QN(csr_io_status_isa[3]) );
  DFFX1_LVT csr_u_T_39_reg_5_ ( .D(csr_N1433), .CLK(csr_n593), .Q(
        csr_n_T_45_5_) );
  DFFX1_LVT csr_reg_stval_reg_5_ ( .D(csr_N1387), .CLK(csr_net34930), .Q(
        csr_n_T_444[5]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_5_ ( .D(csr_n378), .SETB(csr_wdata_5_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_5_) );
  DFFX1_LVT csr_reg_satp_ppn_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[5]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[5]) );
  DFFX1_LVT csr_reg_sscratch_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[5]) );
  DFFX1_LVT csr_reg_mscratch_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[5]) );
  DFFX1_LVT csr_reg_dscratch_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[5]) );
  DFFX1_LVT csr_reg_mideleg_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_net35167), .Q(
        csr_read_mideleg_5), .QN(csr_n427) );
  DFFX1_LVT csr_reg_stvec_reg_5_ ( .D(csr_wdata_5_), .CLK(csr_n570), .Q(
        csr_reg_stvec_5_) );
  DFFX1_LVT csr_reg_mstatus_spie_reg ( .D(csr_n1914), .CLK(csr_n1915), .Q(
        csr_n1933) );
  DFFX1_LVT csr_reg_mstatus_sie_reg ( .D(csr_n1062), .CLK(csr_n1915), .Q(
        csr_n1935) );
  DFFX1_LVT csr_reg_mcause_reg_1_ ( .D(csr_N882), .CLK(csr_n580), .Q(
        csr_reg_mcause[1]) );
  DFFX1_LVT csr_u_T_47_reg_1_ ( .D(csr_N1823), .CLK(csr_n591), .Q(
        csr_io_time[1]) );
  DFFX1_LVT csr_u_T_39_reg_1_ ( .D(csr_N1429), .CLK(csr_n593), .Q(
        csr_n_T_45_1_) );
  DFFSSRX1_LVT csr_reg_bp_0_control_w_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_1_), .CLK(csr_net35314), .Q(csr_io_bp_0_control_w) );
  DFFX1_LVT csr_reg_stval_reg_1_ ( .D(csr_N1383), .CLK(csr_n561), .Q(
        csr_n_T_444[1]) );
  DFFX1_LVT csr_reg_scause_reg_1_ ( .D(csr_N1271), .CLK(csr_n558), .Q(
        csr_reg_scause[1]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[1]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[1]) );
  DFFX1_LVT csr_reg_sscratch_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[1]) );
  DFFX1_LVT csr_reg_mscratch_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[1]) );
  DFFX1_LVT csr_reg_dscratch_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[1]) );
  DFFX1_LVT csr_reg_mideleg_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_net35167), .Q(
        csr_read_mideleg_1), .QN(csr_n407) );
  DFFX1_LVT csr_reg_mcounteren_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_net34945), 
        .Q(csr_read_mcounteren_1_) );
  DFFX1_LVT csr_reg_scounteren_reg_1_ ( .D(csr_wdata_1_), .CLK(csr_net34940), 
        .Q(csr_read_scounteren_1_) );
  DFFSSRX1_LVT csr_reg_misa_reg_2_ ( .D(csr_n387), .SETB(csr_wdata_2_), .RSTB(
        csr_n590), .CLK(csr_net35137), .QN(csr_io_status_isa[2]) );
  DFFX1_LVT csr_reg_dpc_reg_4_ ( .D(csr_net35292), .CLK(csr_n530), .Q(
        csr_reg_dpc_4_) );
  DFFX1_LVT csr_reg_mepc_reg_4_ ( .D(csr_net35070), .CLK(csr_n547), .Q(
        csr_reg_mepc_4_) );
  DFFX1_LVT csr_reg_sepc_reg_4_ ( .D(csr_net34868), .CLK(csr_n583), .Q(
        csr_reg_sepc_4_) );
  DFFX1_LVT csr_reg_fflags_reg_4_ ( .D(csr_n_GEN_345[4]), .CLK(csr_n594), .Q(
        csr_read_fcsr_4_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_4_ ( .D(csr_n_GEN_307[4]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_7_addr[4]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_4_ ( .D(csr_n_GEN_300[4]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_6_addr[4]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_4_ ( .D(csr_n_GEN_293[4]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_5_addr[4]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_4_ ( .D(csr_n_GEN_286[4]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_4_addr[4]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_4_ ( .D(csr_n_GEN_279[4]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_3_addr[4]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_4_ ( .D(csr_n_GEN_272[4]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_2_addr[4]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_4_ ( .D(csr_n_GEN_265[4]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_1_addr[4]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_4_ ( .D(csr_n_GEN_258[4]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_0_addr[4]) );
  DFFX1_LVT csr_reg_mtval_reg_4_ ( .D(csr_N997), .CLK(csr_n574), .Q(
        csr_n_T_383[4]) );
  DFFX1_LVT csr_u_T_47_reg_4_ ( .D(csr_N1826), .CLK(csr_n591), .Q(
        csr_io_time[4]), .QN(csr_n454) );
  DFFX1_LVT csr_u_T_39_reg_4_ ( .D(csr_N1432), .CLK(csr_n594), .Q(
        csr_n_T_45_4_) );
  DFFSSRX1_LVT csr_reg_pmp_0_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_4_), .CLK(csr_net34905), .Q(io_ptw_pmp_0_cfg_a[1]) );
  DFFX1_LVT csr_reg_stval_reg_4_ ( .D(csr_N1386), .CLK(csr_n561), .Q(
        csr_n_T_444[4]) );
  DFFX1_LVT csr_reg_scause_reg_4_ ( .D(csr_N1274), .CLK(csr_n558), .Q(
        csr_reg_scause[4]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_4_ ( .D(csr_n378), .SETB(csr_wdata_4_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_4_) );
  DFFX1_LVT csr_reg_satp_ppn_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[4]) );
  DFFX1_LVT csr_reg_bp_0_control_s_reg ( .D(csr_wdata_4_), .CLK(csr_net35319), 
        .Q(csr_io_bp_0_control_s) );
  DFFX1_LVT csr_reg_bp_0_address_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[4]) );
  DFFX1_LVT csr_reg_sscratch_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[4]) );
  DFFX1_LVT csr_reg_mscratch_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[4]) );
  DFFX1_LVT csr_reg_dscratch_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[4]) );
  DFFX1_LVT csr_reg_medeleg_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_net35172), .Q(
        csr_read_medeleg_4_) );
  DFFX1_LVT csr_reg_stvec_reg_4_ ( .D(csr_wdata_4_), .CLK(csr_n570), .Q(
        csr_reg_stvec_4_) );
  DFFX1_LVT csr_reg_dpc_reg_8_ ( .D(csr_net35280), .CLK(csr_n530), .Q(
        csr_reg_dpc_8_) );
  DFFX1_LVT csr_reg_mepc_reg_8_ ( .D(csr_net35058), .CLK(csr_n547), .Q(
        csr_reg_mepc_8_) );
  DFFX1_LVT csr_reg_sepc_reg_8_ ( .D(csr_net34856), .CLK(csr_n583), .Q(
        csr_reg_sepc_8_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_8_ ( .D(csr_n_GEN_307[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_7_addr[8]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_8_ ( .D(csr_n_GEN_300[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_6_addr[8]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_8_ ( .D(csr_n_GEN_293[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_5_addr[8]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_8_ ( .D(csr_n_GEN_286[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_4_addr[8]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_8_ ( .D(csr_n_GEN_279[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_3_addr[8]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_8_ ( .D(csr_n_GEN_272[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_2_addr[8]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_8_ ( .D(csr_n_GEN_265[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_1_addr[8]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_8_ ( .D(csr_n_GEN_258[8]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_0_addr[8]) );
  DFFX1_LVT csr_u_T_1196_reg_0_ ( .D(csr_N1691), .CLK(csr_n594), .Q(
        io_dmem_req_bits_dprv[0]) );
  DFFX1_LVT csr_reg_dpc_reg_11_ ( .D(csr_net35271), .CLK(csr_n530), .Q(
        csr_reg_dpc_11_) );
  DFFX1_LVT csr_reg_mepc_reg_11_ ( .D(csr_net35049), .CLK(csr_n547), .Q(
        csr_reg_mepc_11_) );
  DFFX1_LVT csr_reg_sepc_reg_11_ ( .D(csr_net34847), .CLK(csr_n583), .Q(
        csr_reg_sepc_11_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_11_ ( .D(csr_n_GEN_307[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_7_addr[11]), .QN(csr_n403) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_11_ ( .D(csr_n_GEN_300[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_6_addr[11]), .QN(csr_n404) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_11_ ( .D(csr_n_GEN_293[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_5_addr[11]), .QN(csr_n399) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_11_ ( .D(csr_n_GEN_286[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_4_addr[11]), .QN(csr_n400) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_11_ ( .D(csr_n_GEN_279[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_3_addr[11]), .QN(csr_n401) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_11_ ( .D(csr_n_GEN_272[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_2_addr[11]), .QN(csr_n405) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_11_ ( .D(csr_n_GEN_265[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_1_addr[11]), .QN(csr_n402) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_11_ ( .D(csr_n_GEN_258[11]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_0_addr[11]), .QN(csr_n406) );
  DFFX1_LVT csr_reg_mie_reg_11_ ( .D(csr_N617), .CLK(csr_net34728), .Q(
        csr_reg_mie_11_) );
  DFFX1_LVT csr_u_T_49_reg_5_ ( .D(csr_N1896), .CLK(csr_n517), .Q(
        csr_io_time[11]) );
  DFFX1_LVT csr_u_T_41_reg_5_ ( .D(csr_N1502), .CLK(csr_n575), .Q(
        csr_n_T_45_11_) );
  DFFSSRX1_LVT csr_reg_pmp_1_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_11_), .CLK(csr_net35132), .Q(io_ptw_pmp_1_cfg_a[0]) );
  DFFX1_LVT csr_reg_stval_reg_11_ ( .D(csr_N1393), .CLK(csr_n561), .Q(
        csr_n_T_444[11]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_11_ ( .D(csr_n378), .SETB(csr_wdata_11_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_11_) );
  DFFX1_LVT csr_reg_mtval_reg_11_ ( .D(csr_N1004), .CLK(csr_n574), .Q(
        csr_n_T_383[11]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_11_ ( .D(csr_wdata_11_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[11]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_11_ ( .D(csr_wdata_11_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[11]) );
  DFFX1_LVT csr_reg_sscratch_reg_11_ ( .D(csr_wdata_11_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[11]) );
  DFFX1_LVT csr_reg_mscratch_reg_11_ ( .D(csr_wdata_11_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[11]) );
  DFFX1_LVT csr_reg_dscratch_reg_11_ ( .D(csr_wdata_11_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[11]) );
  DFFX1_LVT csr_reg_stvec_reg_11_ ( .D(csr_wdata_11_), .CLK(csr_n570), .Q(
        csr_reg_stvec_11_) );
  DFFX1_LVT csr_reg_mstatus_mpp_reg_0_ ( .D(csr_N333), .CLK(csr_net35147), .Q(
        csr_n_1930_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[0]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_7_ ( .D(csr_wdata_7_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[7]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[8]) );
  DFFX1_LVT csr_reg_dpc_reg_10_ ( .D(csr_net35274), .CLK(csr_n530), .Q(
        csr_reg_dpc_10_) );
  DFFX1_LVT csr_reg_mepc_reg_10_ ( .D(csr_net35052), .CLK(csr_n547), .Q(
        csr_reg_mepc_10_) );
  DFFX1_LVT csr_reg_sepc_reg_10_ ( .D(csr_net34850), .CLK(csr_n583), .Q(
        csr_reg_sepc_10_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_10_ ( .D(csr_n_GEN_307[10]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_7_addr[10]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_10_ ( .D(csr_n_GEN_300[10]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_6_addr[10]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_10_ ( .D(csr_n_GEN_293[10]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_5_addr[10]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_10_ ( .D(csr_n_GEN_286[10]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_4_addr[10]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_10_ ( .D(csr_n_GEN_279[10]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_3_addr[10]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_10_ ( .D(csr_n_GEN_272[10]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_2_addr[10]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_10_ ( .D(csr_n_GEN_265[10]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_1_addr[10]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_10_ ( .D(csr_n_GEN_258[10]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_0_addr[10]) );
  DFFX1_LVT csr_u_T_49_reg_4_ ( .D(csr_N1895), .CLK(csr_n517), .Q(
        csr_io_time[10]) );
  DFFX1_LVT csr_u_T_41_reg_4_ ( .D(csr_N1501), .CLK(csr_n575), .Q(
        csr_n_T_45_10_) );
  DFFX1_LVT csr_reg_stval_reg_10_ ( .D(csr_N1392), .CLK(csr_n561), .Q(
        csr_n_T_444[10]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_10_ ( .D(csr_n378), .SETB(csr_wdata_10_), 
        .RSTB(1'b1), .CLK(csr_n556), .QN(csr_reg_mtvec_10_) );
  DFFX1_LVT csr_reg_mtval_reg_10_ ( .D(csr_N1003), .CLK(csr_n574), .Q(
        csr_n_T_383[10]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_10_ ( .D(csr_wdata_10_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[10]) );
  DFFX1_LVT csr_reg_sscratch_reg_10_ ( .D(csr_wdata_10_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[10]) );
  DFFX1_LVT csr_reg_mscratch_reg_10_ ( .D(csr_wdata_10_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[10]) );
  DFFX1_LVT csr_reg_pmp_1_cfg_x_reg ( .D(csr_wdata_10_), .CLK(csr_net35087), 
        .Q(io_ptw_pmp_1_cfg_x) );
  DFFX1_LVT csr_reg_dscratch_reg_10_ ( .D(csr_wdata_10_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[10]) );
  DFFX1_LVT csr_reg_stvec_reg_10_ ( .D(csr_wdata_10_), .CLK(csr_n570), .Q(
        csr_reg_stvec_10_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_10_ ( .D(csr_wdata_10_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[10]) );
  DFFX1_LVT csr_reg_dpc_reg_13_ ( .D(csr_net35265), .CLK(csr_n530), .Q(
        csr_reg_dpc_13_) );
  DFFX1_LVT csr_reg_mepc_reg_13_ ( .D(csr_net35043), .CLK(csr_n547), .Q(
        csr_reg_mepc_13_) );
  DFFX1_LVT csr_reg_sepc_reg_13_ ( .D(csr_net34841), .CLK(csr_n583), .Q(
        csr_reg_sepc_13_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_13_ ( .D(csr_n_GEN_307[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_7_addr[13]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_13_ ( .D(csr_n_GEN_300[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_6_addr[13]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_13_ ( .D(csr_n_GEN_293[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_5_addr[13]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_13_ ( .D(csr_n_GEN_286[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_4_addr[13]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_13_ ( .D(csr_n_GEN_279[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_3_addr[13]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_13_ ( .D(csr_n_GEN_272[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_2_addr[13]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_13_ ( .D(csr_n_GEN_265[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_1_addr[13]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_13_ ( .D(csr_n_GEN_258[13]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_0_addr[13]) );
  DFFX1_LVT csr_reg_dpc_reg_14_ ( .D(csr_net35262), .CLK(csr_n530), .Q(
        csr_reg_dpc_14_) );
  DFFX1_LVT csr_reg_mepc_reg_14_ ( .D(csr_net35040), .CLK(csr_n547), .Q(
        csr_reg_mepc_14_) );
  DFFX1_LVT csr_reg_sepc_reg_14_ ( .D(csr_net34838), .CLK(csr_n583), .Q(
        csr_reg_sepc_14_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_14_ ( .D(csr_n_GEN_307[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_7_addr[14]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_14_ ( .D(csr_n_GEN_300[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_6_addr[14]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_14_ ( .D(csr_n_GEN_293[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_5_addr[14]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_14_ ( .D(csr_n_GEN_286[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_4_addr[14]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_14_ ( .D(csr_n_GEN_279[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_3_addr[14]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_14_ ( .D(csr_n_GEN_272[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_2_addr[14]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_14_ ( .D(csr_n_GEN_265[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_1_addr[14]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_14_ ( .D(csr_n_GEN_258[14]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_0_addr[14]) );
  DFFX1_LVT csr_u_T_49_reg_8_ ( .D(csr_N1899), .CLK(csr_n517), .Q(
        csr_io_time[14]) );
  DFFX1_LVT csr_u_T_41_reg_8_ ( .D(csr_N1505), .CLK(csr_n575), .Q(
        csr_n_T_45_14_) );
  DFFX1_LVT csr_reg_stval_reg_14_ ( .D(csr_N1396), .CLK(csr_n561), .Q(
        csr_n_T_444[14]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_14_ ( .D(csr_n378), .SETB(csr_wdata_14_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_14_) );
  DFFX1_LVT csr_reg_mtval_reg_14_ ( .D(csr_N1007), .CLK(csr_n574), .Q(
        csr_n_T_383[14]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_14_ ( .D(csr_n51), .CLK(csr_net34915), .QN(
        io_ptw_ptbr_ppn[14]) );
  DFFX1_LVT csr_reg_sscratch_reg_14_ ( .D(csr_n51), .CLK(csr_n562), .QN(
        csr_reg_sscratch[14]) );
  DFFX1_LVT csr_reg_mscratch_reg_14_ ( .D(csr_n51), .CLK(csr_n548), .QN(
        csr_reg_mscratch[14]) );
  DFFX1_LVT csr_reg_dscratch_reg_14_ ( .D(csr_n51), .CLK(csr_n522), .QN(
        csr_reg_dscratch[14]) );
  DFFX1_LVT csr_reg_stvec_reg_14_ ( .D(csr_n51), .CLK(csr_n570), .QN(
        csr_reg_stvec_14_) );
  DFFX1_LVT csr_reg_mcause_reg_63_ ( .D(csr_N944), .CLK(csr_n580), .Q(
        csr_reg_mcause[63]) );
  DFFX1_LVT csr_u_T_49_reg_57_ ( .D(csr_N1948), .CLK(csr_n517), .Q(csr_n1936)
         );
  DFFX1_LVT csr_u_T_41_reg_57_ ( .D(csr_N1554), .CLK(csr_n575), .Q(
        csr_n_T_45_63_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_2_ ( .D(csr_n_GEN_307[2]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_7_addr[2]) );
  DFFX1_LVT csr_reg_dpc_reg_29_ ( .D(csr_net35217), .CLK(csr_n530), .Q(
        csr_reg_dpc_29_) );
  DFFX1_LVT csr_reg_mepc_reg_29_ ( .D(csr_net34995), .CLK(csr_n547), .Q(
        csr_reg_mepc_29_) );
  DFFX1_LVT csr_reg_sepc_reg_29_ ( .D(csr_net34793), .CLK(csr_n583), .Q(
        csr_reg_sepc_29_) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_29_ ( .D(csr_n_GEN_300[29]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_6_addr[29]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_29_ ( .D(csr_n_GEN_293[29]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_5_addr[29]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_29_ ( .D(csr_n_GEN_286[29]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_4_addr[29]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_29_ ( .D(csr_n_GEN_279[29]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_3_addr[29]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_29_ ( .D(csr_n_GEN_272[29]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_2_addr[29]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_29_ ( .D(csr_n_GEN_265[29]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_1_addr[29]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_29_ ( .D(csr_n_GEN_258[29]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_0_addr[29]) );
  DFFX1_LVT csr_u_T_49_reg_23_ ( .D(csr_N1914), .CLK(csr_n517), .Q(
        csr_io_time[29]) );
  DFFX1_LVT csr_u_T_41_reg_23_ ( .D(csr_N1520), .CLK(csr_n575), .Q(
        csr_n_T_45_29_) );
  DFFX1_LVT csr_reg_stval_reg_29_ ( .D(csr_N1411), .CLK(csr_n561), .Q(
        csr_n_T_444[29]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_29_ ( .D(csr_n378), .SETB(csr_wdata_29_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_29_) );
  DFFX1_LVT csr_reg_mtval_reg_29_ ( .D(csr_N1022), .CLK(csr_n574), .Q(
        csr_n_T_383[29]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_29_ ( .D(csr_wdata_29_), .CLK(csr_n586), 
        .Q(csr_io_bp_0_address[29]) );
  DFFX1_LVT csr_reg_sscratch_reg_29_ ( .D(csr_wdata_29_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[29]) );
  DFFX1_LVT csr_reg_mscratch_reg_29_ ( .D(csr_wdata_29_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[29]) );
  DFFX1_LVT csr_reg_dscratch_reg_29_ ( .D(csr_wdata_29_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[29]) );
  DFFX1_LVT csr_reg_stvec_reg_29_ ( .D(csr_wdata_29_), .CLK(csr_n570), .Q(
        csr_reg_stvec_29_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_29_ ( .D(csr_n_GEN_307[29]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_7_addr[29]) );
  DFFX1_LVT csr_reg_dpc_reg_28_ ( .D(csr_net35220), .CLK(csr_n530), .Q(
        csr_reg_dpc_28_) );
  DFFX1_LVT csr_reg_mepc_reg_28_ ( .D(csr_net34998), .CLK(csr_n547), .Q(
        csr_reg_mepc_28_) );
  DFFX1_LVT csr_reg_sepc_reg_28_ ( .D(csr_net34796), .CLK(csr_n583), .Q(
        csr_reg_sepc_28_) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_28_ ( .D(csr_n_GEN_300[28]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_6_addr[28]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_28_ ( .D(csr_n_GEN_293[28]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_5_addr[28]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_28_ ( .D(csr_n_GEN_286[28]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_4_addr[28]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_28_ ( .D(csr_n_GEN_279[28]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_3_addr[28]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_28_ ( .D(csr_n_GEN_272[28]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_2_addr[28]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_28_ ( .D(csr_n_GEN_265[28]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_1_addr[28]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_28_ ( .D(csr_n_GEN_258[28]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_0_addr[28]) );
  DFFX1_LVT csr_u_T_49_reg_22_ ( .D(csr_N1913), .CLK(csr_n517), .Q(
        csr_io_time[28]) );
  DFFX1_LVT csr_u_T_41_reg_22_ ( .D(csr_N1519), .CLK(csr_n575), .Q(
        csr_n_T_45_28_) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_2_ ( .D(csr_n_GEN_272[2]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_2_addr[2]) );
  DFFX1_LVT csr_reg_dpc_reg_27_ ( .D(csr_net35223), .CLK(csr_n529), .Q(
        csr_reg_dpc_27_) );
  DFFX1_LVT csr_reg_mepc_reg_27_ ( .D(csr_net35001), .CLK(csr_n546), .Q(
        csr_reg_mepc_27_) );
  DFFX1_LVT csr_reg_sepc_reg_27_ ( .D(csr_net34799), .CLK(csr_n582), .Q(
        csr_reg_sepc_27_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_27_ ( .D(csr_n_GEN_307[27]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_7_addr[27]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_27_ ( .D(csr_n_GEN_300[27]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_6_addr[27]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_27_ ( .D(csr_n_GEN_293[27]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_5_addr[27]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_27_ ( .D(csr_n_GEN_286[27]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_4_addr[27]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_27_ ( .D(csr_n_GEN_279[27]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_3_addr[27]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_27_ ( .D(csr_n_GEN_265[27]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_1_addr[27]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_27_ ( .D(csr_n_GEN_258[27]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_0_addr[27]) );
  DFFX1_LVT csr_u_T_49_reg_21_ ( .D(csr_N1912), .CLK(csr_n517), .Q(
        csr_io_time[27]) );
  DFFX1_LVT csr_u_T_41_reg_21_ ( .D(csr_N1518), .CLK(csr_n575), .Q(
        csr_n_T_45_27_) );
  DFFSSRX1_LVT csr_reg_pmp_3_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_27_), .CLK(csr_net35127), .Q(io_ptw_pmp_3_cfg_a[0]) );
  DFFX1_LVT csr_reg_stval_reg_27_ ( .D(csr_N1409), .CLK(csr_n561), .Q(
        csr_n_T_444[27]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_27_ ( .D(csr_n378), .SETB(csr_wdata_27_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_27_) );
  DFFX1_LVT csr_reg_mtval_reg_27_ ( .D(csr_N1020), .CLK(csr_n574), .Q(
        csr_n_T_383[27]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_27_ ( .D(csr_wdata_27_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[27]) );
  DFFX1_LVT csr_reg_sscratch_reg_27_ ( .D(csr_wdata_27_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[27]) );
  DFFX1_LVT csr_reg_mscratch_reg_27_ ( .D(csr_wdata_27_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[27]) );
  DFFX1_LVT csr_reg_dscratch_reg_27_ ( .D(csr_wdata_27_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[27]) );
  DFFX1_LVT csr_reg_stvec_reg_27_ ( .D(csr_wdata_27_), .CLK(csr_n570), .Q(
        csr_reg_stvec_27_) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_27_ ( .D(csr_n_GEN_272[27]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_2_addr[27]) );
  DFFX1_LVT csr_reg_dpc_reg_26_ ( .D(csr_net35226), .CLK(csr_n529), .Q(
        csr_reg_dpc_26_) );
  DFFX1_LVT csr_reg_mepc_reg_26_ ( .D(csr_net35004), .CLK(csr_n546), .Q(
        csr_reg_mepc_26_) );
  DFFX1_LVT csr_reg_sepc_reg_26_ ( .D(csr_net34802), .CLK(csr_n582), .Q(
        csr_reg_sepc_26_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_26_ ( .D(csr_n_GEN_307[26]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_7_addr[26]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_26_ ( .D(csr_n_GEN_300[26]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_6_addr[26]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_26_ ( .D(csr_n_GEN_293[26]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_5_addr[26]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_26_ ( .D(csr_n_GEN_286[26]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_4_addr[26]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_26_ ( .D(csr_n_GEN_279[26]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_3_addr[26]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_26_ ( .D(csr_n_GEN_265[26]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_1_addr[26]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_26_ ( .D(csr_n_GEN_258[26]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_0_addr[26]) );
  DFFX1_LVT csr_u_T_49_reg_20_ ( .D(csr_N1911), .CLK(csr_n517), .Q(
        csr_io_time[26]) );
  DFFX1_LVT csr_u_T_41_reg_20_ ( .D(csr_N1517), .CLK(csr_n575), .Q(
        csr_n_T_45_26_) );
  DFFX1_LVT csr_reg_stval_reg_26_ ( .D(csr_N1408), .CLK(csr_n561), .Q(
        csr_n_T_444[26]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_26_ ( .D(csr_n378), .SETB(csr_wdata_26_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_26_) );
  DFFX1_LVT csr_reg_mtval_reg_26_ ( .D(csr_N1019), .CLK(csr_n574), .Q(
        csr_n_T_383[26]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_26_ ( .D(csr_wdata_26_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[26]) );
  DFFX1_LVT csr_reg_sscratch_reg_26_ ( .D(csr_wdata_26_), .CLK(csr_n562), .Q(
        csr_reg_sscratch[26]) );
  DFFX1_LVT csr_reg_mscratch_reg_26_ ( .D(csr_wdata_26_), .CLK(csr_n548), .Q(
        csr_reg_mscratch[26]) );
  DFFX1_LVT csr_reg_pmp_3_cfg_x_reg ( .D(csr_wdata_26_), .CLK(csr_net35122), 
        .Q(io_ptw_pmp_3_cfg_x) );
  DFFX1_LVT csr_reg_dscratch_reg_26_ ( .D(csr_wdata_26_), .CLK(csr_n522), .Q(
        csr_reg_dscratch[26]) );
  DFFX1_LVT csr_reg_stvec_reg_26_ ( .D(csr_wdata_26_), .CLK(csr_n570), .Q(
        csr_reg_stvec_26_) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_26_ ( .D(csr_n_GEN_272[26]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_2_addr[26]) );
  DFFX1_LVT csr_reg_dpc_reg_25_ ( .D(csr_net35229), .CLK(csr_n529), .Q(
        csr_reg_dpc_25_) );
  DFFX1_LVT csr_reg_mepc_reg_25_ ( .D(csr_net35007), .CLK(csr_n546), .Q(
        csr_reg_mepc_25_) );
  DFFX1_LVT csr_reg_sepc_reg_25_ ( .D(csr_net34805), .CLK(csr_n582), .Q(
        csr_reg_sepc_25_) );
  DFFSSRX1_LVT csr_reg_pmp_3_cfg_w_reg ( .D(csr_wdata_24_), .SETB(1'b1), 
        .RSTB(csr_wdata_25_), .CLK(csr_net35122), .Q(io_ptw_pmp_3_cfg_w) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_25_ ( .D(csr_n_GEN_307[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_7_addr[25]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_25_ ( .D(csr_n_GEN_300[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_6_addr[25]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_25_ ( .D(csr_n_GEN_293[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_5_addr[25]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_25_ ( .D(csr_n_GEN_286[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_4_addr[25]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_25_ ( .D(csr_n_GEN_279[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_3_addr[25]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_25_ ( .D(csr_n_GEN_265[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_1_addr[25]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_25_ ( .D(csr_n_GEN_258[25]), .CLK(csr_n541), 
        .Q(io_ptw_pmp_0_addr[25]) );
  DFFX1_LVT csr_u_T_49_reg_19_ ( .D(csr_N1910), .CLK(csr_n517), .Q(
        csr_io_time[25]) );
  DFFX1_LVT csr_u_T_41_reg_19_ ( .D(csr_N1516), .CLK(csr_n575), .Q(
        csr_n_T_45_25_) );
  DFFX1_LVT csr_reg_stval_reg_25_ ( .D(csr_N1407), .CLK(csr_n561), .Q(
        csr_n_T_444[25]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_25_ ( .D(csr_n378), .SETB(csr_wdata_25_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_25_) );
  DFFX1_LVT csr_reg_mtval_reg_25_ ( .D(csr_N1018), .CLK(csr_n574), .Q(
        csr_n_T_383[25]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_25_ ( .D(csr_wdata_25_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[25]) );
  DFFX1_LVT csr_reg_sscratch_reg_25_ ( .D(csr_wdata_25_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[25]) );
  DFFX1_LVT csr_reg_mscratch_reg_25_ ( .D(csr_wdata_25_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[25]) );
  DFFX1_LVT csr_reg_dscratch_reg_25_ ( .D(csr_wdata_25_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[25]) );
  DFFX1_LVT csr_reg_stvec_reg_25_ ( .D(csr_wdata_25_), .CLK(csr_n570), .Q(
        csr_reg_stvec_25_) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_25_ ( .D(csr_n_GEN_272[25]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_2_addr[25]) );
  DFFX1_LVT csr_reg_dpc_reg_24_ ( .D(csr_net35232), .CLK(csr_n529), .Q(
        csr_reg_dpc_24_) );
  DFFX1_LVT csr_reg_mepc_reg_24_ ( .D(csr_net35010), .CLK(csr_n546), .Q(
        csr_reg_mepc_24_) );
  DFFX1_LVT csr_reg_sepc_reg_24_ ( .D(csr_net34808), .CLK(csr_n582), .Q(
        csr_reg_sepc_24_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_24_ ( .D(csr_n_GEN_307[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_7_addr[24]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_24_ ( .D(csr_n_GEN_300[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_6_addr[24]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_24_ ( .D(csr_n_GEN_293[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_5_addr[24]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_24_ ( .D(csr_n_GEN_286[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_4_addr[24]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_24_ ( .D(csr_n_GEN_279[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_3_addr[24]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_24_ ( .D(csr_n_GEN_265[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_1_addr[24]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_24_ ( .D(csr_n_GEN_258[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_0_addr[24]) );
  DFFX1_LVT csr_u_T_49_reg_18_ ( .D(csr_N1909), .CLK(csr_n517), .Q(
        csr_io_time[24]) );
  DFFX1_LVT csr_u_T_41_reg_18_ ( .D(csr_N1515), .CLK(csr_n575), .Q(
        csr_n_T_45_24_) );
  DFFX1_LVT csr_reg_stval_reg_24_ ( .D(csr_N1406), .CLK(csr_n561), .Q(
        csr_n_T_444[24]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_24_ ( .D(csr_n378), .SETB(csr_wdata_24_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_24_) );
  DFFX1_LVT csr_reg_mtval_reg_24_ ( .D(csr_N1017), .CLK(csr_n574), .Q(
        csr_n_T_383[24]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_24_ ( .D(csr_wdata_24_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[24]) );
  DFFX1_LVT csr_reg_sscratch_reg_24_ ( .D(csr_wdata_24_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[24]) );
  DFFX1_LVT csr_reg_mscratch_reg_24_ ( .D(csr_wdata_24_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[24]) );
  DFFX1_LVT csr_reg_pmp_3_cfg_r_reg ( .D(csr_wdata_24_), .CLK(csr_net35122), 
        .Q(io_ptw_pmp_3_cfg_r) );
  DFFX1_LVT csr_reg_dscratch_reg_24_ ( .D(csr_wdata_24_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[24]) );
  DFFX1_LVT csr_reg_stvec_reg_24_ ( .D(csr_wdata_24_), .CLK(csr_n570), .Q(
        csr_reg_stvec_24_) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_24_ ( .D(csr_n_GEN_272[24]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_2_addr[24]) );
  DFFX1_LVT csr_reg_dpc_reg_23_ ( .D(csr_net35235), .CLK(csr_n529), .Q(
        csr_reg_dpc_23_) );
  DFFX1_LVT csr_reg_mepc_reg_23_ ( .D(csr_net35013), .CLK(csr_n546), .Q(
        csr_reg_mepc_23_) );
  DFFX1_LVT csr_reg_sepc_reg_23_ ( .D(csr_net34811), .CLK(csr_n582), .Q(
        csr_reg_sepc_23_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_23_ ( .D(csr_n_GEN_307[23]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_7_addr[23]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_23_ ( .D(csr_n_GEN_300[23]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_6_addr[23]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_23_ ( .D(csr_n_GEN_293[23]), .CLK(csr_n542), 
        .Q(io_ptw_pmp_5_addr[23]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_23_ ( .D(csr_n_GEN_286[23]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_4_addr[23]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_23_ ( .D(csr_n_GEN_279[23]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_3_addr[23]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_23_ ( .D(csr_n_GEN_265[23]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_1_addr[23]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_23_ ( .D(csr_n_GEN_258[23]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_0_addr[23]) );
  DFFX1_LVT csr_u_T_49_reg_17_ ( .D(csr_N1908), .CLK(csr_n518), .Q(
        csr_io_time[23]) );
  DFFX1_LVT csr_u_T_41_reg_17_ ( .D(csr_N1514), .CLK(csr_n576), .Q(
        csr_n_T_45_23_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_2_ ( .D(csr_n_GEN_265[2]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_1_addr[2]) );
  DFFX1_LVT csr_reg_dpc_reg_22_ ( .D(csr_net35238), .CLK(csr_n529), .Q(
        csr_reg_dpc_22_) );
  DFFX1_LVT csr_reg_mepc_reg_22_ ( .D(csr_net35016), .CLK(csr_n546), .Q(
        csr_reg_mepc_22_) );
  DFFX1_LVT csr_reg_sepc_reg_22_ ( .D(csr_net34814), .CLK(csr_n582), .Q(
        csr_reg_sepc_22_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_22_ ( .D(csr_n_GEN_307[22]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_7_addr[22]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_22_ ( .D(csr_n_GEN_300[22]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_6_addr[22]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_22_ ( .D(csr_n_GEN_293[22]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_5_addr[22]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_22_ ( .D(csr_n_GEN_286[22]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_4_addr[22]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_22_ ( .D(csr_n_GEN_279[22]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_3_addr[22]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_22_ ( .D(csr_n_GEN_272[22]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_2_addr[22]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_22_ ( .D(csr_n_GEN_258[22]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_0_addr[22]) );
  DFFX1_LVT csr_u_T_49_reg_16_ ( .D(csr_N1907), .CLK(csr_n518), .Q(
        csr_io_time[22]) );
  DFFX1_LVT csr_u_T_41_reg_16_ ( .D(csr_N1513), .CLK(csr_n576), .Q(
        csr_n_T_45_22_) );
  DFFSSRX1_LVT csr_reg_mstatus_tsr_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_22_), .CLK(csr_net35152), .Q(csr_n1924) );
  DFFX1_LVT csr_reg_stval_reg_22_ ( .D(csr_N1404), .CLK(csr_n561), .Q(
        csr_n_T_444[22]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_22_ ( .D(csr_n378), .SETB(csr_wdata_22_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_22_) );
  DFFX1_LVT csr_reg_mtval_reg_22_ ( .D(csr_N1015), .CLK(csr_n574), .Q(
        csr_n_T_383[22]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_22_ ( .D(csr_wdata_22_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[22]) );
  DFFX1_LVT csr_reg_sscratch_reg_22_ ( .D(csr_wdata_22_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[22]) );
  DFFX1_LVT csr_reg_mscratch_reg_22_ ( .D(csr_wdata_22_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[22]) );
  DFFX1_LVT csr_reg_dscratch_reg_22_ ( .D(csr_wdata_22_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[22]) );
  DFFX1_LVT csr_reg_stvec_reg_22_ ( .D(csr_wdata_22_), .CLK(csr_n570), .Q(
        csr_reg_stvec_22_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_22_ ( .D(csr_n_GEN_265[22]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_1_addr[22]) );
  DFFX1_LVT csr_reg_dpc_reg_21_ ( .D(csr_net35241), .CLK(csr_n529), .Q(
        csr_reg_dpc_21_) );
  DFFX1_LVT csr_reg_mepc_reg_21_ ( .D(csr_net35019), .CLK(csr_n546), .Q(
        csr_reg_mepc_21_) );
  DFFX1_LVT csr_reg_sepc_reg_21_ ( .D(csr_net34817), .CLK(csr_n582), .Q(
        csr_reg_sepc_21_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_21_ ( .D(csr_n_GEN_307[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_7_addr[21]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_21_ ( .D(csr_n_GEN_300[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_6_addr[21]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_21_ ( .D(csr_n_GEN_293[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_5_addr[21]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_21_ ( .D(csr_n_GEN_286[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_4_addr[21]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_21_ ( .D(csr_n_GEN_279[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_3_addr[21]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_21_ ( .D(csr_n_GEN_272[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_2_addr[21]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_21_ ( .D(csr_n_GEN_258[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_0_addr[21]) );
  DFFX1_LVT csr_u_T_49_reg_15_ ( .D(csr_N1906), .CLK(csr_n518), .Q(
        csr_io_time[21]) );
  DFFX1_LVT csr_u_T_41_reg_15_ ( .D(csr_N1512), .CLK(csr_n576), .Q(
        csr_n_T_45_21_) );
  DFFSSRX1_LVT csr_reg_mstatus_tw_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_21_), .CLK(csr_net35152), .Q(csr_n1925) );
  DFFX1_LVT csr_reg_stval_reg_21_ ( .D(csr_N1403), .CLK(csr_n561), .Q(
        csr_n_T_444[21]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_21_ ( .D(csr_n378), .SETB(csr_wdata_21_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_21_) );
  DFFX1_LVT csr_reg_mtval_reg_21_ ( .D(csr_N1014), .CLK(csr_n574), .Q(
        csr_n_T_383[21]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_21_ ( .D(csr_wdata_21_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[21]) );
  DFFX1_LVT csr_reg_sscratch_reg_21_ ( .D(csr_wdata_21_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[21]) );
  DFFX1_LVT csr_reg_mscratch_reg_21_ ( .D(csr_wdata_21_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[21]) );
  DFFX1_LVT csr_reg_dscratch_reg_21_ ( .D(csr_wdata_21_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[21]) );
  DFFX1_LVT csr_reg_stvec_reg_21_ ( .D(csr_wdata_21_), .CLK(csr_n570), .Q(
        csr_reg_stvec_21_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_21_ ( .D(csr_n_GEN_265[21]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_1_addr[21]) );
  DFFX1_LVT csr_reg_dpc_reg_20_ ( .D(csr_net35244), .CLK(csr_n529), .Q(
        csr_reg_dpc_20_) );
  DFFX1_LVT csr_reg_mepc_reg_20_ ( .D(csr_net35022), .CLK(csr_n546), .Q(
        csr_reg_mepc_20_) );
  DFFX1_LVT csr_reg_sepc_reg_20_ ( .D(csr_net34820), .CLK(csr_n582), .Q(
        csr_reg_sepc_20_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_20_ ( .D(csr_n_GEN_307[20]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_7_addr[20]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_20_ ( .D(csr_n_GEN_300[20]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_6_addr[20]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_20_ ( .D(csr_n_GEN_293[20]), .CLK(csr_n543), 
        .Q(io_ptw_pmp_5_addr[20]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_20_ ( .D(csr_n_GEN_286[20]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_4_addr[20]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_20_ ( .D(csr_n_GEN_279[20]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_3_addr[20]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_20_ ( .D(csr_n_GEN_272[20]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_2_addr[20]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_20_ ( .D(csr_n_GEN_258[20]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_0_addr[20]) );
  DFFSSRX1_LVT csr_reg_mstatus_tvm_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_20_), .CLK(csr_net35152), .Q(csr_n1926), .QN(csr_n447) );
  DFFX1_LVT csr_u_T_41_reg_14_ ( .D(csr_N1511), .CLK(csr_n576), .Q(
        csr_n_T_45_20_) );
  DFFX1_LVT csr_u_T_49_reg_14_ ( .D(csr_N1905), .CLK(csr_n518), .Q(
        csr_io_time[20]) );
  DFFSSRX1_LVT csr_reg_pmp_2_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_20_), .CLK(csr_net34753), .Q(io_ptw_pmp_2_cfg_a[1]), .QN(
        csr_n463) );
  DFFX1_LVT csr_reg_stval_reg_20_ ( .D(csr_N1402), .CLK(csr_n560), .Q(
        csr_n_T_444[20]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_20_ ( .D(csr_n378), .SETB(csr_wdata_20_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_20_) );
  DFFX1_LVT csr_reg_mtval_reg_20_ ( .D(csr_N1013), .CLK(csr_n573), .Q(
        csr_n_T_383[20]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_20_ ( .D(csr_wdata_20_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[20]) );
  DFFX1_LVT csr_reg_sscratch_reg_20_ ( .D(csr_wdata_20_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[20]) );
  DFFX1_LVT csr_reg_mscratch_reg_20_ ( .D(csr_wdata_20_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[20]) );
  DFFX1_LVT csr_reg_dscratch_reg_20_ ( .D(csr_wdata_20_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[20]) );
  DFFX1_LVT csr_reg_stvec_reg_20_ ( .D(csr_wdata_20_), .CLK(csr_n569), .Q(
        csr_reg_stvec_20_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_20_ ( .D(csr_n_GEN_265[20]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_1_addr[20]) );
  DFFX1_LVT csr_reg_dpc_reg_19_ ( .D(csr_net35247), .CLK(csr_n529), .Q(
        csr_reg_dpc_19_) );
  DFFX1_LVT csr_reg_mepc_reg_19_ ( .D(csr_net35025), .CLK(csr_n546), .Q(
        csr_reg_mepc_19_) );
  DFFX1_LVT csr_reg_sepc_reg_19_ ( .D(csr_net34823), .CLK(csr_n582), .Q(
        csr_reg_sepc_19_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_19_ ( .D(csr_n_GEN_307[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_7_addr[19]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_19_ ( .D(csr_n_GEN_300[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_6_addr[19]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_19_ ( .D(csr_n_GEN_293[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_5_addr[19]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_19_ ( .D(csr_n_GEN_286[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_4_addr[19]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_19_ ( .D(csr_n_GEN_279[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_3_addr[19]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_19_ ( .D(csr_n_GEN_272[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_2_addr[19]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_19_ ( .D(csr_n_GEN_258[19]), .CLK(csr_n544), 
        .Q(io_ptw_pmp_0_addr[19]) );
  DFFSSRX1_LVT csr_reg_mstatus_mxr_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_19_), .CLK(csr_net35157), .Q(io_ptw_status_mxr) );
  DFFX1_LVT csr_u_T_41_reg_13_ ( .D(csr_N1510), .CLK(csr_n576), .Q(
        csr_n_T_45_19_) );
  DFFX1_LVT csr_u_T_49_reg_13_ ( .D(csr_N1904), .CLK(csr_n518), .Q(
        csr_io_time[19]) );
  DFFX1_LVT csr_reg_stval_reg_19_ ( .D(csr_N1401), .CLK(csr_n560), .Q(
        csr_n_T_444[19]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_19_ ( .D(csr_n378), .SETB(csr_wdata_19_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_19_) );
  DFFX1_LVT csr_reg_mtval_reg_19_ ( .D(csr_N1012), .CLK(csr_n573), .Q(
        csr_n_T_383[19]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_19_ ( .D(csr_wdata_19_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[19]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_19_ ( .D(csr_wdata_19_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[19]) );
  DFFX1_LVT csr_reg_sscratch_reg_19_ ( .D(csr_wdata_19_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[19]) );
  DFFX1_LVT csr_reg_mscratch_reg_19_ ( .D(csr_wdata_19_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[19]) );
  DFFX1_LVT csr_reg_dscratch_reg_19_ ( .D(csr_wdata_19_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[19]) );
  DFFX1_LVT csr_reg_stvec_reg_19_ ( .D(csr_wdata_19_), .CLK(csr_n569), .Q(
        csr_reg_stvec_19_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_19_ ( .D(csr_n_GEN_265[19]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_1_addr[19]) );
  DFFX1_LVT csr_reg_dpc_reg_18_ ( .D(csr_net35250), .CLK(csr_n529), .Q(
        csr_reg_dpc_18_) );
  DFFX1_LVT csr_reg_mepc_reg_18_ ( .D(csr_net35028), .CLK(csr_n546), .Q(
        csr_reg_mepc_18_) );
  DFFX1_LVT csr_reg_sepc_reg_18_ ( .D(csr_net34826), .CLK(csr_n582), .Q(
        csr_reg_sepc_18_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_18_ ( .D(csr_n_GEN_307[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_7_addr[18]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_18_ ( .D(csr_n_GEN_300[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_6_addr[18]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_18_ ( .D(csr_n_GEN_293[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_5_addr[18]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_18_ ( .D(csr_n_GEN_286[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_4_addr[18]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_18_ ( .D(csr_n_GEN_279[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_3_addr[18]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_18_ ( .D(csr_n_GEN_272[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_2_addr[18]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_18_ ( .D(csr_n_GEN_258[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_0_addr[18]) );
  DFFX1_LVT csr_u_T_49_reg_12_ ( .D(csr_N1903), .CLK(csr_n518), .Q(
        csr_io_time[18]) );
  DFFX1_LVT csr_u_T_41_reg_12_ ( .D(csr_N1509), .CLK(csr_n576), .Q(
        csr_n_T_45_18_) );
  DFFSSRX1_LVT csr_reg_mstatus_sum_reg ( .D(csr_n503), .SETB(1'b1), .RSTB(
        csr_wdata_18_), .CLK(csr_net35157), .Q(io_ptw_status_sum) );
  DFFX1_LVT csr_reg_stval_reg_18_ ( .D(csr_N1400), .CLK(csr_n560), .Q(
        csr_n_T_444[18]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_18_ ( .D(csr_n378), .SETB(csr_wdata_18_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_18_) );
  DFFX1_LVT csr_reg_mtval_reg_18_ ( .D(csr_N1011), .CLK(csr_n573), .Q(
        csr_n_T_383[18]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_18_ ( .D(csr_wdata_18_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[18]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_18_ ( .D(csr_wdata_18_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[18]) );
  DFFX1_LVT csr_reg_sscratch_reg_18_ ( .D(csr_wdata_18_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[18]) );
  DFFX1_LVT csr_reg_mscratch_reg_18_ ( .D(csr_wdata_18_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[18]) );
  DFFX1_LVT csr_reg_pmp_2_cfg_x_reg ( .D(csr_wdata_18_), .CLK(csr_net34748), 
        .Q(io_ptw_pmp_2_cfg_x) );
  DFFX1_LVT csr_reg_dscratch_reg_18_ ( .D(csr_wdata_18_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[18]) );
  DFFX1_LVT csr_reg_stvec_reg_18_ ( .D(csr_wdata_18_), .CLK(csr_n569), .Q(
        csr_reg_stvec_18_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_18_ ( .D(csr_n_GEN_265[18]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_1_addr[18]) );
  DFFX1_LVT csr_reg_dpc_reg_17_ ( .D(csr_net35253), .CLK(csr_n529), .Q(
        csr_reg_dpc_17_) );
  DFFX1_LVT csr_reg_mepc_reg_17_ ( .D(csr_net35031), .CLK(csr_n546), .Q(
        csr_reg_mepc_17_) );
  DFFX1_LVT csr_reg_sepc_reg_17_ ( .D(csr_net34829), .CLK(csr_n582), .Q(
        csr_reg_sepc_17_) );
  DFFSSRX1_LVT csr_reg_pmp_2_cfg_w_reg ( .D(csr_wdata_17_), .SETB(1'b1), 
        .RSTB(csr_wdata_16_), .CLK(csr_net34748), .Q(io_ptw_pmp_2_cfg_w) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_17_ ( .D(csr_n_GEN_307[17]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_7_addr[17]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_17_ ( .D(csr_n_GEN_300[17]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_6_addr[17]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_17_ ( .D(csr_n_GEN_293[17]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_5_addr[17]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_17_ ( .D(csr_n_GEN_286[17]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_4_addr[17]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_17_ ( .D(csr_n_GEN_279[17]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_3_addr[17]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_17_ ( .D(csr_n_GEN_272[17]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_2_addr[17]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_17_ ( .D(csr_n_GEN_258[17]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_0_addr[17]) );
  DFFX1_LVT csr_u_T_49_reg_11_ ( .D(csr_N1902), .CLK(csr_n518), .Q(
        csr_io_time[17]) );
  DFFX1_LVT csr_u_T_41_reg_11_ ( .D(csr_N1508), .CLK(csr_n576), .Q(
        csr_n_T_45_17_) );
  DFFSSRX1_LVT csr_reg_mstatus_mprv_reg ( .D(csr_n503), .SETB(1'b1), .RSTB(
        csr_wdata_17_), .CLK(csr_net35152), .Q(csr_n1927) );
  DFFX1_LVT csr_reg_stval_reg_17_ ( .D(csr_N1399), .CLK(csr_n560), .Q(
        csr_n_T_444[17]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_17_ ( .D(csr_n378), .SETB(csr_wdata_17_), 
        .RSTB(1'b1), .CLK(csr_n555), .QN(csr_reg_mtvec_17_) );
  DFFX1_LVT csr_reg_mtval_reg_17_ ( .D(csr_N1010), .CLK(csr_n573), .Q(
        csr_n_T_383[17]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_17_ ( .D(csr_wdata_17_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[17]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_17_ ( .D(csr_wdata_17_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[17]) );
  DFFX1_LVT csr_reg_sscratch_reg_17_ ( .D(csr_wdata_17_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[17]) );
  DFFX1_LVT csr_reg_mscratch_reg_17_ ( .D(csr_wdata_17_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[17]) );
  DFFX1_LVT csr_reg_dscratch_reg_17_ ( .D(csr_wdata_17_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[17]) );
  DFFX1_LVT csr_reg_stvec_reg_17_ ( .D(csr_wdata_17_), .CLK(csr_n569), .Q(
        csr_reg_stvec_17_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_17_ ( .D(csr_n_GEN_265[17]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_1_addr[17]) );
  DFFX1_LVT csr_reg_dpc_reg_16_ ( .D(csr_net35256), .CLK(csr_n529), .Q(
        csr_reg_dpc_16_) );
  DFFX1_LVT csr_reg_mepc_reg_16_ ( .D(csr_net35034), .CLK(csr_n546), .Q(
        csr_reg_mepc_16_) );
  DFFX1_LVT csr_reg_sepc_reg_16_ ( .D(csr_net34832), .CLK(csr_n582), .Q(
        csr_reg_sepc_16_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_16_ ( .D(csr_n_GEN_307[16]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_7_addr[16]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_16_ ( .D(csr_n_GEN_300[16]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_6_addr[16]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_16_ ( .D(csr_n_GEN_293[16]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_5_addr[16]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_16_ ( .D(csr_n_GEN_286[16]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_4_addr[16]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_16_ ( .D(csr_n_GEN_279[16]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_3_addr[16]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_16_ ( .D(csr_n_GEN_272[16]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_2_addr[16]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_16_ ( .D(csr_n_GEN_258[16]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_0_addr[16]) );
  DFFX1_LVT csr_u_T_49_reg_10_ ( .D(csr_N1901), .CLK(csr_n518), .Q(
        csr_io_time[16]) );
  DFFX1_LVT csr_u_T_41_reg_10_ ( .D(csr_N1507), .CLK(csr_n576), .Q(
        csr_n_T_45_16_) );
  DFFX1_LVT csr_reg_stval_reg_16_ ( .D(csr_N1398), .CLK(csr_n560), .Q(
        csr_n_T_444[16]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_16_ ( .D(csr_n378), .SETB(csr_wdata_16_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_16_) );
  DFFX1_LVT csr_reg_mtval_reg_16_ ( .D(csr_N1009), .CLK(csr_n573), .Q(
        csr_n_T_383[16]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_16_ ( .D(csr_wdata_16_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[16]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_16_ ( .D(csr_wdata_16_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[16]) );
  DFFX1_LVT csr_reg_sscratch_reg_16_ ( .D(csr_wdata_16_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[16]) );
  DFFX1_LVT csr_reg_mscratch_reg_16_ ( .D(csr_wdata_16_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[16]) );
  DFFX1_LVT csr_reg_pmp_2_cfg_r_reg ( .D(csr_wdata_16_), .CLK(csr_net34748), 
        .Q(io_ptw_pmp_2_cfg_r) );
  DFFX1_LVT csr_reg_dscratch_reg_16_ ( .D(csr_wdata_16_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[16]) );
  DFFX1_LVT csr_reg_stvec_reg_16_ ( .D(csr_wdata_16_), .CLK(csr_n569), .Q(
        csr_reg_stvec_16_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_16_ ( .D(csr_n_GEN_265[16]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_1_addr[16]) );
  DFFX1_LVT csr_reg_dpc_reg_15_ ( .D(csr_net35259), .CLK(csr_n528), .Q(
        csr_reg_dpc_15_) );
  DFFX1_LVT csr_reg_mepc_reg_15_ ( .D(csr_net35037), .CLK(csr_n545), .Q(
        csr_reg_mepc_15_) );
  DFFX1_LVT csr_reg_sepc_reg_15_ ( .D(csr_net34835), .CLK(csr_n581), .Q(
        csr_reg_sepc_15_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_15_ ( .D(csr_n_GEN_307[15]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_7_addr[15]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_15_ ( .D(csr_n_GEN_300[15]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_6_addr[15]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_15_ ( .D(csr_n_GEN_293[15]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_5_addr[15]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_15_ ( .D(csr_n_GEN_286[15]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_4_addr[15]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_15_ ( .D(csr_n_GEN_279[15]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_3_addr[15]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_15_ ( .D(csr_n_GEN_272[15]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_2_addr[15]) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_15_ ( .D(csr_n_GEN_258[15]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_0_addr[15]) );
  DFFSSRX1_LVT csr_reg_dcsr_ebreakm_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_15_), .CLK(csr_net35162), .Q(csr_n_T_1155_3) );
  DFFX1_LVT csr_u_T_41_reg_9_ ( .D(csr_N1506), .CLK(csr_n576), .Q(
        csr_n_T_45_15_) );
  DFFX1_LVT csr_u_T_49_reg_9_ ( .D(csr_N1900), .CLK(csr_n518), .Q(
        csr_io_time[15]) );
  DFFX1_LVT csr_reg_pmp_1_cfg_r_reg ( .D(csr_wdata_8_), .CLK(csr_net35087), 
        .Q(io_ptw_pmp_1_cfg_r) );
  DFFSSRX1_LVT csr_reg_pmp_1_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_15_), .CLK(csr_net35132), .Q(io_ptw_pmp_1_cfg_l), .QN(
        csr_n440) );
  DFFX1_LVT csr_reg_stval_reg_15_ ( .D(csr_N1397), .CLK(csr_n560), .Q(
        csr_n_T_444[15]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_15_ ( .D(csr_n376), .SETB(csr_wdata_15_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_15_) );
  DFFX1_LVT csr_reg_mtval_reg_15_ ( .D(csr_N1008), .CLK(csr_n573), .Q(
        csr_n_T_383[15]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[15]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_n585), 
        .Q(csr_io_bp_0_address[15]) );
  DFFX1_LVT csr_reg_sscratch_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[15]) );
  DFFX1_LVT csr_reg_mscratch_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[15]) );
  DFFX1_LVT csr_reg_dscratch_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[15]) );
  DFFX1_LVT csr_reg_medeleg_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_net35172), 
        .Q(csr_read_medeleg_15) );
  DFFX1_LVT csr_reg_stvec_reg_15_ ( .D(csr_wdata_15_), .CLK(csr_n569), .Q(
        csr_reg_stvec_15_) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_15_ ( .D(csr_n_GEN_265[15]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_1_addr[15]) );
  DFFX1_LVT csr_reg_pmp_1_addr_reg_0_ ( .D(csr_n_GEN_265[0]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_1_addr[0]) );
  DFFSSRX1_LVT csr_reg_pmp_2_cfg_a_reg_0_ ( .D(csr_n503), .SETB(1'b1), .RSTB(
        csr_wdata_19_), .CLK(csr_net34753), .Q(io_ptw_pmp_2_cfg_a[0]) );
  DFFSSRX1_LVT csr_reg_pmp_2_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_23_), .CLK(csr_net34753), .Q(io_ptw_pmp_2_cfg_l), .QN(
        csr_n441) );
  DFFX1_LVT csr_reg_stval_reg_23_ ( .D(csr_N1405), .CLK(csr_n560), .Q(
        csr_n_T_444[23]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_23_ ( .D(csr_n376), .SETB(csr_wdata_23_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_23_) );
  DFFX1_LVT csr_reg_mtval_reg_23_ ( .D(csr_N1016), .CLK(csr_n573), .Q(
        csr_n_T_383[23]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_23_ ( .D(csr_wdata_23_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[23]) );
  DFFX1_LVT csr_reg_sscratch_reg_23_ ( .D(csr_wdata_23_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[23]) );
  DFFX1_LVT csr_reg_mscratch_reg_23_ ( .D(csr_wdata_23_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[23]) );
  DFFX1_LVT csr_reg_dscratch_reg_23_ ( .D(csr_wdata_23_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[23]) );
  DFFX1_LVT csr_reg_stvec_reg_23_ ( .D(csr_wdata_23_), .CLK(csr_n569), .Q(
        csr_reg_stvec_23_) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_23_ ( .D(csr_n_GEN_272[23]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_2_addr[23]) );
  DFFX1_LVT csr_reg_pmp_2_addr_reg_0_ ( .D(csr_n_GEN_272[0]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_2_addr[0]) );
  DFFSSRX1_LVT csr_reg_pmp_3_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_28_), .CLK(csr_net35127), .Q(io_ptw_pmp_3_cfg_a[1]), .QN(
        csr_n460) );
  DFFX1_LVT csr_reg_stval_reg_28_ ( .D(csr_N1410), .CLK(csr_n560), .Q(
        csr_n_T_444[28]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_28_ ( .D(csr_n376), .SETB(csr_wdata_28_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_28_) );
  DFFX1_LVT csr_reg_mtval_reg_28_ ( .D(csr_N1021), .CLK(csr_n573), .Q(
        csr_n_T_383[28]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_28_ ( .D(csr_wdata_28_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[28]) );
  DFFX1_LVT csr_reg_sscratch_reg_28_ ( .D(csr_wdata_28_), .CLK(csr_n563), .Q(
        csr_reg_sscratch[28]) );
  DFFX1_LVT csr_reg_mscratch_reg_28_ ( .D(csr_wdata_28_), .CLK(csr_n549), .Q(
        csr_reg_mscratch[28]) );
  DFFX1_LVT csr_reg_dscratch_reg_28_ ( .D(csr_wdata_28_), .CLK(csr_n523), .Q(
        csr_reg_dscratch[28]) );
  DFFX1_LVT csr_reg_stvec_reg_28_ ( .D(csr_wdata_28_), .CLK(csr_n569), .Q(
        csr_reg_stvec_28_) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_28_ ( .D(csr_n_GEN_307[28]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_7_addr[28]) );
  DFFX1_LVT csr_reg_pmp_7_addr_reg_0_ ( .D(csr_n_GEN_307[0]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_7_addr[0]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_2_ ( .D(csr_n_GEN_300[2]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_6_addr[2]) );
  DFFX1_LVT csr_reg_pmp_6_addr_reg_0_ ( .D(csr_n_GEN_300[0]), .CLK(csr_n535), 
        .Q(io_ptw_pmp_6_addr[0]) );
  DFFX1_LVT csr_u_T_49_reg_53_ ( .D(csr_N1944), .CLK(csr_n518), .Q(csr_n1940)
         );
  DFFX1_LVT csr_u_T_41_reg_53_ ( .D(csr_N1550), .CLK(csr_n576), .Q(
        csr_n_T_45_59_) );
  DFFX1_LVT csr_reg_sscratch_reg_59_ ( .D(csr_wdata_59_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[59]) );
  DFFX1_LVT csr_reg_mscratch_reg_59_ ( .D(csr_wdata_59_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[59]) );
  DFFX1_LVT csr_reg_dscratch_reg_59_ ( .D(csr_wdata_59_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[59]) );
  DFFSSRX1_LVT csr_reg_pmp_7_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_59_), .CLK(csr_net34743), .Q(io_ptw_pmp_7_cfg_a[0]) );
  DFFX1_LVT csr_u_T_49_reg_54_ ( .D(csr_N1945), .CLK(csr_n518), .Q(csr_n1939)
         );
  DFFX1_LVT csr_u_T_41_reg_54_ ( .D(csr_N1551), .CLK(csr_n576), .Q(
        csr_n_T_45_60_) );
  DFFX1_LVT csr_reg_satp_mode_reg_3_ ( .D(csr_wdata_63_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_mode[3]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[0]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_2_ ( .D(csr_n1483), .CLK(csr_net34915), .QN(
        io_ptw_ptbr_ppn[2]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_7_ ( .D(csr_wdata_7_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[7]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[8]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_12_ ( .D(csr_n367), .CLK(csr_net34915), .QN(
        io_ptw_ptbr_ppn[12]) );
  DFFX1_LVT csr_reg_satp_ppn_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_net34915), 
        .Q(io_ptw_ptbr_ppn[13]) );
  DFFX1_LVT csr_reg_sscratch_reg_60_ ( .D(csr_wdata_60_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[60]) );
  DFFX1_LVT csr_reg_mscratch_reg_60_ ( .D(csr_wdata_60_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[60]) );
  DFFX1_LVT csr_reg_dscratch_reg_60_ ( .D(csr_wdata_60_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[60]) );
  DFFSSRX1_LVT csr_reg_pmp_7_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_60_), .CLK(csr_net34743), .Q(io_ptw_pmp_7_cfg_a[1]), .QN(
        csr_n459) );
  DFFX1_LVT csr_u_T_49_reg_52_ ( .D(csr_N1943), .CLK(csr_n518), .Q(csr_n1941)
         );
  DFFX1_LVT csr_u_T_41_reg_52_ ( .D(csr_N1549), .CLK(csr_n576), .Q(
        csr_n_T_45_58_) );
  DFFX1_LVT csr_reg_sscratch_reg_58_ ( .D(csr_wdata_58_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[58]) );
  DFFX1_LVT csr_reg_mscratch_reg_58_ ( .D(csr_wdata_58_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[58]) );
  DFFX1_LVT csr_reg_dscratch_reg_58_ ( .D(csr_wdata_58_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[58]) );
  DFFX1_LVT csr_reg_pmp_7_cfg_x_reg ( .D(csr_wdata_58_), .CLK(csr_net34738), 
        .Q(io_ptw_pmp_7_cfg_x) );
  DFFX1_LVT csr_u_T_49_reg_51_ ( .D(csr_N1942), .CLK(csr_n519), .Q(csr_n1942)
         );
  DFFX1_LVT csr_u_T_41_reg_51_ ( .D(csr_N1548), .CLK(csr_n577), .Q(
        csr_n_T_45_57_) );
  DFFX1_LVT csr_reg_sscratch_reg_57_ ( .D(csr_wdata_57_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[57]) );
  DFFX1_LVT csr_reg_mscratch_reg_57_ ( .D(csr_wdata_57_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[57]) );
  DFFX1_LVT csr_reg_dscratch_reg_57_ ( .D(csr_wdata_57_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[57]) );
  DFFSSRX1_LVT csr_reg_pmp_7_cfg_w_reg ( .D(csr_wdata_56_), .SETB(1'b1), 
        .RSTB(csr_wdata_57_), .CLK(csr_net34738), .Q(io_ptw_pmp_7_cfg_w) );
  DFFX1_LVT csr_u_T_49_reg_50_ ( .D(csr_N1941), .CLK(csr_n519), .Q(csr_n1943)
         );
  DFFX1_LVT csr_u_T_41_reg_50_ ( .D(csr_N1547), .CLK(csr_n577), .Q(
        csr_n_T_45_56_) );
  DFFX1_LVT csr_reg_sscratch_reg_56_ ( .D(csr_wdata_56_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[56]) );
  DFFX1_LVT csr_reg_mscratch_reg_56_ ( .D(csr_wdata_56_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[56]) );
  DFFX1_LVT csr_reg_dscratch_reg_56_ ( .D(csr_wdata_56_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[56]) );
  DFFX1_LVT csr_reg_pmp_7_cfg_r_reg ( .D(csr_wdata_56_), .CLK(csr_net34738), 
        .Q(io_ptw_pmp_7_cfg_r) );
  DFFSSRX1_LVT csr_reg_pmp_7_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_63_), .CLK(csr_net34743), .Q(io_ptw_pmp_7_cfg_l), .QN(
        csr_n442) );
  DFFX1_LVT csr_reg_scause_reg_63_ ( .D(csr_N1333), .CLK(csr_n558), .Q(
        csr_reg_scause[63]) );
  DFFX1_LVT csr_reg_sscratch_reg_63_ ( .D(csr_wdata_63_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[63]) );
  DFFX1_LVT csr_reg_mscratch_reg_63_ ( .D(csr_wdata_63_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[63]) );
  DFFX1_LVT csr_reg_dscratch_reg_63_ ( .D(csr_wdata_63_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[63]) );
  DFFSSRX1_LVT csr_reg_mstatus_fs_reg_1_ ( .D(csr_wdata_13_), .SETB(csr_n51), 
        .RSTB(csr_n375), .CLK(csr_net35157), .Q(csr_n1928) );
  DFFX1_LVT csr_u_T_49_reg_7_ ( .D(csr_N1898), .CLK(csr_n519), .Q(
        csr_io_time[13]) );
  DFFX1_LVT csr_u_T_41_reg_7_ ( .D(csr_N1504), .CLK(csr_n577), .Q(
        csr_n_T_45_13_) );
  DFFSSRX1_LVT csr_reg_dcsr_ebreaks_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_13_), .CLK(csr_net35162), .Q(csr_n_T_1155_1_) );
  DFFX1_LVT csr_reg_stval_reg_13_ ( .D(csr_N1395), .CLK(csr_n560), .Q(
        csr_n_T_444[13]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_13_ ( .D(csr_n376), .SETB(csr_wdata_13_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_13_) );
  DFFX1_LVT csr_reg_mtval_reg_13_ ( .D(csr_N1006), .CLK(csr_n573), .Q(
        csr_n_T_383[13]) );
  DFFX1_LVT csr_reg_sscratch_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[13]) );
  DFFX1_LVT csr_reg_mscratch_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[13]) );
  DFFX1_LVT csr_reg_dscratch_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[13]) );
  DFFX1_LVT csr_reg_medeleg_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_net35172), 
        .Q(csr_read_medeleg_13) );
  DFFX1_LVT csr_reg_stvec_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_n569), .Q(
        csr_reg_stvec_13_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_13_ ( .D(csr_wdata_13_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[13]) );
  DFFX1_LVT csr_reg_dpc_reg_30_ ( .D(csr_net35214), .CLK(csr_n528), .Q(
        csr_reg_dpc_30_) );
  DFFX1_LVT csr_reg_mepc_reg_30_ ( .D(csr_net34992), .CLK(csr_n545), .Q(
        csr_reg_mepc_30_) );
  DFFX1_LVT csr_reg_sepc_reg_30_ ( .D(csr_net34790), .CLK(csr_n581), .Q(
        csr_reg_sepc_30_) );
  DFFX1_LVT csr_u_T_49_reg_24_ ( .D(csr_N1915), .CLK(csr_n519), .Q(
        csr_io_time[30]) );
  DFFX1_LVT csr_u_T_41_reg_24_ ( .D(csr_N1521), .CLK(csr_n577), .Q(
        csr_n_T_45_30_) );
  DFFX1_LVT csr_reg_stval_reg_30_ ( .D(csr_N1412), .CLK(csr_n560), .Q(
        csr_n_T_444[30]) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_30_ ( .D(csr_n376), .SETB(csr_wdata_30_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_30_) );
  DFFX1_LVT csr_reg_mtval_reg_30_ ( .D(csr_N1023), .CLK(csr_n573), .Q(
        csr_n_T_383[30]) );
  DFFX1_LVT csr_reg_sscratch_reg_30_ ( .D(csr_wdata_30_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[30]) );
  DFFX1_LVT csr_reg_mscratch_reg_30_ ( .D(csr_wdata_30_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[30]) );
  DFFX1_LVT csr_reg_dscratch_reg_30_ ( .D(csr_wdata_30_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[30]) );
  DFFX1_LVT csr_reg_stvec_reg_30_ ( .D(csr_wdata_30_), .CLK(csr_n569), .Q(
        csr_reg_stvec_30_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_30_ ( .D(csr_wdata_30_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[30]) );
  DFFX1_LVT csr_reg_dpc_reg_31_ ( .D(csr_net35211), .CLK(csr_n528), .Q(
        csr_reg_dpc_31_) );
  DFFX1_LVT csr_reg_mepc_reg_31_ ( .D(csr_net34989), .CLK(csr_n545), .Q(
        csr_reg_mepc_31_) );
  DFFX1_LVT csr_reg_sepc_reg_31_ ( .D(csr_net34787), .CLK(csr_n581), .Q(
        csr_reg_sepc_31_) );
  DFFX1_LVT csr_u_T_49_reg_25_ ( .D(csr_N1916), .CLK(csr_n519), .Q(
        csr_io_time[31]) );
  DFFX1_LVT csr_u_T_41_reg_25_ ( .D(csr_N1522), .CLK(csr_n577), .Q(
        csr_n_T_45_31_) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_2_ ( .D(csr_n_GEN_279[2]), .CLK(csr_n536), 
        .Q(io_ptw_pmp_3_addr[2]) );
  DFFX1_LVT csr_reg_pmp_3_addr_reg_0_ ( .D(csr_n_GEN_279[0]), .CLK(csr_n537), 
        .Q(io_ptw_pmp_3_addr[0]) );
  DFFSSRX1_LVT csr_reg_pmp_3_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_31_), .CLK(csr_net35127), .Q(io_ptw_pmp_3_cfg_l), .QN(
        csr_n443) );
  DFFX1_LVT csr_reg_stval_reg_31_ ( .D(csr_N1413), .CLK(csr_n560), .Q(
        csr_n_T_444[31]) );
  DFFX1_LVT csr_reg_mtval_reg_31_ ( .D(csr_N1024), .CLK(csr_n573), .Q(
        csr_n_T_383[31]) );
  DFFX1_LVT csr_reg_sscratch_reg_31_ ( .D(csr_wdata_31_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[31]) );
  DFFX1_LVT csr_reg_mscratch_reg_31_ ( .D(csr_wdata_31_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[31]) );
  DFFX1_LVT csr_reg_dscratch_reg_31_ ( .D(csr_wdata_31_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[31]) );
  DFFX1_LVT csr_reg_stvec_reg_31_ ( .D(csr_wdata_31_), .CLK(csr_n569), .Q(
        csr_reg_stvec_31_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_31_ ( .D(csr_wdata_31_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[31]) );
  DFFX1_LVT csr_reg_dpc_reg_32_ ( .D(csr_net35208), .CLK(csr_n528), .Q(
        csr_reg_dpc_32_) );
  DFFX1_LVT csr_reg_mepc_reg_32_ ( .D(csr_net34986), .CLK(csr_n545), .Q(
        csr_reg_mepc_32_) );
  DFFX1_LVT csr_reg_sepc_reg_32_ ( .D(csr_net34784), .CLK(csr_n581), .Q(
        csr_reg_sepc_32_) );
  DFFX1_LVT csr_reg_dpc_reg_33_ ( .D(csr_net35205), .CLK(csr_n528), .Q(
        csr_reg_dpc_33_) );
  DFFX1_LVT csr_reg_mepc_reg_33_ ( .D(csr_net34983), .CLK(csr_n545), .Q(
        csr_reg_mepc_33_) );
  DFFX1_LVT csr_reg_sepc_reg_33_ ( .D(csr_net34781), .CLK(csr_n581), .Q(
        csr_reg_sepc_33_) );
  DFFX1_LVT csr_u_T_49_reg_27_ ( .D(csr_N1918), .CLK(csr_n519), .Q(csr_n1966)
         );
  DFFX1_LVT csr_u_T_41_reg_27_ ( .D(csr_N1524), .CLK(csr_n577), .Q(
        csr_n_T_45_33_) );
  DFFX1_LVT csr_reg_stval_reg_33_ ( .D(csr_N1415), .CLK(csr_n560), .Q(
        csr_n_T_444[33]) );
  DFFX1_LVT csr_reg_mtval_reg_33_ ( .D(csr_N1026), .CLK(csr_n573), .Q(
        csr_n_T_383[33]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_33_ ( .D(csr_wdata_33_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[33]) );
  DFFX1_LVT csr_reg_sscratch_reg_33_ ( .D(csr_wdata_33_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[33]) );
  DFFX1_LVT csr_reg_mscratch_reg_33_ ( .D(csr_wdata_33_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[33]) );
  DFFX1_LVT csr_reg_dscratch_reg_33_ ( .D(csr_wdata_33_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[33]) );
  DFFX1_LVT csr_reg_stvec_reg_33_ ( .D(csr_wdata_33_), .CLK(csr_n569), .Q(
        csr_reg_stvec_33_) );
  DFFSSRX1_LVT csr_reg_pmp_4_cfg_w_reg ( .D(csr_wdata_32_), .SETB(1'b1), 
        .RSTB(csr_wdata_33_), .CLK(csr_net35117), .Q(io_ptw_pmp_4_cfg_w) );
  DFFX1_LVT csr_u_T_49_reg_26_ ( .D(csr_N1917), .CLK(csr_n519), .Q(csr_n1967)
         );
  DFFX1_LVT csr_u_T_41_reg_26_ ( .D(csr_N1523), .CLK(csr_n577), .Q(
        csr_n_T_45_32_) );
  DFFX1_LVT csr_reg_stval_reg_32_ ( .D(csr_N1414), .CLK(csr_n559), .Q(
        csr_n_T_444[32]) );
  DFFX1_LVT csr_reg_mtval_reg_32_ ( .D(csr_N1025), .CLK(csr_n572), .Q(
        csr_n_T_383[32]) );
  DFFX1_LVT csr_reg_sscratch_reg_32_ ( .D(csr_wdata_32_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[32]) );
  DFFX1_LVT csr_reg_mscratch_reg_32_ ( .D(csr_wdata_32_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[32]) );
  DFFX1_LVT csr_reg_pmp_4_cfg_r_reg ( .D(csr_wdata_32_), .CLK(csr_net35117), 
        .Q(io_ptw_pmp_4_cfg_r) );
  DFFX1_LVT csr_reg_dscratch_reg_32_ ( .D(csr_wdata_32_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[32]) );
  DFFX1_LVT csr_reg_stvec_reg_32_ ( .D(csr_wdata_32_), .CLK(csr_n568), .Q(
        csr_reg_stvec_32_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_32_ ( .D(csr_wdata_32_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[32]) );
  DFFX1_LVT csr_reg_dpc_reg_34_ ( .D(csr_net35202), .CLK(csr_n528), .Q(
        csr_reg_dpc_34_) );
  DFFX1_LVT csr_reg_mepc_reg_34_ ( .D(csr_net34980), .CLK(csr_n545), .Q(
        csr_reg_mepc_34_) );
  DFFX1_LVT csr_reg_sepc_reg_34_ ( .D(csr_net34778), .CLK(csr_n581), .Q(
        csr_reg_sepc_34_) );
  DFFX1_LVT csr_u_T_49_reg_28_ ( .D(csr_N1919), .CLK(csr_n519), .Q(csr_n1965)
         );
  DFFX1_LVT csr_u_T_41_reg_28_ ( .D(csr_N1525), .CLK(csr_n577), .Q(
        csr_n_T_45_34_) );
  DFFX1_LVT csr_reg_stval_reg_34_ ( .D(csr_N1416), .CLK(csr_n559), .Q(
        csr_n_T_444[34]) );
  DFFX1_LVT csr_reg_mtval_reg_34_ ( .D(csr_N1027), .CLK(csr_n572), .Q(
        csr_n_T_383[34]) );
  DFFX1_LVT csr_reg_sscratch_reg_34_ ( .D(csr_wdata_34_), .CLK(csr_n564), .Q(
        csr_reg_sscratch[34]) );
  DFFX1_LVT csr_reg_mscratch_reg_34_ ( .D(csr_wdata_34_), .CLK(csr_n550), .Q(
        csr_reg_mscratch[34]) );
  DFFX1_LVT csr_reg_pmp_4_cfg_x_reg ( .D(csr_wdata_34_), .CLK(csr_net35117), 
        .Q(io_ptw_pmp_4_cfg_x) );
  DFFX1_LVT csr_reg_dscratch_reg_34_ ( .D(csr_wdata_34_), .CLK(csr_n524), .Q(
        csr_reg_dscratch[34]) );
  DFFX1_LVT csr_reg_stvec_reg_34_ ( .D(csr_wdata_34_), .CLK(csr_n568), .Q(
        csr_reg_stvec_34_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_34_ ( .D(csr_wdata_34_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[34]) );
  DFFX1_LVT csr_reg_dpc_reg_35_ ( .D(csr_net35199), .CLK(csr_n528), .Q(
        csr_reg_dpc_35_) );
  DFFX1_LVT csr_reg_mepc_reg_35_ ( .D(csr_net34977), .CLK(csr_n545), .Q(
        csr_reg_mepc_35_) );
  DFFX1_LVT csr_reg_sepc_reg_35_ ( .D(csr_net34775), .CLK(csr_n581), .Q(
        csr_reg_sepc_35_) );
  DFFX1_LVT csr_u_T_49_reg_29_ ( .D(csr_N1920), .CLK(csr_n519), .Q(csr_n1964)
         );
  DFFX1_LVT csr_u_T_41_reg_29_ ( .D(csr_N1526), .CLK(csr_n577), .Q(
        csr_n_T_45_35_) );
  DFFSSRX1_LVT csr_reg_pmp_4_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_35_), .CLK(csr_net34910), .Q(io_ptw_pmp_4_cfg_a[0]) );
  DFFX1_LVT csr_reg_stval_reg_35_ ( .D(csr_N1417), .CLK(csr_n559), .Q(
        csr_n_T_444[35]) );
  DFFX1_LVT csr_reg_mtval_reg_35_ ( .D(csr_N1028), .CLK(csr_n572), .Q(
        csr_n_T_383[35]) );
  DFFX1_LVT csr_reg_sscratch_reg_35_ ( .D(csr_wdata_35_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[35]) );
  DFFX1_LVT csr_reg_mscratch_reg_35_ ( .D(csr_wdata_35_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[35]) );
  DFFX1_LVT csr_reg_dscratch_reg_35_ ( .D(csr_wdata_35_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[35]) );
  DFFX1_LVT csr_reg_stvec_reg_35_ ( .D(csr_wdata_35_), .CLK(csr_n568), .Q(
        csr_reg_stvec_35_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_35_ ( .D(csr_wdata_35_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[35]) );
  DFFX1_LVT csr_reg_dpc_reg_36_ ( .D(csr_net35196), .CLK(csr_n528), .Q(
        csr_reg_dpc_36_) );
  DFFX1_LVT csr_reg_mepc_reg_36_ ( .D(csr_net34974), .CLK(csr_n545), .Q(
        csr_reg_mepc_36_) );
  DFFX1_LVT csr_reg_sepc_reg_36_ ( .D(csr_net34772), .CLK(csr_n581), .Q(
        csr_reg_sepc_36_) );
  DFFX1_LVT csr_u_T_49_reg_30_ ( .D(csr_N1921), .CLK(csr_n519), .Q(csr_n1963)
         );
  DFFX1_LVT csr_u_T_41_reg_30_ ( .D(csr_N1527), .CLK(csr_n577), .Q(
        csr_n_T_45_36_) );
  DFFSSRX1_LVT csr_reg_pmp_4_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_36_), .CLK(csr_net34910), .Q(io_ptw_pmp_4_cfg_a[1]), .QN(
        csr_n464) );
  DFFX1_LVT csr_reg_stval_reg_36_ ( .D(csr_N1418), .CLK(csr_n559), .Q(
        csr_n_T_444[36]) );
  DFFX1_LVT csr_reg_mtval_reg_36_ ( .D(csr_N1029), .CLK(csr_n572), .Q(
        csr_n_T_383[36]) );
  DFFX1_LVT csr_reg_sscratch_reg_36_ ( .D(csr_wdata_36_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[36]) );
  DFFX1_LVT csr_reg_mscratch_reg_36_ ( .D(csr_wdata_36_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[36]) );
  DFFX1_LVT csr_reg_dscratch_reg_36_ ( .D(csr_wdata_36_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[36]) );
  DFFX1_LVT csr_reg_stvec_reg_36_ ( .D(csr_wdata_36_), .CLK(csr_n568), .Q(
        csr_reg_stvec_36_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_36_ ( .D(csr_wdata_36_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[36]) );
  DFFX1_LVT csr_reg_dpc_reg_37_ ( .D(csr_net35193), .CLK(csr_n528), .Q(
        csr_reg_dpc_37_) );
  DFFX1_LVT csr_reg_mepc_reg_37_ ( .D(csr_net34971), .CLK(csr_n545), .Q(
        csr_reg_mepc_37_) );
  DFFX1_LVT csr_reg_sepc_reg_37_ ( .D(csr_net34769), .CLK(csr_n581), .Q(
        csr_reg_sepc_37_) );
  DFFX1_LVT csr_u_T_49_reg_31_ ( .D(csr_N1922), .CLK(csr_n519), .Q(csr_n1962)
         );
  DFFX1_LVT csr_u_T_41_reg_31_ ( .D(csr_N1528), .CLK(csr_n577), .Q(
        csr_n_T_45_37_) );
  DFFX1_LVT csr_reg_stval_reg_37_ ( .D(csr_N1419), .CLK(csr_n559), .Q(
        csr_n_T_444[37]) );
  DFFX1_LVT csr_reg_mtval_reg_37_ ( .D(csr_N1030), .CLK(csr_n572), .Q(
        csr_n_T_383[37]) );
  DFFX1_LVT csr_reg_sscratch_reg_37_ ( .D(csr_wdata_37_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[37]) );
  DFFX1_LVT csr_reg_mscratch_reg_37_ ( .D(csr_wdata_37_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[37]) );
  DFFX1_LVT csr_reg_dscratch_reg_37_ ( .D(csr_wdata_37_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[37]) );
  DFFX1_LVT csr_reg_stvec_reg_37_ ( .D(csr_wdata_37_), .CLK(csr_n568), .Q(
        csr_reg_stvec_37_) );
  DFFX1_LVT csr_reg_bp_0_address_reg_37_ ( .D(csr_wdata_37_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[37]) );
  DFFX1_LVT csr_reg_dpc_reg_38_ ( .D(csr_net35190), .CLK(csr_n528), .Q(
        csr_reg_dpc_38_) );
  DFFX1_LVT csr_reg_mepc_reg_38_ ( .D(csr_net34968), .CLK(csr_n545), .Q(
        csr_reg_mepc_38_) );
  DFFX1_LVT csr_reg_sepc_reg_38_ ( .D(csr_net34766), .CLK(csr_n581), .Q(
        csr_reg_sepc_38_) );
  DFFX1_LVT csr_u_T_49_reg_32_ ( .D(csr_N1923), .CLK(csr_n519), .Q(csr_n1961)
         );
  DFFX1_LVT csr_u_T_41_reg_32_ ( .D(csr_N1529), .CLK(csr_n577), .Q(
        csr_n_T_45_38_) );
  DFFX1_LVT csr_reg_stval_reg_38_ ( .D(csr_N1420), .CLK(csr_n559), .Q(
        csr_n_T_444[38]) );
  DFFX1_LVT csr_reg_mtval_reg_38_ ( .D(csr_N1031), .CLK(csr_n572), .Q(
        csr_n_T_383[38]) );
  DFFX1_LVT csr_reg_sscratch_reg_38_ ( .D(csr_wdata_38_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[38]) );
  DFFX1_LVT csr_reg_mscratch_reg_38_ ( .D(csr_wdata_38_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[38]) );
  DFFX1_LVT csr_reg_dscratch_reg_38_ ( .D(csr_wdata_38_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[38]) );
  DFFX1_LVT csr_reg_stvec_reg_38_ ( .D(csr_wdata_38_), .CLK(csr_n568), .Q(
        csr_reg_stvec_38_), .QN(csr_n465) );
  DFFX1_LVT csr_u_T_49_reg_49_ ( .D(csr_N1940), .CLK(csr_n520), .Q(csr_n1944)
         );
  DFFX1_LVT csr_u_T_41_reg_49_ ( .D(csr_N1546), .CLK(csr_n578), .Q(
        csr_n_T_45_55_) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_2_ ( .D(csr_n_GEN_293[2]), .CLK(csr_n539), 
        .Q(io_ptw_pmp_5_addr[2]) );
  DFFX1_LVT csr_reg_pmp_5_addr_reg_0_ ( .D(csr_n_GEN_293[0]), .CLK(csr_n540), 
        .Q(io_ptw_pmp_5_addr[0]) );
  DFFX1_LVT csr_u_T_49_reg_45_ ( .D(csr_N1936), .CLK(csr_n520), .Q(csr_n1948)
         );
  DFFX1_LVT csr_u_T_41_reg_45_ ( .D(csr_N1542), .CLK(csr_n578), .Q(
        csr_n_T_45_51_) );
  DFFX1_LVT csr_reg_sscratch_reg_51_ ( .D(csr_wdata_51_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[51]) );
  DFFX1_LVT csr_reg_mscratch_reg_51_ ( .D(csr_wdata_51_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[51]) );
  DFFX1_LVT csr_reg_dscratch_reg_51_ ( .D(csr_wdata_51_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[51]) );
  DFFSSRX1_LVT csr_reg_pmp_6_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_51_), .CLK(csr_net35102), .Q(io_ptw_pmp_6_cfg_a[0]) );
  DFFX1_LVT csr_u_T_49_reg_46_ ( .D(csr_N1937), .CLK(csr_n520), .Q(csr_n1947)
         );
  DFFX1_LVT csr_u_T_41_reg_46_ ( .D(csr_N1543), .CLK(csr_n578), .Q(
        csr_n_T_45_52_) );
  DFFX1_LVT csr_reg_sscratch_reg_52_ ( .D(csr_wdata_52_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[52]) );
  DFFX1_LVT csr_reg_mscratch_reg_52_ ( .D(csr_wdata_52_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[52]) );
  DFFX1_LVT csr_reg_dscratch_reg_52_ ( .D(csr_wdata_52_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[52]) );
  DFFSSRX1_LVT csr_reg_pmp_6_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_52_), .CLK(csr_net35102), .Q(io_ptw_pmp_6_cfg_a[1]), .QN(
        csr_n458) );
  DFFX1_LVT csr_u_T_49_reg_44_ ( .D(csr_N1935), .CLK(csr_n520), .Q(csr_n1949)
         );
  DFFX1_LVT csr_u_T_41_reg_44_ ( .D(csr_N1541), .CLK(csr_n578), .Q(
        csr_n_T_45_50_) );
  DFFX1_LVT csr_reg_sscratch_reg_50_ ( .D(csr_wdata_50_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[50]) );
  DFFX1_LVT csr_reg_mscratch_reg_50_ ( .D(csr_wdata_50_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[50]) );
  DFFX1_LVT csr_reg_dscratch_reg_50_ ( .D(csr_wdata_50_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[50]) );
  DFFX1_LVT csr_reg_pmp_6_cfg_x_reg ( .D(csr_wdata_50_), .CLK(csr_net35107), 
        .Q(io_ptw_pmp_6_cfg_x) );
  DFFX1_LVT csr_u_T_49_reg_43_ ( .D(csr_N1934), .CLK(csr_n520), .Q(csr_n1950)
         );
  DFFX1_LVT csr_u_T_41_reg_43_ ( .D(csr_N1540), .CLK(csr_n578), .Q(
        csr_n_T_45_49_) );
  DFFX1_LVT csr_reg_sscratch_reg_49_ ( .D(csr_wdata_49_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[49]) );
  DFFX1_LVT csr_reg_mscratch_reg_49_ ( .D(csr_wdata_49_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[49]) );
  DFFX1_LVT csr_reg_dscratch_reg_49_ ( .D(csr_wdata_49_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[49]) );
  DFFX1_LVT csr_u_T_49_reg_42_ ( .D(csr_N1933), .CLK(csr_n520), .Q(csr_n1951)
         );
  DFFX1_LVT csr_u_T_41_reg_42_ ( .D(csr_N1539), .CLK(csr_n578), .Q(
        csr_n_T_45_48_) );
  DFFX1_LVT csr_reg_sscratch_reg_48_ ( .D(csr_wdata_48_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[48]) );
  DFFX1_LVT csr_reg_mscratch_reg_48_ ( .D(csr_wdata_48_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[48]) );
  DFFX1_LVT csr_reg_dscratch_reg_48_ ( .D(csr_wdata_48_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[48]) );
  DFFX1_LVT csr_reg_pmp_6_cfg_r_reg ( .D(csr_wdata_48_), .CLK(csr_net35107), 
        .Q(io_ptw_pmp_6_cfg_r) );
  DFFX1_LVT csr_reg_sscratch_reg_55_ ( .D(csr_wdata_55_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[55]) );
  DFFX1_LVT csr_reg_mscratch_reg_55_ ( .D(csr_wdata_55_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[55]) );
  DFFX1_LVT csr_reg_dscratch_reg_55_ ( .D(csr_wdata_55_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[55]) );
  DFFX1_LVT csr_u_T_49_reg_55_ ( .D(csr_N1946), .CLK(csr_n520), .Q(csr_n1938)
         );
  DFFX1_LVT csr_u_T_41_reg_55_ ( .D(csr_N1552), .CLK(csr_n578), .Q(
        csr_n_T_45_61_) );
  DFFX1_LVT csr_reg_sscratch_reg_61_ ( .D(csr_wdata_61_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[61]) );
  DFFX1_LVT csr_reg_mscratch_reg_61_ ( .D(csr_wdata_61_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[61]) );
  DFFX1_LVT csr_reg_dscratch_reg_61_ ( .D(csr_wdata_61_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[61]) );
  DFFX1_LVT csr_reg_dpc_reg_39_ ( .D(csr_net35187), .CLK(csr_n528), .Q(
        csr_reg_dpc_39_) );
  DFFX1_LVT csr_reg_mepc_reg_39_ ( .D(csr_net34965), .CLK(csr_n545), .Q(
        csr_reg_mepc_39_) );
  DFFX1_LVT csr_reg_sepc_reg_39_ ( .D(csr_net34763), .CLK(csr_n581), .Q(
        csr_reg_sepc_39_) );
  DFFX1_LVT csr_u_T_49_reg_33_ ( .D(csr_N1924), .CLK(csr_n520), .Q(csr_n1960)
         );
  DFFX1_LVT csr_u_T_41_reg_33_ ( .D(csr_N1530), .CLK(csr_n578), .Q(
        csr_n_T_45_39_) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_2_ ( .D(csr_n_GEN_286[2]), .CLK(csr_n538), 
        .Q(io_ptw_pmp_4_addr[2]) );
  DFFX1_LVT csr_reg_pmp_4_addr_reg_0_ ( .D(csr_n_GEN_286[0]), .CLK(csr_n532), 
        .Q(io_ptw_pmp_4_addr[0]) );
  DFFSSRX1_LVT csr_reg_pmp_4_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_39_), .CLK(csr_net34910), .Q(io_ptw_pmp_4_cfg_l), .QN(
        csr_n438) );
  DFFX1_LVT csr_reg_stval_reg_39_ ( .D(csr_N1421), .CLK(csr_n559), .Q(
        csr_n_T_444[39]) );
  DFFX1_LVT csr_reg_mtval_reg_39_ ( .D(csr_N1032), .CLK(csr_n572), .Q(
        csr_n_T_383[39]) );
  DFFX1_LVT csr_reg_sscratch_reg_39_ ( .D(csr_wdata_39_), .CLK(csr_n565), .Q(
        csr_reg_sscratch[39]) );
  DFFX1_LVT csr_reg_mscratch_reg_39_ ( .D(csr_wdata_39_), .CLK(csr_n551), .Q(
        csr_reg_mscratch[39]) );
  DFFX1_LVT csr_reg_dscratch_reg_39_ ( .D(csr_wdata_39_), .CLK(csr_n525), .Q(
        csr_reg_dscratch[39]) );
  DFFX1_LVT csr_u_T_49_reg_56_ ( .D(csr_N1947), .CLK(csr_n520), .Q(csr_n1937)
         );
  DFFX1_LVT csr_u_T_41_reg_56_ ( .D(csr_N1553), .CLK(csr_n578), .Q(
        csr_n_T_45_62_) );
  DFFX1_LVT csr_reg_sscratch_reg_62_ ( .D(csr_wdata_62_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[62]) );
  DFFX1_LVT csr_reg_mscratch_reg_62_ ( .D(csr_wdata_62_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[62]) );
  DFFX1_LVT csr_reg_dscratch_reg_62_ ( .D(csr_wdata_62_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[62]) );
  DFFX1_LVT csr_u_T_49_reg_35_ ( .D(csr_N1926), .CLK(csr_n520), .Q(csr_n1958)
         );
  DFFX1_LVT csr_u_T_41_reg_35_ ( .D(csr_N1532), .CLK(csr_n578), .Q(
        csr_n_T_45_41_) );
  DFFX1_LVT csr_reg_sscratch_reg_41_ ( .D(csr_wdata_41_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[41]) );
  DFFX1_LVT csr_reg_mscratch_reg_41_ ( .D(csr_wdata_41_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[41]) );
  DFFX1_LVT csr_reg_dscratch_reg_41_ ( .D(csr_wdata_41_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[41]) );
  DFFSSRX1_LVT csr_reg_pmp_5_cfg_w_reg ( .D(csr_wdata_40_), .SETB(1'b1), 
        .RSTB(csr_wdata_41_), .CLK(csr_net35097), .Q(io_ptw_pmp_5_cfg_w) );
  DFFX1_LVT csr_u_T_49_reg_34_ ( .D(csr_N1925), .CLK(csr_n520), .Q(csr_n1959)
         );
  DFFX1_LVT csr_u_T_41_reg_34_ ( .D(csr_N1531), .CLK(csr_n578), .Q(
        csr_n_T_45_40_) );
  DFFX1_LVT csr_reg_sscratch_reg_40_ ( .D(csr_wdata_40_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[40]) );
  DFFX1_LVT csr_reg_mscratch_reg_40_ ( .D(csr_wdata_40_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[40]) );
  DFFX1_LVT csr_reg_pmp_5_cfg_r_reg ( .D(csr_wdata_40_), .CLK(csr_net35097), 
        .Q(io_ptw_pmp_5_cfg_r) );
  DFFX1_LVT csr_reg_dscratch_reg_40_ ( .D(csr_wdata_40_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[40]) );
  DFFX1_LVT csr_u_T_49_reg_36_ ( .D(csr_N1927), .CLK(csr_n520), .Q(csr_n1957)
         );
  DFFX1_LVT csr_u_T_41_reg_36_ ( .D(csr_N1533), .CLK(csr_n578), .Q(
        csr_n_T_45_42_) );
  DFFX1_LVT csr_reg_sscratch_reg_42_ ( .D(csr_wdata_42_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[42]) );
  DFFX1_LVT csr_reg_mscratch_reg_42_ ( .D(csr_wdata_42_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[42]) );
  DFFX1_LVT csr_reg_pmp_5_cfg_x_reg ( .D(csr_wdata_42_), .CLK(csr_net35097), 
        .Q(io_ptw_pmp_5_cfg_x) );
  DFFX1_LVT csr_reg_dscratch_reg_42_ ( .D(csr_wdata_42_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[42]) );
  DFFX1_LVT csr_u_T_49_reg_37_ ( .D(csr_N1928), .CLK(csr_n521), .Q(csr_n1956)
         );
  DFFX1_LVT csr_u_T_41_reg_37_ ( .D(csr_N1534), .CLK(csr_n579), .Q(
        csr_n_T_45_43_) );
  DFFSSRX1_LVT csr_reg_pmp_5_cfg_a_reg_0_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_43_), .CLK(csr_net35112), .Q(io_ptw_pmp_5_cfg_a[0]) );
  DFFX1_LVT csr_reg_sscratch_reg_43_ ( .D(csr_wdata_43_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[43]) );
  DFFX1_LVT csr_reg_mscratch_reg_43_ ( .D(csr_wdata_43_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[43]) );
  DFFX1_LVT csr_reg_dscratch_reg_43_ ( .D(csr_wdata_43_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[43]) );
  DFFX1_LVT csr_u_T_49_reg_38_ ( .D(csr_N1929), .CLK(csr_n521), .Q(csr_n1955)
         );
  DFFX1_LVT csr_u_T_41_reg_38_ ( .D(csr_N1535), .CLK(csr_n579), .Q(
        csr_n_T_45_44_) );
  DFFSSRX1_LVT csr_reg_pmp_5_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_44_), .CLK(csr_net35112), .Q(io_ptw_pmp_5_cfg_a[1]), .QN(
        csr_n461) );
  DFFX1_LVT csr_reg_sscratch_reg_44_ ( .D(csr_wdata_44_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[44]) );
  DFFX1_LVT csr_reg_mscratch_reg_44_ ( .D(csr_wdata_44_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[44]) );
  DFFX1_LVT csr_reg_dscratch_reg_44_ ( .D(csr_wdata_44_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[44]) );
  DFFX1_LVT csr_u_T_49_reg_39_ ( .D(csr_N1930), .CLK(csr_n521), .Q(csr_n1954)
         );
  DFFX1_LVT csr_u_T_41_reg_39_ ( .D(csr_N1536), .CLK(csr_n579), .Q(
        csr_n_T_45_45_) );
  DFFX1_LVT csr_reg_sscratch_reg_45_ ( .D(csr_wdata_45_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[45]) );
  DFFX1_LVT csr_reg_mscratch_reg_45_ ( .D(csr_wdata_45_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[45]) );
  DFFX1_LVT csr_reg_dscratch_reg_45_ ( .D(csr_wdata_45_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[45]) );
  DFFX1_LVT csr_u_T_49_reg_40_ ( .D(csr_N1931), .CLK(csr_n521), .Q(csr_n1953)
         );
  DFFX1_LVT csr_u_T_41_reg_40_ ( .D(csr_N1537), .CLK(csr_n579), .Q(
        csr_n_T_45_46_) );
  DFFX1_LVT csr_reg_sscratch_reg_46_ ( .D(csr_wdata_46_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[46]) );
  DFFX1_LVT csr_reg_mscratch_reg_46_ ( .D(csr_wdata_46_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[46]) );
  DFFX1_LVT csr_reg_dscratch_reg_46_ ( .D(csr_wdata_46_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[46]) );
  DFFX1_LVT csr_u_T_49_reg_41_ ( .D(csr_N1932), .CLK(csr_n521), .Q(csr_n1952)
         );
  DFFX1_LVT csr_u_T_41_reg_41_ ( .D(csr_N1538), .CLK(csr_n579), .Q(
        csr_n_T_45_47_) );
  DFFSSRX1_LVT csr_reg_pmp_5_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_47_), .CLK(csr_net35112), .Q(io_ptw_pmp_5_cfg_l), .QN(
        csr_n437) );
  DFFX1_LVT csr_reg_sscratch_reg_47_ ( .D(csr_wdata_47_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[47]) );
  DFFX1_LVT csr_reg_mscratch_reg_47_ ( .D(csr_wdata_47_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[47]) );
  DFFX1_LVT csr_reg_dscratch_reg_47_ ( .D(csr_wdata_47_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[47]) );
  DFFX1_LVT csr_u_T_49_reg_47_ ( .D(csr_N1938), .CLK(csr_n521), .Q(csr_n1946)
         );
  DFFX1_LVT csr_u_T_41_reg_47_ ( .D(csr_N1544), .CLK(csr_n579), .Q(
        csr_n_T_45_53_) );
  DFFX1_LVT csr_reg_sscratch_reg_53_ ( .D(csr_wdata_53_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[53]) );
  DFFX1_LVT csr_reg_mscratch_reg_53_ ( .D(csr_wdata_53_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[53]) );
  DFFX1_LVT csr_reg_dscratch_reg_53_ ( .D(csr_wdata_53_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[53]) );
  DFFX1_LVT csr_u_T_49_reg_48_ ( .D(csr_N1939), .CLK(csr_n521), .Q(csr_n1945)
         );
  DFFX1_LVT csr_reg_sscratch_reg_54_ ( .D(csr_wdata_54_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[54]) );
  DFFX1_LVT csr_reg_mscratch_reg_54_ ( .D(csr_wdata_54_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[54]) );
  DFFX1_LVT csr_reg_dscratch_reg_54_ ( .D(csr_wdata_54_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[54]) );
  DFFX1_LVT csr_reg_bp_0_address_reg_38_ ( .D(csr_wdata_38_), .CLK(csr_n584), 
        .Q(csr_io_bp_0_address[38]) );
  DFFSSRX1_LVT csr_reg_bp_0_control_r_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_0_), .CLK(csr_net35314), .Q(csr_io_bp_0_control_r) );
  DFFSSRX1_LVT csr_reg_bp_0_control_x_reg ( .D(csr_n503), .SETB(1'b1), .RSTB(
        csr_wdata_2_), .CLK(csr_net35314), .Q(csr_io_bp_0_control_x) );
  DFFX1_LVT csr_reg_bp_0_control_action_reg ( .D(csr_N485), .CLK(csr_net35314), 
        .Q(csr_io_bp_0_control_action) );
  DFFX1_LVT csr_reg_bp_0_control_dmode_reg ( .D(csr_n1482), .CLK(csr_net35314), 
        .Q(csr_n_T_366_59_), .QN(csr_n457) );
  DFFX1_LVT csr_reg_bp_0_control_tmatch_reg_0_ ( .D(csr_wdata_7_), .CLK(
        csr_net35319), .Q(csr_io_bp_0_control_tmatch[0]) );
  DFFX1_LVT csr_reg_bp_0_control_tmatch_reg_1_ ( .D(csr_wdata_8_), .CLK(
        csr_net35319), .Q(csr_io_bp_0_control_tmatch[1]) );
  DFFX1_LVT csr_reg_dcsr_cause_reg_1_ ( .D(csr_N469), .CLK(csr_net35177), .Q(
        csr_n_T_389[7]) );
  DFFX1_LVT csr_reg_dpc_reg_2_ ( .D(csr_net35298), .CLK(csr_n528), .Q(
        csr_reg_dpc_2_) );
  DFFX1_LVT csr_reg_singleStepped_reg ( .D(csr_N435), .CLK(csr_n594), .Q(
        csr_n426), .QN(csr_n860) );
  DFFX1_LVT csr_reg_debug_reg ( .D(csr_n2161), .CLK(csr_n594), .Q(
        csr_io_status_debug), .QN(n9516) );
  DFFX1_LVT csr_reg_sepc_reg_2_ ( .D(csr_net34874), .CLK(csr_n581), .Q(
        csr_reg_sepc_2_) );
  DFFX1_LVT csr_reg_mepc_reg_2_ ( .D(csr_net35076), .CLK(csr_n545), .Q(
        csr_reg_mepc_2_) );
  DFFX1_LVT csr_reg_mcause_reg_0_ ( .D(csr_N881), .CLK(csr_n580), .Q(
        csr_reg_mcause[0]) );
  DFFX1_LVT csr_reg_mcause_reg_2_ ( .D(csr_N883), .CLK(csr_net34885), .Q(
        csr_reg_mcause[2]) );
  DFFX1_LVT csr_reg_mtval_reg_0_ ( .D(csr_N993), .CLK(csr_n572), .Q(
        csr_n_T_383[0]) );
  DFFX1_LVT csr_reg_mtval_reg_2_ ( .D(csr_N995), .CLK(csr_n572), .Q(
        csr_n_T_383[2]) );
  DFFX1_LVT csr_reg_mtval_reg_7_ ( .D(csr_N1000), .CLK(csr_n572), .Q(
        csr_n_T_383[7]) );
  DFFX1_LVT csr_reg_mtval_reg_8_ ( .D(csr_N1001), .CLK(csr_n572), .Q(
        csr_n_T_383[8]) );
  DFFX1_LVT csr_reg_mtval_reg_12_ ( .D(csr_N1005), .CLK(csr_n572), .Q(
        csr_n_T_383[12]) );
  DFFX1_LVT csr_reg_stval_reg_0_ ( .D(csr_N1382), .CLK(csr_n559), .Q(
        csr_n_T_444[0]) );
  DFFX1_LVT csr_reg_stval_reg_2_ ( .D(csr_N1384), .CLK(csr_n559), .Q(
        csr_n_T_444[2]) );
  DFFX1_LVT csr_reg_stval_reg_7_ ( .D(csr_N1389), .CLK(csr_n559), .Q(
        csr_n_T_444[7]) );
  DFFX1_LVT csr_reg_stval_reg_8_ ( .D(csr_N1390), .CLK(csr_n559), .Q(
        csr_n_T_444[8]) );
  DFFX1_LVT csr_reg_stval_reg_12_ ( .D(csr_N1394), .CLK(csr_n559), .Q(
        csr_n_T_444[12]) );
  DFFX1_LVT csr_reg_scause_reg_0_ ( .D(csr_N1270), .CLK(csr_n557), .Q(
        csr_reg_scause[0]) );
  DFFX1_LVT csr_reg_scause_reg_2_ ( .D(csr_N1272), .CLK(csr_n557), .Q(
        csr_reg_scause[2]) );
  DFFX1_LVT csr_reg_mstatus_spp_reg ( .D(csr_n1913), .CLK(csr_n1915), .Q(
        csr_n1931) );
  DFFX1_LVT csr_u_T_49_reg_2_ ( .D(csr_N1893), .CLK(csr_n521), .Q(
        csr_io_time[8]) );
  DFFX1_LVT csr_u_T_41_reg_2_ ( .D(csr_N1499), .CLK(csr_n579), .Q(
        csr_n_T_45_8_) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_8_ ( .D(csr_n376), .SETB(csr_wdata_8_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_8_) );
  DFFX1_LVT csr_reg_sscratch_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_n566), .Q(
        csr_reg_sscratch[8]) );
  DFFX1_LVT csr_reg_mscratch_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_n552), .Q(
        csr_reg_mscratch[8]) );
  DFFX1_LVT csr_reg_dscratch_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_n526), .Q(
        csr_reg_dscratch[8]) );
  DFFX1_LVT csr_reg_medeleg_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_net35172), .Q(
        csr_read_medeleg_8) );
  DFFX1_LVT csr_reg_stvec_reg_8_ ( .D(csr_wdata_8_), .CLK(csr_n568), .Q(
        csr_reg_stvec_8_) );
  DFFX1_LVT csr_reg_misa_reg_8_ ( .D(csr_N1567), .CLK(csr_net35137), .Q(
        csr_n1922) );
  DFFX1_LVT csr_reg_misa_reg_18_ ( .D(csr_N1577), .CLK(csr_net35137), .Q(
        csr_n1921) );
  DFFX1_LVT csr_reg_misa_reg_20_ ( .D(csr_N1579), .CLK(csr_net35137), .Q(
        csr_n1920) );
  DFFX1_LVT csr_reg_misa_reg_23_ ( .D(csr_N1582), .CLK(csr_net35137), .Q(
        csr_n1919) );
  DFFX1_LVT csr_reg_misa_reg_63_ ( .D(csr_N1622), .CLK(csr_net35137), .Q(
        csr_n_T_3678_63_) );
  DFFX1_LVT csr_reg_fflags_reg_2_ ( .D(csr_n_GEN_345[2]), .CLK(csr_n594), .Q(
        csr_read_fcsr_2_), .QN(csr_n477) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_2_ ( .D(csr_n_GEN_258[2]), .CLK(csr_n533), 
        .Q(io_ptw_pmp_0_addr[2]) );
  DFFX1_LVT csr_u_T_47_reg_2_ ( .D(csr_N1824), .CLK(csr_n591), .Q(
        csr_io_time[2]) );
  DFFX1_LVT csr_u_T_39_reg_2_ ( .D(csr_N1430), .CLK(csr_n594), .Q(
        csr_n_T_45_2_) );
  DFFSSRX1_LVT csr_reg_dcsr_step_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_2_), .CLK(csr_net35162), .Q(csr_n_T_389_2), .QN(csr_n452) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_2_ ( .D(csr_n376), .SETB(csr_wdata_2_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_2_) );
  DFFX1_LVT csr_reg_stvec_reg_2_ ( .D(csr_n1483), .CLK(csr_n568), .QN(
        csr_reg_stvec_2_) );
  DFFX1_LVT csr_reg_frm_reg_2_ ( .D(csr_n_GEN_155[2]), .CLK(csr_net34900), .Q(
        io_fpu_fcsr_rm[2]) );
  DFFX1_LVT csr_reg_mie_reg_7_ ( .D(csr_N613), .CLK(csr_net34728), .Q(
        csr_reg_mie_7_) );
  DFFX1_LVT csr_u_T_49_reg_1_ ( .D(csr_N1892), .CLK(csr_n521), .Q(
        csr_io_time[7]) );
  DFFX1_LVT csr_u_T_41_reg_1_ ( .D(csr_N1498), .CLK(csr_n579), .Q(
        csr_n_T_45_7_) );
  DFFX1_LVT csr_reg_pmp_0_cfg_r_reg ( .D(csr_wdata_0_), .CLK(csr_net34733), 
        .Q(io_ptw_pmp_0_cfg_r) );
  DFFSSRX1_LVT csr_reg_pmp_0_cfg_l_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_7_), .CLK(csr_net34905), .Q(io_ptw_pmp_0_cfg_l), .QN(
        csr_n453) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_7_ ( .D(csr_n376), .SETB(csr_wdata_7_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_7_) );
  DFFX1_LVT csr_reg_sscratch_reg_7_ ( .D(csr_wdata_7_), .CLK(csr_n567), .Q(
        csr_reg_sscratch[7]) );
  DFFX1_LVT csr_reg_mscratch_reg_7_ ( .D(csr_wdata_7_), .CLK(csr_n553), .Q(
        csr_reg_mscratch[7]) );
  DFFX1_LVT csr_reg_dscratch_reg_7_ ( .D(csr_wdata_7_), .CLK(csr_n527), .Q(
        csr_reg_dscratch[7]) );
  DFFX1_LVT csr_reg_stvec_reg_7_ ( .D(csr_wdata_7_), .CLK(csr_n568), .Q(
        csr_reg_stvec_7_) );
  DFFX1_LVT csr_reg_mstatus_mpie_reg ( .D(csr_N360), .CLK(csr_net35147), .Q(
        csr_n1932) );
  DFFX1_LVT csr_reg_mideleg_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_net35167), .Q(
        csr_read_mideleg_9_), .QN(csr_n446) );
  DFFX1_LVT csr_reg_stvec_reg_9_ ( .D(csr_wdata_9_), .CLK(csr_n568), .Q(
        csr_reg_stvec_9_) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_9_ ( .D(csr_n_GEN_258[9]), .CLK(csr_n534), 
        .Q(io_ptw_pmp_0_addr[9]), .QN(csr_n419) );
  DFFX1_LVT csr_reg_pmp_0_addr_reg_0_ ( .D(csr_n_GEN_258[0]), .CLK(csr_n531), 
        .Q(io_ptw_pmp_0_addr[0]) );
  DFFSSRX1_LVT csr_reg_pmp_1_cfg_a_reg_1_ ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_12_), .CLK(csr_net35132), .Q(io_ptw_pmp_1_cfg_a[1]), .QN(
        csr_n462) );
  DFFX1_LVT csr_u_T_49_reg_6_ ( .D(csr_N1897), .CLK(csr_n521), .Q(
        csr_io_time[12]) );
  DFFX1_LVT csr_u_T_41_reg_6_ ( .D(csr_N1503), .CLK(csr_n579), .Q(
        csr_n_T_45_12_) );
  DFFSSRX1_LVT csr_reg_dcsr_ebreaku_reg ( .D(csr_n375), .SETB(1'b1), .RSTB(
        csr_wdata_12_), .CLK(csr_net35162), .Q(csr_n_T_1155_0_) );
  DFFSSRX1_LVT csr_reg_mtvec_reg_12_ ( .D(csr_n378), .SETB(csr_wdata_12_), 
        .RSTB(1'b1), .CLK(csr_n554), .QN(csr_reg_mtvec_12_) );
  DFFX1_LVT csr_reg_stvec_reg_12_ ( .D(csr_n367), .CLK(csr_n568), .QN(
        csr_reg_stvec_12_) );
  DFFX1_LVT csr_reg_mstatus_mpp_reg_1_ ( .D(csr_N334), .CLK(csr_net35147), .Q(
        csr_n_1929_) );
  DFFX1_LVT csr_reg_dcsr_prv_reg_0_ ( .D(csr_n2156), .CLK(csr_n594), .Q(
        csr_n_T_389_0) );
  DFFX1_LVT csr_reg_fflags_reg_0_ ( .D(csr_n_GEN_345[0]), .CLK(csr_n594), .Q(
        csr_read_fcsr_0_) );
  DFFX1_LVT csr_u_T_39_reg_0_ ( .D(csr_N1428), .CLK(csr_n594), .Q(
        csr_n_T_45_0_) );
  DFFX1_LVT csr_reg_sscratch_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_n567), .Q(
        csr_reg_sscratch[0]) );
  DFFX1_LVT csr_reg_mscratch_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_n553), .Q(
        csr_reg_mscratch[0]) );
  DFFX1_LVT csr_reg_dscratch_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_n527), .Q(
        csr_reg_dscratch[0]) );
  DFFX1_LVT csr_reg_medeleg_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_net35172), .Q(
        csr_read_medeleg_0) );
  DFFX1_LVT csr_reg_mcounteren_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_net34945), 
        .Q(csr_read_mcounteren_0_), .QN(csr_n470) );
  DFFX1_LVT csr_reg_scounteren_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_net34940), 
        .Q(csr_read_scounteren_0_) );
  DFFX1_LVT csr_reg_stvec_reg_0_ ( .D(csr_wdata_0_), .CLK(csr_n568), .Q(
        csr_n428), .QN(csr_n658) );
  DFFX1_LVT csr_u_T_47_reg_0_ ( .D(csr_N1822), .CLK(csr_n591), .Q(
        csr_io_time[0]), .QN(csr_n417) );
  DFFX1_LVT csr_u_T_1579_reg ( .D(csr_N1693), .CLK(csr_net35147), .Q(csr_n1918) );
  DFFX1_LVT csr_reg_mip_stip_reg ( .D(csr_n199), .CLK(csr_n531), .Q(
        csr_n_T_61_5_) );
  DFFX1_LVT csr_reg_mip_seip_reg ( .D(csr_n200), .CLK(csr_n531), .Q(
        csr_n_T_3694_9_) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_1 csr_clk_gate__T_49_reg ( .CLK(csr_n591), .EN(
        csr_N1890), .ENCLK(csr_net35324), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_2 csr_clk_gate_reg_bp_0_control_tmatch_reg ( 
        .CLK(csr_n593), .EN(csr_N487), .ENCLK(csr_net35319), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_3 csr_clk_gate_reg_bp_0_control_dmode_reg ( 
        .CLK(csr_n593), .EN(csr_N479), .ENCLK(csr_net35314), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_4 csr_clk_gate_reg_dscratch_reg ( .CLK(csr_n593), .EN(csr_N475), .ENCLK(csr_net35309), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_5 csr_clk_gate_reg_dpc_reg ( .CLK(csr_n593), 
        .EN(csr_net35183), .ENCLK(csr_net35304), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_6 csr_clk_gate_reg_dcsr_cause_reg ( .CLK(
        csr_n593), .EN(csr_N467), .ENCLK(csr_net35177), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_7 csr_clk_gate_reg_medeleg_reg ( .CLK(csr_n593), 
        .EN(csr_N460), .ENCLK(csr_net35172), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_8 csr_clk_gate_reg_mideleg_reg ( .CLK(csr_n593), 
        .EN(csr_N459), .ENCLK(csr_net35167), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_9 csr_clk_gate_reg_dcsr_ebreakm_reg ( .CLK(
        csr_n593), .EN(csr_N438), .ENCLK(csr_net35162), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_10 csr_clk_gate_reg_mstatus_mxr_reg ( .CLK(
        csr_n593), .EN(csr_N290), .ENCLK(csr_net35157), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_11 csr_clk_gate_reg_mstatus_tsr_reg ( .CLK(
        csr_n593), .EN(csr_N276), .ENCLK(csr_net35152), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_12 csr_clk_gate_reg_mstatus_mpp_reg ( .CLK(
        csr_n592), .EN(csr_N335), .ENCLK(csr_net35147), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_14 csr_clk_gate_reg_misa_reg ( .CLK(csr_n592), 
        .EN(csr_N1558), .ENCLK(csr_net35137), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_15 csr_clk_gate_reg_pmp_1_cfg_a_reg ( .CLK(
        csr_n592), .EN(csr_N527), .ENCLK(csr_net35132), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_16 csr_clk_gate_reg_pmp_3_cfg_a_reg ( .CLK(
        csr_n592), .EN(csr_N551), .ENCLK(csr_net35127), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_17 csr_clk_gate_reg_pmp_3_cfg_r_reg ( .CLK(
        csr_n592), .EN(csr_N556), .ENCLK(csr_net35122), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_18 csr_clk_gate_reg_pmp_4_cfg_r_reg ( .CLK(
        csr_n592), .EN(csr_N568), .ENCLK(csr_net35117), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_19 csr_clk_gate_reg_pmp_5_cfg_a_reg ( .CLK(
        csr_n592), .EN(csr_N575), .ENCLK(csr_net35112), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_20 csr_clk_gate_reg_pmp_6_cfg_r_reg ( .CLK(
        csr_n592), .EN(csr_N592), .ENCLK(csr_net35107), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_21 csr_clk_gate_reg_pmp_6_cfg_a_reg ( .CLK(
        csr_n592), .EN(csr_N587), .ENCLK(csr_net35102), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_22 csr_clk_gate_reg_pmp_5_cfg_r_reg ( .CLK(
        csr_n592), .EN(csr_N580), .ENCLK(csr_net35097), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_23 csr_clk_gate_reg_pmp_6_addr_reg ( .CLK(
        csr_n592), .EN(csr_n504), .ENCLK(csr_net35092), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_24 csr_clk_gate_reg_pmp_1_cfg_w_reg ( .CLK(
        csr_n593), .EN(csr_N531), .ENCLK(csr_net35087), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_25 csr_clk_gate_reg_mepc_reg ( .CLK(csr_n593), 
        .EN(csr_net34961), .ENCLK(csr_net35082), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_26 csr_clk_gate_reg_mscratch_reg ( .CLK(
        csr_n593), .EN(csr_N1033), .ENCLK(csr_net34955), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_27 csr_clk_gate_reg_mtvec_reg ( .CLK(csr_n593), 
        .EN(csr_n2165), .ENCLK(csr_net34950), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_28 csr_clk_gate_reg_mcounteren_reg ( .CLK(
        csr_n593), .EN(csr_n2169), .ENCLK(csr_net34945), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_29 csr_clk_gate_reg_scounteren_reg ( .CLK(
        csr_n593), .EN(csr_n2168), .ENCLK(csr_net34940), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_30 csr_clk_gate_reg_scause_reg ( .CLK(csr_n593), 
        .EN(csr_N1269), .ENCLK(csr_net34935), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_31 csr_clk_gate_reg_stval_reg ( .CLK(csr_n593), 
        .EN(csr_N1381), .ENCLK(csr_net34930), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_32 csr_clk_gate_reg_sscratch_reg ( .CLK(
        csr_n593), .EN(csr_N1422), .ENCLK(csr_net34925), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_33 csr_clk_gate_reg_stvec_reg ( .CLK(csr_n593), 
        .EN(csr_n2167), .ENCLK(csr_net34920), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_34 csr_clk_gate_reg_satp_ppn_reg ( .CLK(
        csr_n593), .EN(csr_N1426), .ENCLK(csr_net34915), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_35 csr_clk_gate_reg_pmp_4_cfg_l_reg ( .CLK(
        csr_n593), .EN(csr_N559), .ENCLK(csr_net34910), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_36 csr_clk_gate_reg_pmp_0_cfg_a_reg ( .CLK(
        csr_n593), .EN(csr_N515), .ENCLK(csr_net34905), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_37 csr_clk_gate_reg_frm_reg ( .CLK(csr_n593), 
        .EN(csr_n2166), .ENCLK(csr_net34900), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_38 csr_clk_gate_reg_mtval_reg ( .CLK(csr_n593), 
        .EN(csr_N992), .ENCLK(csr_net34895), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_39 csr_clk_gate__T_41_reg ( .CLK(csr_n593), 
        .EN(csr_N1496), .ENCLK(csr_net34890), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_40 csr_clk_gate_reg_mcause_reg ( .CLK(csr_n593), 
        .EN(csr_N880), .ENCLK(csr_net34885), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_41 csr_clk_gate_reg_sepc_reg ( .CLK(csr_n593), 
        .EN(csr_net34759), .ENCLK(csr_net34880), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_42 csr_clk_gate_reg_pmp_2_cfg_a_reg ( .CLK(
        csr_n593), .EN(csr_N539), .ENCLK(csr_net34753), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_43 csr_clk_gate_reg_pmp_2_cfg_x_reg ( .CLK(
        csr_n593), .EN(csr_N542), .ENCLK(csr_net34748), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_44 csr_clk_gate_reg_pmp_7_cfg_l_reg ( .CLK(
        csr_n593), .EN(csr_N595), .ENCLK(csr_net34743), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_45 csr_clk_gate_reg_pmp_7_cfg_r_reg ( .CLK(
        csr_n593), .EN(csr_N604), .ENCLK(csr_net34738), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_46 csr_clk_gate_reg_pmp_0_cfg_x_reg ( .CLK(
        csr_n594), .EN(csr_N518), .ENCLK(csr_net34733), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_47 csr_clk_gate_reg_mie_reg ( .CLK(csr_n594), 
        .EN(csr_N670), .ENCLK(csr_net34728), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_0 csr_clk_gate_reg_bp_0_address_reg ( .CLK(
        csr_n594), .EN(csr_n2163), .ENCLK(csr_net34722), .TE(1'b0) );
  NAND3X0_LVT csr_add_x_427_U194 ( .A1(csr_add_x_427_n93), .A2(
        io_ptw_pmp_7_addr[1]), .A3(io_ptw_pmp_7_addr[2]), .Y(
        csr_add_x_427_n176) );
  AND3X1_LVT csr_add_x_427_U193 ( .A1(io_ptw_pmp_7_addr[3]), .A2(
        io_ptw_pmp_7_addr[4]), .A3(csr_add_x_427_n170), .Y(csr_add_x_427_n174)
         );
  NAND3X0_LVT csr_add_x_427_U192 ( .A1(io_ptw_pmp_7_addr[5]), .A2(
        io_ptw_pmp_7_addr[6]), .A3(csr_add_x_427_n174), .Y(csr_add_x_427_n172)
         );
  AND3X1_LVT csr_add_x_427_U191 ( .A1(csr_add_x_427_n168), .A2(
        io_ptw_pmp_7_addr[8]), .A3(io_ptw_pmp_7_addr[7]), .Y(
        csr_add_x_427_n199) );
  HADDX1_LVT csr_add_x_427_U190 ( .A0(io_ptw_pmp_7_addr[9]), .B0(
        csr_add_x_427_n199), .SO(csr_n_T_304[10]) );
  AND4X1_LVT csr_add_x_427_U189 ( .A1(csr_add_x_427_n168), .A2(
        io_ptw_pmp_7_addr[8]), .A3(io_ptw_pmp_7_addr[7]), .A4(
        io_ptw_pmp_7_addr[9]), .Y(csr_add_x_427_n198) );
  HADDX1_LVT csr_add_x_427_U188 ( .A0(io_ptw_pmp_7_addr[10]), .B0(
        csr_add_x_427_n198), .SO(csr_n_T_304[11]) );
  AND4X1_LVT csr_add_x_427_U187 ( .A1(io_ptw_pmp_7_addr[8]), .A2(
        io_ptw_pmp_7_addr[7]), .A3(io_ptw_pmp_7_addr[10]), .A4(
        io_ptw_pmp_7_addr[9]), .Y(csr_add_x_427_n197) );
  NAND2X0_LVT csr_add_x_427_U186 ( .A1(csr_add_x_427_n168), .A2(
        csr_add_x_427_n197), .Y(csr_add_x_427_n196) );
  AO22X1_LVT csr_add_x_427_U185 ( .A1(io_ptw_pmp_7_addr[11]), .A2(
        csr_add_x_427_n196), .A3(csr_add_x_427_n165), .A4(csr_add_x_427_n166), 
        .Y(csr_n_T_304[12]) );
  AND2X1_LVT csr_add_x_427_U184 ( .A1(csr_add_x_427_n166), .A2(
        io_ptw_pmp_7_addr[11]), .Y(csr_add_x_427_n195) );
  HADDX1_LVT csr_add_x_427_U183 ( .A0(csr_add_x_427_n195), .B0(
        io_ptw_pmp_7_addr[12]), .SO(csr_n_T_304[13]) );
  AND3X1_LVT csr_add_x_427_U182 ( .A1(io_ptw_pmp_7_addr[11]), .A2(
        io_ptw_pmp_7_addr[12]), .A3(csr_add_x_427_n166), .Y(csr_add_x_427_n193) );
  HADDX1_LVT csr_add_x_427_U181 ( .A0(io_ptw_pmp_7_addr[13]), .B0(
        csr_add_x_427_n193), .SO(csr_n_T_304[14]) );
  AND4X1_LVT csr_add_x_427_U180 ( .A1(io_ptw_pmp_7_addr[11]), .A2(
        io_ptw_pmp_7_addr[12]), .A3(io_ptw_pmp_7_addr[13]), .A4(
        csr_add_x_427_n166), .Y(csr_add_x_427_n194) );
  HADDX1_LVT csr_add_x_427_U179 ( .A0(io_ptw_pmp_7_addr[14]), .B0(
        csr_add_x_427_n194), .SO(csr_n_T_304[15]) );
  NAND3X0_LVT csr_add_x_427_U178 ( .A1(io_ptw_pmp_7_addr[13]), .A2(
        io_ptw_pmp_7_addr[14]), .A3(csr_add_x_427_n193), .Y(csr_add_x_427_n192) );
  AO22X1_LVT csr_add_x_427_U177 ( .A1(io_ptw_pmp_7_addr[15]), .A2(
        csr_add_x_427_n192), .A3(csr_add_x_427_n163), .A4(csr_add_x_427_n164), 
        .Y(csr_n_T_304[16]) );
  AND2X1_LVT csr_add_x_427_U176 ( .A1(csr_add_x_427_n164), .A2(
        io_ptw_pmp_7_addr[15]), .Y(csr_add_x_427_n191) );
  HADDX1_LVT csr_add_x_427_U175 ( .A0(csr_add_x_427_n191), .B0(
        io_ptw_pmp_7_addr[16]), .SO(csr_n_T_304[17]) );
  AND3X1_LVT csr_add_x_427_U174 ( .A1(io_ptw_pmp_7_addr[15]), .A2(
        io_ptw_pmp_7_addr[16]), .A3(csr_add_x_427_n164), .Y(csr_add_x_427_n190) );
  HADDX1_LVT csr_add_x_427_U173 ( .A0(io_ptw_pmp_7_addr[17]), .B0(
        csr_add_x_427_n190), .SO(csr_n_T_304[18]) );
  AND4X1_LVT csr_add_x_427_U172 ( .A1(io_ptw_pmp_7_addr[15]), .A2(
        io_ptw_pmp_7_addr[16]), .A3(io_ptw_pmp_7_addr[17]), .A4(
        csr_add_x_427_n164), .Y(csr_add_x_427_n189) );
  HADDX1_LVT csr_add_x_427_U171 ( .A0(io_ptw_pmp_7_addr[18]), .B0(
        csr_add_x_427_n189), .SO(csr_n_T_304[19]) );
  AND4X1_LVT csr_add_x_427_U170 ( .A1(io_ptw_pmp_7_addr[15]), .A2(
        io_ptw_pmp_7_addr[16]), .A3(io_ptw_pmp_7_addr[18]), .A4(
        io_ptw_pmp_7_addr[17]), .Y(csr_add_x_427_n188) );
  NAND2X0_LVT csr_add_x_427_U169 ( .A1(csr_add_x_427_n188), .A2(
        csr_add_x_427_n164), .Y(csr_add_x_427_n187) );
  AO22X1_LVT csr_add_x_427_U168 ( .A1(io_ptw_pmp_7_addr[19]), .A2(
        csr_add_x_427_n187), .A3(csr_add_x_427_n161), .A4(csr_add_x_427_n162), 
        .Y(csr_n_T_304[20]) );
  AND2X1_LVT csr_add_x_427_U167 ( .A1(csr_add_x_427_n162), .A2(
        io_ptw_pmp_7_addr[19]), .Y(csr_add_x_427_n186) );
  HADDX1_LVT csr_add_x_427_U166 ( .A0(csr_add_x_427_n186), .B0(
        io_ptw_pmp_7_addr[20]), .SO(csr_n_T_304[21]) );
  AND3X1_LVT csr_add_x_427_U165 ( .A1(io_ptw_pmp_7_addr[19]), .A2(
        io_ptw_pmp_7_addr[20]), .A3(csr_add_x_427_n162), .Y(csr_add_x_427_n184) );
  HADDX1_LVT csr_add_x_427_U164 ( .A0(io_ptw_pmp_7_addr[21]), .B0(
        csr_add_x_427_n184), .SO(csr_n_T_304[22]) );
  AND2X1_LVT csr_add_x_427_U163 ( .A1(csr_add_x_427_n184), .A2(
        io_ptw_pmp_7_addr[21]), .Y(csr_add_x_427_n185) );
  HADDX1_LVT csr_add_x_427_U162 ( .A0(csr_add_x_427_n185), .B0(
        io_ptw_pmp_7_addr[22]), .SO(csr_n_T_304[23]) );
  NAND3X0_LVT csr_add_x_427_U161 ( .A1(io_ptw_pmp_7_addr[22]), .A2(
        io_ptw_pmp_7_addr[21]), .A3(csr_add_x_427_n184), .Y(csr_add_x_427_n183) );
  AO22X1_LVT csr_add_x_427_U160 ( .A1(io_ptw_pmp_7_addr[23]), .A2(
        csr_add_x_427_n183), .A3(csr_add_x_427_n159), .A4(csr_add_x_427_n160), 
        .Y(csr_n_T_304[24]) );
  AND2X1_LVT csr_add_x_427_U159 ( .A1(csr_add_x_427_n160), .A2(
        io_ptw_pmp_7_addr[23]), .Y(csr_add_x_427_n182) );
  HADDX1_LVT csr_add_x_427_U158 ( .A0(csr_add_x_427_n182), .B0(
        io_ptw_pmp_7_addr[24]), .SO(csr_n_T_304[25]) );
  AND3X1_LVT csr_add_x_427_U157 ( .A1(io_ptw_pmp_7_addr[23]), .A2(
        io_ptw_pmp_7_addr[24]), .A3(csr_add_x_427_n160), .Y(csr_add_x_427_n181) );
  HADDX1_LVT csr_add_x_427_U156 ( .A0(io_ptw_pmp_7_addr[25]), .B0(
        csr_add_x_427_n181), .SO(csr_n_T_304[26]) );
  AND2X1_LVT csr_add_x_427_U155 ( .A1(io_ptw_pmp_7_addr[25]), .A2(
        csr_add_x_427_n181), .Y(csr_add_x_427_n179) );
  HADDX1_LVT csr_add_x_427_U154 ( .A0(io_ptw_pmp_7_addr[26]), .B0(
        csr_add_x_427_n179), .SO(csr_n_T_304[27]) );
  AND2X1_LVT csr_add_x_427_U153 ( .A1(io_ptw_pmp_7_addr[26]), .A2(
        csr_add_x_427_n179), .Y(csr_add_x_427_n180) );
  HADDX1_LVT csr_add_x_427_U152 ( .A0(csr_add_x_427_n180), .B0(
        io_ptw_pmp_7_addr[27]), .SO(csr_n_T_304[28]) );
  AND3X1_LVT csr_add_x_427_U151 ( .A1(csr_add_x_427_n179), .A2(
        io_ptw_pmp_7_addr[26]), .A3(io_ptw_pmp_7_addr[27]), .Y(
        csr_add_x_427_n178) );
  HADDX1_LVT csr_add_x_427_U150 ( .A0(csr_add_x_427_n178), .B0(
        io_ptw_pmp_7_addr[28]), .SO(csr_n_T_304[29]) );
  HADDX1_LVT csr_add_x_427_U149 ( .A0(csr_add_x_427_n93), .B0(
        io_ptw_pmp_7_addr[1]), .SO(csr_n_T_304[2]) );
  AND2X1_LVT csr_add_x_427_U148 ( .A1(csr_add_x_427_n93), .A2(
        io_ptw_pmp_7_addr[1]), .Y(csr_add_x_427_n177) );
  HADDX1_LVT csr_add_x_427_U147 ( .A0(io_ptw_pmp_7_addr[2]), .B0(
        csr_add_x_427_n177), .SO(csr_n_T_304[3]) );
  AO22X1_LVT csr_add_x_427_U146 ( .A1(io_ptw_pmp_7_addr[3]), .A2(
        csr_add_x_427_n176), .A3(csr_add_x_427_n169), .A4(csr_add_x_427_n170), 
        .Y(csr_n_T_304[4]) );
  AND2X1_LVT csr_add_x_427_U145 ( .A1(csr_add_x_427_n170), .A2(
        io_ptw_pmp_7_addr[3]), .Y(csr_add_x_427_n175) );
  HADDX1_LVT csr_add_x_427_U144 ( .A0(csr_add_x_427_n175), .B0(
        io_ptw_pmp_7_addr[4]), .SO(csr_n_T_304[5]) );
  HADDX1_LVT csr_add_x_427_U143 ( .A0(io_ptw_pmp_7_addr[5]), .B0(
        csr_add_x_427_n174), .SO(csr_n_T_304[6]) );
  AND2X1_LVT csr_add_x_427_U142 ( .A1(io_ptw_pmp_7_addr[5]), .A2(
        csr_add_x_427_n174), .Y(csr_add_x_427_n173) );
  HADDX1_LVT csr_add_x_427_U141 ( .A0(io_ptw_pmp_7_addr[6]), .B0(
        csr_add_x_427_n173), .SO(csr_n_T_304[7]) );
  AO22X1_LVT csr_add_x_427_U140 ( .A1(csr_add_x_427_n168), .A2(
        csr_add_x_427_n167), .A3(csr_add_x_427_n172), .A4(io_ptw_pmp_7_addr[7]), .Y(csr_n_T_304[8]) );
  AND2X1_LVT csr_add_x_427_U139 ( .A1(io_ptw_pmp_7_addr[7]), .A2(
        csr_add_x_427_n168), .Y(csr_add_x_427_n171) );
  HADDX1_LVT csr_add_x_427_U138 ( .A0(csr_add_x_427_n171), .B0(
        io_ptw_pmp_7_addr[8]), .SO(csr_n_T_304[9]) );
  INVX1_LVT csr_add_x_427_U137 ( .A(csr_add_x_427_n176), .Y(csr_add_x_427_n170) );
  INVX1_LVT csr_add_x_427_U136 ( .A(io_ptw_pmp_7_addr[3]), .Y(
        csr_add_x_427_n169) );
  INVX1_LVT csr_add_x_427_U135 ( .A(csr_add_x_427_n172), .Y(csr_add_x_427_n168) );
  INVX1_LVT csr_add_x_427_U134 ( .A(io_ptw_pmp_7_addr[7]), .Y(
        csr_add_x_427_n167) );
  INVX1_LVT csr_add_x_427_U133 ( .A(csr_add_x_427_n196), .Y(csr_add_x_427_n166) );
  INVX1_LVT csr_add_x_427_U132 ( .A(io_ptw_pmp_7_addr[11]), .Y(
        csr_add_x_427_n165) );
  INVX1_LVT csr_add_x_427_U131 ( .A(csr_add_x_427_n192), .Y(csr_add_x_427_n164) );
  INVX1_LVT csr_add_x_427_U130 ( .A(io_ptw_pmp_7_addr[15]), .Y(
        csr_add_x_427_n163) );
  INVX1_LVT csr_add_x_427_U129 ( .A(csr_add_x_427_n187), .Y(csr_add_x_427_n162) );
  INVX1_LVT csr_add_x_427_U128 ( .A(io_ptw_pmp_7_addr[19]), .Y(
        csr_add_x_427_n161) );
  INVX1_LVT csr_add_x_427_U127 ( .A(csr_add_x_427_n183), .Y(csr_add_x_427_n160) );
  INVX1_LVT csr_add_x_427_U126 ( .A(io_ptw_pmp_7_addr[23]), .Y(
        csr_add_x_427_n159) );
  HADDX1_LVT csr_add_x_427_U121 ( .A0(io_ptw_pmp_7_addr[0]), .B0(
        io_ptw_pmp_7_cfg_a[0]), .C1(csr_add_x_427_n93), .SO(csr_n_T_304[1]) );
  NAND3X0_LVT csr_add_x_426_U194 ( .A1(csr_add_x_426_n93), .A2(
        io_ptw_pmp_6_addr[1]), .A3(io_ptw_pmp_6_addr[2]), .Y(
        csr_add_x_426_n176) );
  AND3X1_LVT csr_add_x_426_U193 ( .A1(io_ptw_pmp_6_addr[3]), .A2(
        io_ptw_pmp_6_addr[4]), .A3(csr_add_x_426_n170), .Y(csr_add_x_426_n174)
         );
  NAND3X0_LVT csr_add_x_426_U192 ( .A1(io_ptw_pmp_6_addr[5]), .A2(
        io_ptw_pmp_6_addr[6]), .A3(csr_add_x_426_n174), .Y(csr_add_x_426_n172)
         );
  AND3X1_LVT csr_add_x_426_U191 ( .A1(csr_add_x_426_n168), .A2(
        io_ptw_pmp_6_addr[8]), .A3(io_ptw_pmp_6_addr[7]), .Y(
        csr_add_x_426_n199) );
  HADDX1_LVT csr_add_x_426_U190 ( .A0(io_ptw_pmp_6_addr[9]), .B0(
        csr_add_x_426_n199), .SO(csr_n_T_295[10]) );
  AND4X1_LVT csr_add_x_426_U189 ( .A1(csr_add_x_426_n168), .A2(
        io_ptw_pmp_6_addr[8]), .A3(io_ptw_pmp_6_addr[7]), .A4(
        io_ptw_pmp_6_addr[9]), .Y(csr_add_x_426_n198) );
  HADDX1_LVT csr_add_x_426_U188 ( .A0(io_ptw_pmp_6_addr[10]), .B0(
        csr_add_x_426_n198), .SO(csr_n_T_295[11]) );
  AND4X1_LVT csr_add_x_426_U187 ( .A1(io_ptw_pmp_6_addr[8]), .A2(
        io_ptw_pmp_6_addr[7]), .A3(io_ptw_pmp_6_addr[10]), .A4(
        io_ptw_pmp_6_addr[9]), .Y(csr_add_x_426_n197) );
  NAND2X0_LVT csr_add_x_426_U186 ( .A1(csr_add_x_426_n168), .A2(
        csr_add_x_426_n197), .Y(csr_add_x_426_n196) );
  AO22X1_LVT csr_add_x_426_U185 ( .A1(io_ptw_pmp_6_addr[11]), .A2(
        csr_add_x_426_n196), .A3(csr_add_x_426_n165), .A4(csr_add_x_426_n166), 
        .Y(csr_n_T_295[12]) );
  AND2X1_LVT csr_add_x_426_U184 ( .A1(csr_add_x_426_n166), .A2(
        io_ptw_pmp_6_addr[11]), .Y(csr_add_x_426_n195) );
  HADDX1_LVT csr_add_x_426_U183 ( .A0(csr_add_x_426_n195), .B0(
        io_ptw_pmp_6_addr[12]), .SO(csr_n_T_295[13]) );
  AND3X1_LVT csr_add_x_426_U182 ( .A1(io_ptw_pmp_6_addr[11]), .A2(
        io_ptw_pmp_6_addr[12]), .A3(csr_add_x_426_n166), .Y(csr_add_x_426_n193) );
  HADDX1_LVT csr_add_x_426_U181 ( .A0(io_ptw_pmp_6_addr[13]), .B0(
        csr_add_x_426_n193), .SO(csr_n_T_295[14]) );
  AND4X1_LVT csr_add_x_426_U180 ( .A1(io_ptw_pmp_6_addr[11]), .A2(
        io_ptw_pmp_6_addr[12]), .A3(io_ptw_pmp_6_addr[13]), .A4(
        csr_add_x_426_n166), .Y(csr_add_x_426_n194) );
  HADDX1_LVT csr_add_x_426_U179 ( .A0(io_ptw_pmp_6_addr[14]), .B0(
        csr_add_x_426_n194), .SO(csr_n_T_295[15]) );
  NAND3X0_LVT csr_add_x_426_U178 ( .A1(io_ptw_pmp_6_addr[13]), .A2(
        io_ptw_pmp_6_addr[14]), .A3(csr_add_x_426_n193), .Y(csr_add_x_426_n192) );
  AO22X1_LVT csr_add_x_426_U177 ( .A1(io_ptw_pmp_6_addr[15]), .A2(
        csr_add_x_426_n192), .A3(csr_add_x_426_n163), .A4(csr_add_x_426_n164), 
        .Y(csr_n_T_295[16]) );
  AND2X1_LVT csr_add_x_426_U176 ( .A1(csr_add_x_426_n164), .A2(
        io_ptw_pmp_6_addr[15]), .Y(csr_add_x_426_n191) );
  HADDX1_LVT csr_add_x_426_U175 ( .A0(csr_add_x_426_n191), .B0(
        io_ptw_pmp_6_addr[16]), .SO(csr_n_T_295[17]) );
  AND3X1_LVT csr_add_x_426_U174 ( .A1(io_ptw_pmp_6_addr[15]), .A2(
        io_ptw_pmp_6_addr[16]), .A3(csr_add_x_426_n164), .Y(csr_add_x_426_n190) );
  HADDX1_LVT csr_add_x_426_U173 ( .A0(io_ptw_pmp_6_addr[17]), .B0(
        csr_add_x_426_n190), .SO(csr_n_T_295[18]) );
  AND4X1_LVT csr_add_x_426_U172 ( .A1(io_ptw_pmp_6_addr[15]), .A2(
        io_ptw_pmp_6_addr[16]), .A3(io_ptw_pmp_6_addr[17]), .A4(
        csr_add_x_426_n164), .Y(csr_add_x_426_n189) );
  HADDX1_LVT csr_add_x_426_U171 ( .A0(io_ptw_pmp_6_addr[18]), .B0(
        csr_add_x_426_n189), .SO(csr_n_T_295[19]) );
  AND4X1_LVT csr_add_x_426_U170 ( .A1(io_ptw_pmp_6_addr[15]), .A2(
        io_ptw_pmp_6_addr[16]), .A3(io_ptw_pmp_6_addr[18]), .A4(
        io_ptw_pmp_6_addr[17]), .Y(csr_add_x_426_n188) );
  NAND2X0_LVT csr_add_x_426_U169 ( .A1(csr_add_x_426_n188), .A2(
        csr_add_x_426_n164), .Y(csr_add_x_426_n187) );
  AO22X1_LVT csr_add_x_426_U168 ( .A1(io_ptw_pmp_6_addr[19]), .A2(
        csr_add_x_426_n187), .A3(csr_add_x_426_n161), .A4(csr_add_x_426_n162), 
        .Y(csr_n_T_295[20]) );
  AND2X1_LVT csr_add_x_426_U167 ( .A1(csr_add_x_426_n162), .A2(
        io_ptw_pmp_6_addr[19]), .Y(csr_add_x_426_n186) );
  HADDX1_LVT csr_add_x_426_U166 ( .A0(csr_add_x_426_n186), .B0(
        io_ptw_pmp_6_addr[20]), .SO(csr_n_T_295[21]) );
  AND3X1_LVT csr_add_x_426_U165 ( .A1(io_ptw_pmp_6_addr[19]), .A2(
        io_ptw_pmp_6_addr[20]), .A3(csr_add_x_426_n162), .Y(csr_add_x_426_n184) );
  HADDX1_LVT csr_add_x_426_U164 ( .A0(io_ptw_pmp_6_addr[21]), .B0(
        csr_add_x_426_n184), .SO(csr_n_T_295[22]) );
  AND2X1_LVT csr_add_x_426_U163 ( .A1(csr_add_x_426_n184), .A2(
        io_ptw_pmp_6_addr[21]), .Y(csr_add_x_426_n185) );
  HADDX1_LVT csr_add_x_426_U162 ( .A0(csr_add_x_426_n185), .B0(
        io_ptw_pmp_6_addr[22]), .SO(csr_n_T_295[23]) );
  NAND3X0_LVT csr_add_x_426_U161 ( .A1(io_ptw_pmp_6_addr[22]), .A2(
        io_ptw_pmp_6_addr[21]), .A3(csr_add_x_426_n184), .Y(csr_add_x_426_n183) );
  AO22X1_LVT csr_add_x_426_U160 ( .A1(io_ptw_pmp_6_addr[23]), .A2(
        csr_add_x_426_n183), .A3(csr_add_x_426_n159), .A4(csr_add_x_426_n160), 
        .Y(csr_n_T_295[24]) );
  AND2X1_LVT csr_add_x_426_U159 ( .A1(csr_add_x_426_n160), .A2(
        io_ptw_pmp_6_addr[23]), .Y(csr_add_x_426_n182) );
  HADDX1_LVT csr_add_x_426_U158 ( .A0(csr_add_x_426_n182), .B0(
        io_ptw_pmp_6_addr[24]), .SO(csr_n_T_295[25]) );
  AND3X1_LVT csr_add_x_426_U157 ( .A1(io_ptw_pmp_6_addr[23]), .A2(
        io_ptw_pmp_6_addr[24]), .A3(csr_add_x_426_n160), .Y(csr_add_x_426_n181) );
  HADDX1_LVT csr_add_x_426_U156 ( .A0(io_ptw_pmp_6_addr[25]), .B0(
        csr_add_x_426_n181), .SO(csr_n_T_295[26]) );
  AND2X1_LVT csr_add_x_426_U155 ( .A1(io_ptw_pmp_6_addr[25]), .A2(
        csr_add_x_426_n181), .Y(csr_add_x_426_n179) );
  HADDX1_LVT csr_add_x_426_U154 ( .A0(io_ptw_pmp_6_addr[26]), .B0(
        csr_add_x_426_n179), .SO(csr_n_T_295[27]) );
  AND2X1_LVT csr_add_x_426_U153 ( .A1(io_ptw_pmp_6_addr[26]), .A2(
        csr_add_x_426_n179), .Y(csr_add_x_426_n180) );
  HADDX1_LVT csr_add_x_426_U152 ( .A0(csr_add_x_426_n180), .B0(
        io_ptw_pmp_6_addr[27]), .SO(csr_n_T_295[28]) );
  AND3X1_LVT csr_add_x_426_U151 ( .A1(csr_add_x_426_n179), .A2(
        io_ptw_pmp_6_addr[26]), .A3(io_ptw_pmp_6_addr[27]), .Y(
        csr_add_x_426_n178) );
  HADDX1_LVT csr_add_x_426_U150 ( .A0(csr_add_x_426_n178), .B0(
        io_ptw_pmp_6_addr[28]), .SO(csr_n_T_295[29]) );
  HADDX1_LVT csr_add_x_426_U149 ( .A0(csr_add_x_426_n93), .B0(
        io_ptw_pmp_6_addr[1]), .SO(csr_n_T_295[2]) );
  AND2X1_LVT csr_add_x_426_U148 ( .A1(csr_add_x_426_n93), .A2(
        io_ptw_pmp_6_addr[1]), .Y(csr_add_x_426_n177) );
  HADDX1_LVT csr_add_x_426_U147 ( .A0(io_ptw_pmp_6_addr[2]), .B0(
        csr_add_x_426_n177), .SO(csr_n_T_295[3]) );
  AO22X1_LVT csr_add_x_426_U146 ( .A1(io_ptw_pmp_6_addr[3]), .A2(
        csr_add_x_426_n176), .A3(csr_add_x_426_n169), .A4(csr_add_x_426_n170), 
        .Y(csr_n_T_295[4]) );
  AND2X1_LVT csr_add_x_426_U145 ( .A1(csr_add_x_426_n170), .A2(
        io_ptw_pmp_6_addr[3]), .Y(csr_add_x_426_n175) );
  HADDX1_LVT csr_add_x_426_U144 ( .A0(csr_add_x_426_n175), .B0(
        io_ptw_pmp_6_addr[4]), .SO(csr_n_T_295[5]) );
  HADDX1_LVT csr_add_x_426_U143 ( .A0(io_ptw_pmp_6_addr[5]), .B0(
        csr_add_x_426_n174), .SO(csr_n_T_295[6]) );
  AND2X1_LVT csr_add_x_426_U142 ( .A1(io_ptw_pmp_6_addr[5]), .A2(
        csr_add_x_426_n174), .Y(csr_add_x_426_n173) );
  HADDX1_LVT csr_add_x_426_U141 ( .A0(io_ptw_pmp_6_addr[6]), .B0(
        csr_add_x_426_n173), .SO(csr_n_T_295[7]) );
  AO22X1_LVT csr_add_x_426_U140 ( .A1(csr_add_x_426_n168), .A2(
        csr_add_x_426_n167), .A3(csr_add_x_426_n172), .A4(io_ptw_pmp_6_addr[7]), .Y(csr_n_T_295[8]) );
  AND2X1_LVT csr_add_x_426_U139 ( .A1(io_ptw_pmp_6_addr[7]), .A2(
        csr_add_x_426_n168), .Y(csr_add_x_426_n171) );
  HADDX1_LVT csr_add_x_426_U138 ( .A0(csr_add_x_426_n171), .B0(
        io_ptw_pmp_6_addr[8]), .SO(csr_n_T_295[9]) );
  INVX1_LVT csr_add_x_426_U137 ( .A(csr_add_x_426_n176), .Y(csr_add_x_426_n170) );
  INVX1_LVT csr_add_x_426_U136 ( .A(io_ptw_pmp_6_addr[3]), .Y(
        csr_add_x_426_n169) );
  INVX1_LVT csr_add_x_426_U135 ( .A(csr_add_x_426_n172), .Y(csr_add_x_426_n168) );
  INVX1_LVT csr_add_x_426_U134 ( .A(io_ptw_pmp_6_addr[7]), .Y(
        csr_add_x_426_n167) );
  INVX1_LVT csr_add_x_426_U133 ( .A(csr_add_x_426_n196), .Y(csr_add_x_426_n166) );
  INVX1_LVT csr_add_x_426_U132 ( .A(io_ptw_pmp_6_addr[11]), .Y(
        csr_add_x_426_n165) );
  INVX1_LVT csr_add_x_426_U131 ( .A(csr_add_x_426_n192), .Y(csr_add_x_426_n164) );
  INVX1_LVT csr_add_x_426_U130 ( .A(io_ptw_pmp_6_addr[15]), .Y(
        csr_add_x_426_n163) );
  INVX1_LVT csr_add_x_426_U129 ( .A(csr_add_x_426_n187), .Y(csr_add_x_426_n162) );
  INVX1_LVT csr_add_x_426_U128 ( .A(io_ptw_pmp_6_addr[19]), .Y(
        csr_add_x_426_n161) );
  INVX1_LVT csr_add_x_426_U127 ( .A(csr_add_x_426_n183), .Y(csr_add_x_426_n160) );
  INVX1_LVT csr_add_x_426_U126 ( .A(io_ptw_pmp_6_addr[23]), .Y(
        csr_add_x_426_n159) );
  HADDX1_LVT csr_add_x_426_U121 ( .A0(io_ptw_pmp_6_addr[0]), .B0(
        io_ptw_pmp_6_cfg_a[0]), .C1(csr_add_x_426_n93), .SO(csr_n_T_295[1]) );
  NAND3X0_LVT csr_add_x_425_U194 ( .A1(csr_add_x_425_n93), .A2(
        io_ptw_pmp_5_addr[1]), .A3(io_ptw_pmp_5_addr[2]), .Y(
        csr_add_x_425_n176) );
  AND3X1_LVT csr_add_x_425_U193 ( .A1(io_ptw_pmp_5_addr[3]), .A2(
        io_ptw_pmp_5_addr[4]), .A3(csr_add_x_425_n170), .Y(csr_add_x_425_n174)
         );
  NAND3X0_LVT csr_add_x_425_U192 ( .A1(io_ptw_pmp_5_addr[5]), .A2(
        io_ptw_pmp_5_addr[6]), .A3(csr_add_x_425_n174), .Y(csr_add_x_425_n172)
         );
  AND3X1_LVT csr_add_x_425_U191 ( .A1(csr_add_x_425_n168), .A2(
        io_ptw_pmp_5_addr[8]), .A3(io_ptw_pmp_5_addr[7]), .Y(
        csr_add_x_425_n199) );
  HADDX1_LVT csr_add_x_425_U190 ( .A0(io_ptw_pmp_5_addr[9]), .B0(
        csr_add_x_425_n199), .SO(csr_n_T_286[10]) );
  AND4X1_LVT csr_add_x_425_U189 ( .A1(csr_add_x_425_n168), .A2(
        io_ptw_pmp_5_addr[8]), .A3(io_ptw_pmp_5_addr[7]), .A4(
        io_ptw_pmp_5_addr[9]), .Y(csr_add_x_425_n198) );
  HADDX1_LVT csr_add_x_425_U188 ( .A0(io_ptw_pmp_5_addr[10]), .B0(
        csr_add_x_425_n198), .SO(csr_n_T_286[11]) );
  AND4X1_LVT csr_add_x_425_U187 ( .A1(io_ptw_pmp_5_addr[8]), .A2(
        io_ptw_pmp_5_addr[7]), .A3(io_ptw_pmp_5_addr[10]), .A4(
        io_ptw_pmp_5_addr[9]), .Y(csr_add_x_425_n197) );
  NAND2X0_LVT csr_add_x_425_U186 ( .A1(csr_add_x_425_n168), .A2(
        csr_add_x_425_n197), .Y(csr_add_x_425_n196) );
  AO22X1_LVT csr_add_x_425_U185 ( .A1(io_ptw_pmp_5_addr[11]), .A2(
        csr_add_x_425_n196), .A3(csr_add_x_425_n165), .A4(csr_add_x_425_n166), 
        .Y(csr_n_T_286[12]) );
  AND2X1_LVT csr_add_x_425_U184 ( .A1(csr_add_x_425_n166), .A2(
        io_ptw_pmp_5_addr[11]), .Y(csr_add_x_425_n195) );
  HADDX1_LVT csr_add_x_425_U183 ( .A0(csr_add_x_425_n195), .B0(
        io_ptw_pmp_5_addr[12]), .SO(csr_n_T_286[13]) );
  AND3X1_LVT csr_add_x_425_U182 ( .A1(io_ptw_pmp_5_addr[11]), .A2(
        io_ptw_pmp_5_addr[12]), .A3(csr_add_x_425_n166), .Y(csr_add_x_425_n193) );
  HADDX1_LVT csr_add_x_425_U181 ( .A0(io_ptw_pmp_5_addr[13]), .B0(
        csr_add_x_425_n193), .SO(csr_n_T_286[14]) );
  AND4X1_LVT csr_add_x_425_U180 ( .A1(io_ptw_pmp_5_addr[11]), .A2(
        io_ptw_pmp_5_addr[12]), .A3(io_ptw_pmp_5_addr[13]), .A4(
        csr_add_x_425_n166), .Y(csr_add_x_425_n194) );
  HADDX1_LVT csr_add_x_425_U179 ( .A0(io_ptw_pmp_5_addr[14]), .B0(
        csr_add_x_425_n194), .SO(csr_n_T_286[15]) );
  NAND3X0_LVT csr_add_x_425_U178 ( .A1(io_ptw_pmp_5_addr[13]), .A2(
        io_ptw_pmp_5_addr[14]), .A3(csr_add_x_425_n193), .Y(csr_add_x_425_n192) );
  AO22X1_LVT csr_add_x_425_U177 ( .A1(io_ptw_pmp_5_addr[15]), .A2(
        csr_add_x_425_n192), .A3(csr_add_x_425_n163), .A4(csr_add_x_425_n164), 
        .Y(csr_n_T_286[16]) );
  AND2X1_LVT csr_add_x_425_U176 ( .A1(csr_add_x_425_n164), .A2(
        io_ptw_pmp_5_addr[15]), .Y(csr_add_x_425_n191) );
  HADDX1_LVT csr_add_x_425_U175 ( .A0(csr_add_x_425_n191), .B0(
        io_ptw_pmp_5_addr[16]), .SO(csr_n_T_286[17]) );
  AND3X1_LVT csr_add_x_425_U174 ( .A1(io_ptw_pmp_5_addr[15]), .A2(
        io_ptw_pmp_5_addr[16]), .A3(csr_add_x_425_n164), .Y(csr_add_x_425_n190) );
  HADDX1_LVT csr_add_x_425_U173 ( .A0(io_ptw_pmp_5_addr[17]), .B0(
        csr_add_x_425_n190), .SO(csr_n_T_286[18]) );
  AND4X1_LVT csr_add_x_425_U172 ( .A1(io_ptw_pmp_5_addr[15]), .A2(
        io_ptw_pmp_5_addr[16]), .A3(io_ptw_pmp_5_addr[17]), .A4(
        csr_add_x_425_n164), .Y(csr_add_x_425_n189) );
  HADDX1_LVT csr_add_x_425_U171 ( .A0(io_ptw_pmp_5_addr[18]), .B0(
        csr_add_x_425_n189), .SO(csr_n_T_286[19]) );
  AND4X1_LVT csr_add_x_425_U170 ( .A1(io_ptw_pmp_5_addr[15]), .A2(
        io_ptw_pmp_5_addr[16]), .A3(io_ptw_pmp_5_addr[18]), .A4(
        io_ptw_pmp_5_addr[17]), .Y(csr_add_x_425_n188) );
  NAND2X0_LVT csr_add_x_425_U169 ( .A1(csr_add_x_425_n188), .A2(
        csr_add_x_425_n164), .Y(csr_add_x_425_n187) );
  AO22X1_LVT csr_add_x_425_U168 ( .A1(io_ptw_pmp_5_addr[19]), .A2(
        csr_add_x_425_n187), .A3(csr_add_x_425_n161), .A4(csr_add_x_425_n162), 
        .Y(csr_n_T_286[20]) );
  AND2X1_LVT csr_add_x_425_U167 ( .A1(csr_add_x_425_n162), .A2(
        io_ptw_pmp_5_addr[19]), .Y(csr_add_x_425_n186) );
  HADDX1_LVT csr_add_x_425_U166 ( .A0(csr_add_x_425_n186), .B0(
        io_ptw_pmp_5_addr[20]), .SO(csr_n_T_286[21]) );
  AND3X1_LVT csr_add_x_425_U165 ( .A1(io_ptw_pmp_5_addr[19]), .A2(
        io_ptw_pmp_5_addr[20]), .A3(csr_add_x_425_n162), .Y(csr_add_x_425_n184) );
  HADDX1_LVT csr_add_x_425_U164 ( .A0(io_ptw_pmp_5_addr[21]), .B0(
        csr_add_x_425_n184), .SO(csr_n_T_286[22]) );
  AND2X1_LVT csr_add_x_425_U163 ( .A1(csr_add_x_425_n184), .A2(
        io_ptw_pmp_5_addr[21]), .Y(csr_add_x_425_n185) );
  HADDX1_LVT csr_add_x_425_U162 ( .A0(csr_add_x_425_n185), .B0(
        io_ptw_pmp_5_addr[22]), .SO(csr_n_T_286[23]) );
  NAND3X0_LVT csr_add_x_425_U161 ( .A1(io_ptw_pmp_5_addr[22]), .A2(
        io_ptw_pmp_5_addr[21]), .A3(csr_add_x_425_n184), .Y(csr_add_x_425_n183) );
  AO22X1_LVT csr_add_x_425_U160 ( .A1(io_ptw_pmp_5_addr[23]), .A2(
        csr_add_x_425_n183), .A3(csr_add_x_425_n159), .A4(csr_add_x_425_n160), 
        .Y(csr_n_T_286[24]) );
  AND2X1_LVT csr_add_x_425_U159 ( .A1(csr_add_x_425_n160), .A2(
        io_ptw_pmp_5_addr[23]), .Y(csr_add_x_425_n182) );
  HADDX1_LVT csr_add_x_425_U158 ( .A0(csr_add_x_425_n182), .B0(
        io_ptw_pmp_5_addr[24]), .SO(csr_n_T_286[25]) );
  AND3X1_LVT csr_add_x_425_U157 ( .A1(io_ptw_pmp_5_addr[23]), .A2(
        io_ptw_pmp_5_addr[24]), .A3(csr_add_x_425_n160), .Y(csr_add_x_425_n181) );
  HADDX1_LVT csr_add_x_425_U156 ( .A0(io_ptw_pmp_5_addr[25]), .B0(
        csr_add_x_425_n181), .SO(csr_n_T_286[26]) );
  AND2X1_LVT csr_add_x_425_U155 ( .A1(io_ptw_pmp_5_addr[25]), .A2(
        csr_add_x_425_n181), .Y(csr_add_x_425_n179) );
  HADDX1_LVT csr_add_x_425_U154 ( .A0(io_ptw_pmp_5_addr[26]), .B0(
        csr_add_x_425_n179), .SO(csr_n_T_286[27]) );
  AND2X1_LVT csr_add_x_425_U153 ( .A1(io_ptw_pmp_5_addr[26]), .A2(
        csr_add_x_425_n179), .Y(csr_add_x_425_n180) );
  HADDX1_LVT csr_add_x_425_U152 ( .A0(csr_add_x_425_n180), .B0(
        io_ptw_pmp_5_addr[27]), .SO(csr_n_T_286[28]) );
  AND3X1_LVT csr_add_x_425_U151 ( .A1(csr_add_x_425_n179), .A2(
        io_ptw_pmp_5_addr[26]), .A3(io_ptw_pmp_5_addr[27]), .Y(
        csr_add_x_425_n178) );
  HADDX1_LVT csr_add_x_425_U150 ( .A0(csr_add_x_425_n178), .B0(
        io_ptw_pmp_5_addr[28]), .SO(csr_n_T_286[29]) );
  HADDX1_LVT csr_add_x_425_U149 ( .A0(csr_add_x_425_n93), .B0(
        io_ptw_pmp_5_addr[1]), .SO(csr_n_T_286[2]) );
  AND2X1_LVT csr_add_x_425_U148 ( .A1(csr_add_x_425_n93), .A2(
        io_ptw_pmp_5_addr[1]), .Y(csr_add_x_425_n177) );
  HADDX1_LVT csr_add_x_425_U147 ( .A0(io_ptw_pmp_5_addr[2]), .B0(
        csr_add_x_425_n177), .SO(csr_n_T_286[3]) );
  AO22X1_LVT csr_add_x_425_U146 ( .A1(io_ptw_pmp_5_addr[3]), .A2(
        csr_add_x_425_n176), .A3(csr_add_x_425_n169), .A4(csr_add_x_425_n170), 
        .Y(csr_n_T_286[4]) );
  AND2X1_LVT csr_add_x_425_U145 ( .A1(csr_add_x_425_n170), .A2(
        io_ptw_pmp_5_addr[3]), .Y(csr_add_x_425_n175) );
  HADDX1_LVT csr_add_x_425_U144 ( .A0(csr_add_x_425_n175), .B0(
        io_ptw_pmp_5_addr[4]), .SO(csr_n_T_286[5]) );
  HADDX1_LVT csr_add_x_425_U143 ( .A0(io_ptw_pmp_5_addr[5]), .B0(
        csr_add_x_425_n174), .SO(csr_n_T_286[6]) );
  AND2X1_LVT csr_add_x_425_U142 ( .A1(io_ptw_pmp_5_addr[5]), .A2(
        csr_add_x_425_n174), .Y(csr_add_x_425_n173) );
  HADDX1_LVT csr_add_x_425_U141 ( .A0(io_ptw_pmp_5_addr[6]), .B0(
        csr_add_x_425_n173), .SO(csr_n_T_286[7]) );
  AO22X1_LVT csr_add_x_425_U140 ( .A1(csr_add_x_425_n168), .A2(
        csr_add_x_425_n167), .A3(csr_add_x_425_n172), .A4(io_ptw_pmp_5_addr[7]), .Y(csr_n_T_286[8]) );
  AND2X1_LVT csr_add_x_425_U139 ( .A1(io_ptw_pmp_5_addr[7]), .A2(
        csr_add_x_425_n168), .Y(csr_add_x_425_n171) );
  HADDX1_LVT csr_add_x_425_U138 ( .A0(csr_add_x_425_n171), .B0(
        io_ptw_pmp_5_addr[8]), .SO(csr_n_T_286[9]) );
  INVX1_LVT csr_add_x_425_U137 ( .A(csr_add_x_425_n176), .Y(csr_add_x_425_n170) );
  INVX1_LVT csr_add_x_425_U136 ( .A(io_ptw_pmp_5_addr[3]), .Y(
        csr_add_x_425_n169) );
  INVX1_LVT csr_add_x_425_U135 ( .A(csr_add_x_425_n172), .Y(csr_add_x_425_n168) );
  INVX1_LVT csr_add_x_425_U134 ( .A(io_ptw_pmp_5_addr[7]), .Y(
        csr_add_x_425_n167) );
  INVX1_LVT csr_add_x_425_U133 ( .A(csr_add_x_425_n196), .Y(csr_add_x_425_n166) );
  INVX1_LVT csr_add_x_425_U132 ( .A(io_ptw_pmp_5_addr[11]), .Y(
        csr_add_x_425_n165) );
  INVX1_LVT csr_add_x_425_U131 ( .A(csr_add_x_425_n192), .Y(csr_add_x_425_n164) );
  INVX1_LVT csr_add_x_425_U130 ( .A(io_ptw_pmp_5_addr[15]), .Y(
        csr_add_x_425_n163) );
  INVX1_LVT csr_add_x_425_U129 ( .A(csr_add_x_425_n187), .Y(csr_add_x_425_n162) );
  INVX1_LVT csr_add_x_425_U128 ( .A(io_ptw_pmp_5_addr[19]), .Y(
        csr_add_x_425_n161) );
  INVX1_LVT csr_add_x_425_U127 ( .A(csr_add_x_425_n183), .Y(csr_add_x_425_n160) );
  INVX1_LVT csr_add_x_425_U126 ( .A(io_ptw_pmp_5_addr[23]), .Y(
        csr_add_x_425_n159) );
  HADDX1_LVT csr_add_x_425_U121 ( .A0(io_ptw_pmp_5_addr[0]), .B0(
        io_ptw_pmp_5_cfg_a[0]), .C1(csr_add_x_425_n93), .SO(csr_n_T_286[1]) );
  NAND3X0_LVT csr_add_x_424_U194 ( .A1(csr_add_x_424_n93), .A2(
        io_ptw_pmp_4_addr[1]), .A3(io_ptw_pmp_4_addr[2]), .Y(
        csr_add_x_424_n176) );
  AND3X1_LVT csr_add_x_424_U193 ( .A1(io_ptw_pmp_4_addr[3]), .A2(
        io_ptw_pmp_4_addr[4]), .A3(csr_add_x_424_n170), .Y(csr_add_x_424_n174)
         );
  NAND3X0_LVT csr_add_x_424_U192 ( .A1(io_ptw_pmp_4_addr[5]), .A2(
        io_ptw_pmp_4_addr[6]), .A3(csr_add_x_424_n174), .Y(csr_add_x_424_n172)
         );
  AND3X1_LVT csr_add_x_424_U191 ( .A1(csr_add_x_424_n168), .A2(
        io_ptw_pmp_4_addr[8]), .A3(io_ptw_pmp_4_addr[7]), .Y(
        csr_add_x_424_n199) );
  HADDX1_LVT csr_add_x_424_U190 ( .A0(io_ptw_pmp_4_addr[9]), .B0(
        csr_add_x_424_n199), .SO(csr_n_T_277[10]) );
  AND4X1_LVT csr_add_x_424_U189 ( .A1(csr_add_x_424_n168), .A2(
        io_ptw_pmp_4_addr[8]), .A3(io_ptw_pmp_4_addr[7]), .A4(
        io_ptw_pmp_4_addr[9]), .Y(csr_add_x_424_n198) );
  HADDX1_LVT csr_add_x_424_U188 ( .A0(io_ptw_pmp_4_addr[10]), .B0(
        csr_add_x_424_n198), .SO(csr_n_T_277[11]) );
  AND4X1_LVT csr_add_x_424_U187 ( .A1(io_ptw_pmp_4_addr[8]), .A2(
        io_ptw_pmp_4_addr[7]), .A3(io_ptw_pmp_4_addr[10]), .A4(
        io_ptw_pmp_4_addr[9]), .Y(csr_add_x_424_n197) );
  NAND2X0_LVT csr_add_x_424_U186 ( .A1(csr_add_x_424_n168), .A2(
        csr_add_x_424_n197), .Y(csr_add_x_424_n196) );
  AO22X1_LVT csr_add_x_424_U185 ( .A1(io_ptw_pmp_4_addr[11]), .A2(
        csr_add_x_424_n196), .A3(csr_add_x_424_n165), .A4(csr_add_x_424_n166), 
        .Y(csr_n_T_277[12]) );
  AND2X1_LVT csr_add_x_424_U184 ( .A1(csr_add_x_424_n166), .A2(
        io_ptw_pmp_4_addr[11]), .Y(csr_add_x_424_n195) );
  HADDX1_LVT csr_add_x_424_U183 ( .A0(csr_add_x_424_n195), .B0(
        io_ptw_pmp_4_addr[12]), .SO(csr_n_T_277[13]) );
  AND3X1_LVT csr_add_x_424_U182 ( .A1(io_ptw_pmp_4_addr[11]), .A2(
        io_ptw_pmp_4_addr[12]), .A3(csr_add_x_424_n166), .Y(csr_add_x_424_n193) );
  HADDX1_LVT csr_add_x_424_U181 ( .A0(io_ptw_pmp_4_addr[13]), .B0(
        csr_add_x_424_n193), .SO(csr_n_T_277[14]) );
  AND4X1_LVT csr_add_x_424_U180 ( .A1(io_ptw_pmp_4_addr[11]), .A2(
        io_ptw_pmp_4_addr[12]), .A3(io_ptw_pmp_4_addr[13]), .A4(
        csr_add_x_424_n166), .Y(csr_add_x_424_n194) );
  HADDX1_LVT csr_add_x_424_U179 ( .A0(io_ptw_pmp_4_addr[14]), .B0(
        csr_add_x_424_n194), .SO(csr_n_T_277[15]) );
  NAND3X0_LVT csr_add_x_424_U178 ( .A1(io_ptw_pmp_4_addr[13]), .A2(
        io_ptw_pmp_4_addr[14]), .A3(csr_add_x_424_n193), .Y(csr_add_x_424_n192) );
  AO22X1_LVT csr_add_x_424_U177 ( .A1(io_ptw_pmp_4_addr[15]), .A2(
        csr_add_x_424_n192), .A3(csr_add_x_424_n163), .A4(csr_add_x_424_n164), 
        .Y(csr_n_T_277[16]) );
  AND2X1_LVT csr_add_x_424_U176 ( .A1(csr_add_x_424_n164), .A2(
        io_ptw_pmp_4_addr[15]), .Y(csr_add_x_424_n191) );
  HADDX1_LVT csr_add_x_424_U175 ( .A0(csr_add_x_424_n191), .B0(
        io_ptw_pmp_4_addr[16]), .SO(csr_n_T_277[17]) );
  AND3X1_LVT csr_add_x_424_U174 ( .A1(io_ptw_pmp_4_addr[15]), .A2(
        io_ptw_pmp_4_addr[16]), .A3(csr_add_x_424_n164), .Y(csr_add_x_424_n190) );
  HADDX1_LVT csr_add_x_424_U173 ( .A0(io_ptw_pmp_4_addr[17]), .B0(
        csr_add_x_424_n190), .SO(csr_n_T_277[18]) );
  AND4X1_LVT csr_add_x_424_U172 ( .A1(io_ptw_pmp_4_addr[15]), .A2(
        io_ptw_pmp_4_addr[16]), .A3(io_ptw_pmp_4_addr[17]), .A4(
        csr_add_x_424_n164), .Y(csr_add_x_424_n189) );
  HADDX1_LVT csr_add_x_424_U171 ( .A0(io_ptw_pmp_4_addr[18]), .B0(
        csr_add_x_424_n189), .SO(csr_n_T_277[19]) );
  AND4X1_LVT csr_add_x_424_U170 ( .A1(io_ptw_pmp_4_addr[15]), .A2(
        io_ptw_pmp_4_addr[16]), .A3(io_ptw_pmp_4_addr[18]), .A4(
        io_ptw_pmp_4_addr[17]), .Y(csr_add_x_424_n188) );
  NAND2X0_LVT csr_add_x_424_U169 ( .A1(csr_add_x_424_n188), .A2(
        csr_add_x_424_n164), .Y(csr_add_x_424_n187) );
  AO22X1_LVT csr_add_x_424_U168 ( .A1(io_ptw_pmp_4_addr[19]), .A2(
        csr_add_x_424_n187), .A3(csr_add_x_424_n161), .A4(csr_add_x_424_n162), 
        .Y(csr_n_T_277[20]) );
  AND2X1_LVT csr_add_x_424_U167 ( .A1(csr_add_x_424_n162), .A2(
        io_ptw_pmp_4_addr[19]), .Y(csr_add_x_424_n186) );
  HADDX1_LVT csr_add_x_424_U166 ( .A0(csr_add_x_424_n186), .B0(
        io_ptw_pmp_4_addr[20]), .SO(csr_n_T_277[21]) );
  AND3X1_LVT csr_add_x_424_U165 ( .A1(io_ptw_pmp_4_addr[19]), .A2(
        io_ptw_pmp_4_addr[20]), .A3(csr_add_x_424_n162), .Y(csr_add_x_424_n184) );
  HADDX1_LVT csr_add_x_424_U164 ( .A0(io_ptw_pmp_4_addr[21]), .B0(
        csr_add_x_424_n184), .SO(csr_n_T_277[22]) );
  AND2X1_LVT csr_add_x_424_U163 ( .A1(csr_add_x_424_n184), .A2(
        io_ptw_pmp_4_addr[21]), .Y(csr_add_x_424_n185) );
  HADDX1_LVT csr_add_x_424_U162 ( .A0(csr_add_x_424_n185), .B0(
        io_ptw_pmp_4_addr[22]), .SO(csr_n_T_277[23]) );
  NAND3X0_LVT csr_add_x_424_U161 ( .A1(io_ptw_pmp_4_addr[22]), .A2(
        io_ptw_pmp_4_addr[21]), .A3(csr_add_x_424_n184), .Y(csr_add_x_424_n183) );
  AO22X1_LVT csr_add_x_424_U160 ( .A1(io_ptw_pmp_4_addr[23]), .A2(
        csr_add_x_424_n183), .A3(csr_add_x_424_n159), .A4(csr_add_x_424_n160), 
        .Y(csr_n_T_277[24]) );
  AND2X1_LVT csr_add_x_424_U159 ( .A1(csr_add_x_424_n160), .A2(
        io_ptw_pmp_4_addr[23]), .Y(csr_add_x_424_n182) );
  HADDX1_LVT csr_add_x_424_U158 ( .A0(csr_add_x_424_n182), .B0(
        io_ptw_pmp_4_addr[24]), .SO(csr_n_T_277[25]) );
  AND3X1_LVT csr_add_x_424_U157 ( .A1(io_ptw_pmp_4_addr[23]), .A2(
        io_ptw_pmp_4_addr[24]), .A3(csr_add_x_424_n160), .Y(csr_add_x_424_n181) );
  HADDX1_LVT csr_add_x_424_U156 ( .A0(io_ptw_pmp_4_addr[25]), .B0(
        csr_add_x_424_n181), .SO(csr_n_T_277[26]) );
  AND2X1_LVT csr_add_x_424_U155 ( .A1(io_ptw_pmp_4_addr[25]), .A2(
        csr_add_x_424_n181), .Y(csr_add_x_424_n179) );
  HADDX1_LVT csr_add_x_424_U154 ( .A0(io_ptw_pmp_4_addr[26]), .B0(
        csr_add_x_424_n179), .SO(csr_n_T_277[27]) );
  AND2X1_LVT csr_add_x_424_U153 ( .A1(io_ptw_pmp_4_addr[26]), .A2(
        csr_add_x_424_n179), .Y(csr_add_x_424_n180) );
  HADDX1_LVT csr_add_x_424_U152 ( .A0(csr_add_x_424_n180), .B0(
        io_ptw_pmp_4_addr[27]), .SO(csr_n_T_277[28]) );
  AND3X1_LVT csr_add_x_424_U151 ( .A1(csr_add_x_424_n179), .A2(
        io_ptw_pmp_4_addr[26]), .A3(io_ptw_pmp_4_addr[27]), .Y(
        csr_add_x_424_n178) );
  HADDX1_LVT csr_add_x_424_U150 ( .A0(csr_add_x_424_n178), .B0(
        io_ptw_pmp_4_addr[28]), .SO(csr_n_T_277[29]) );
  HADDX1_LVT csr_add_x_424_U149 ( .A0(csr_add_x_424_n93), .B0(
        io_ptw_pmp_4_addr[1]), .SO(csr_n_T_277[2]) );
  AND2X1_LVT csr_add_x_424_U148 ( .A1(csr_add_x_424_n93), .A2(
        io_ptw_pmp_4_addr[1]), .Y(csr_add_x_424_n177) );
  HADDX1_LVT csr_add_x_424_U147 ( .A0(io_ptw_pmp_4_addr[2]), .B0(
        csr_add_x_424_n177), .SO(csr_n_T_277[3]) );
  AO22X1_LVT csr_add_x_424_U146 ( .A1(io_ptw_pmp_4_addr[3]), .A2(
        csr_add_x_424_n176), .A3(csr_add_x_424_n169), .A4(csr_add_x_424_n170), 
        .Y(csr_n_T_277[4]) );
  AND2X1_LVT csr_add_x_424_U145 ( .A1(csr_add_x_424_n170), .A2(
        io_ptw_pmp_4_addr[3]), .Y(csr_add_x_424_n175) );
  HADDX1_LVT csr_add_x_424_U144 ( .A0(csr_add_x_424_n175), .B0(
        io_ptw_pmp_4_addr[4]), .SO(csr_n_T_277[5]) );
  HADDX1_LVT csr_add_x_424_U143 ( .A0(io_ptw_pmp_4_addr[5]), .B0(
        csr_add_x_424_n174), .SO(csr_n_T_277[6]) );
  AND2X1_LVT csr_add_x_424_U142 ( .A1(io_ptw_pmp_4_addr[5]), .A2(
        csr_add_x_424_n174), .Y(csr_add_x_424_n173) );
  HADDX1_LVT csr_add_x_424_U141 ( .A0(io_ptw_pmp_4_addr[6]), .B0(
        csr_add_x_424_n173), .SO(csr_n_T_277[7]) );
  AO22X1_LVT csr_add_x_424_U140 ( .A1(csr_add_x_424_n168), .A2(
        csr_add_x_424_n167), .A3(csr_add_x_424_n172), .A4(io_ptw_pmp_4_addr[7]), .Y(csr_n_T_277[8]) );
  AND2X1_LVT csr_add_x_424_U139 ( .A1(io_ptw_pmp_4_addr[7]), .A2(
        csr_add_x_424_n168), .Y(csr_add_x_424_n171) );
  HADDX1_LVT csr_add_x_424_U138 ( .A0(csr_add_x_424_n171), .B0(
        io_ptw_pmp_4_addr[8]), .SO(csr_n_T_277[9]) );
  INVX1_LVT csr_add_x_424_U137 ( .A(csr_add_x_424_n176), .Y(csr_add_x_424_n170) );
  INVX1_LVT csr_add_x_424_U136 ( .A(io_ptw_pmp_4_addr[3]), .Y(
        csr_add_x_424_n169) );
  INVX1_LVT csr_add_x_424_U135 ( .A(csr_add_x_424_n172), .Y(csr_add_x_424_n168) );
  INVX1_LVT csr_add_x_424_U134 ( .A(io_ptw_pmp_4_addr[7]), .Y(
        csr_add_x_424_n167) );
  INVX1_LVT csr_add_x_424_U133 ( .A(csr_add_x_424_n196), .Y(csr_add_x_424_n166) );
  INVX1_LVT csr_add_x_424_U132 ( .A(io_ptw_pmp_4_addr[11]), .Y(
        csr_add_x_424_n165) );
  INVX1_LVT csr_add_x_424_U131 ( .A(csr_add_x_424_n192), .Y(csr_add_x_424_n164) );
  INVX1_LVT csr_add_x_424_U130 ( .A(io_ptw_pmp_4_addr[15]), .Y(
        csr_add_x_424_n163) );
  INVX1_LVT csr_add_x_424_U129 ( .A(csr_add_x_424_n187), .Y(csr_add_x_424_n162) );
  INVX1_LVT csr_add_x_424_U128 ( .A(io_ptw_pmp_4_addr[19]), .Y(
        csr_add_x_424_n161) );
  INVX1_LVT csr_add_x_424_U127 ( .A(csr_add_x_424_n183), .Y(csr_add_x_424_n160) );
  INVX1_LVT csr_add_x_424_U126 ( .A(io_ptw_pmp_4_addr[23]), .Y(
        csr_add_x_424_n159) );
  HADDX1_LVT csr_add_x_424_U121 ( .A0(io_ptw_pmp_4_addr[0]), .B0(
        io_ptw_pmp_4_cfg_a[0]), .C1(csr_add_x_424_n93), .SO(csr_n_T_277[1]) );
  NAND3X0_LVT csr_add_x_423_U194 ( .A1(csr_add_x_423_n93), .A2(
        io_ptw_pmp_3_addr[1]), .A3(io_ptw_pmp_3_addr[2]), .Y(
        csr_add_x_423_n176) );
  AND3X1_LVT csr_add_x_423_U193 ( .A1(io_ptw_pmp_3_addr[3]), .A2(
        io_ptw_pmp_3_addr[4]), .A3(csr_add_x_423_n164), .Y(csr_add_x_423_n174)
         );
  NAND3X0_LVT csr_add_x_423_U192 ( .A1(io_ptw_pmp_3_addr[5]), .A2(
        io_ptw_pmp_3_addr[6]), .A3(csr_add_x_423_n174), .Y(csr_add_x_423_n172)
         );
  AND3X1_LVT csr_add_x_423_U191 ( .A1(csr_add_x_423_n163), .A2(
        io_ptw_pmp_3_addr[8]), .A3(io_ptw_pmp_3_addr[7]), .Y(
        csr_add_x_423_n199) );
  HADDX1_LVT csr_add_x_423_U190 ( .A0(io_ptw_pmp_3_addr[9]), .B0(
        csr_add_x_423_n199), .SO(csr_n_T_268[10]) );
  AND4X1_LVT csr_add_x_423_U189 ( .A1(csr_add_x_423_n163), .A2(
        io_ptw_pmp_3_addr[8]), .A3(io_ptw_pmp_3_addr[7]), .A4(
        io_ptw_pmp_3_addr[9]), .Y(csr_add_x_423_n198) );
  HADDX1_LVT csr_add_x_423_U188 ( .A0(io_ptw_pmp_3_addr[10]), .B0(
        csr_add_x_423_n198), .SO(csr_n_T_268[11]) );
  AND4X1_LVT csr_add_x_423_U187 ( .A1(io_ptw_pmp_3_addr[8]), .A2(
        io_ptw_pmp_3_addr[7]), .A3(io_ptw_pmp_3_addr[10]), .A4(
        io_ptw_pmp_3_addr[9]), .Y(csr_add_x_423_n197) );
  NAND2X0_LVT csr_add_x_423_U186 ( .A1(csr_add_x_423_n163), .A2(
        csr_add_x_423_n197), .Y(csr_add_x_423_n196) );
  AO22X1_LVT csr_add_x_423_U185 ( .A1(io_ptw_pmp_3_addr[11]), .A2(
        csr_add_x_423_n196), .A3(csr_add_x_423_n168), .A4(csr_add_x_423_n162), 
        .Y(csr_n_T_268[12]) );
  AND2X1_LVT csr_add_x_423_U184 ( .A1(csr_add_x_423_n162), .A2(
        io_ptw_pmp_3_addr[11]), .Y(csr_add_x_423_n195) );
  HADDX1_LVT csr_add_x_423_U183 ( .A0(csr_add_x_423_n195), .B0(
        io_ptw_pmp_3_addr[12]), .SO(csr_n_T_268[13]) );
  AND3X1_LVT csr_add_x_423_U182 ( .A1(io_ptw_pmp_3_addr[11]), .A2(
        io_ptw_pmp_3_addr[12]), .A3(csr_add_x_423_n162), .Y(csr_add_x_423_n193) );
  HADDX1_LVT csr_add_x_423_U181 ( .A0(io_ptw_pmp_3_addr[13]), .B0(
        csr_add_x_423_n193), .SO(csr_n_T_268[14]) );
  AND4X1_LVT csr_add_x_423_U180 ( .A1(io_ptw_pmp_3_addr[11]), .A2(
        io_ptw_pmp_3_addr[12]), .A3(io_ptw_pmp_3_addr[13]), .A4(
        csr_add_x_423_n162), .Y(csr_add_x_423_n194) );
  HADDX1_LVT csr_add_x_423_U179 ( .A0(io_ptw_pmp_3_addr[14]), .B0(
        csr_add_x_423_n194), .SO(csr_n_T_268[15]) );
  NAND3X0_LVT csr_add_x_423_U178 ( .A1(io_ptw_pmp_3_addr[13]), .A2(
        io_ptw_pmp_3_addr[14]), .A3(csr_add_x_423_n193), .Y(csr_add_x_423_n192) );
  AO22X1_LVT csr_add_x_423_U177 ( .A1(io_ptw_pmp_3_addr[15]), .A2(
        csr_add_x_423_n192), .A3(csr_add_x_423_n167), .A4(csr_add_x_423_n161), 
        .Y(csr_n_T_268[16]) );
  AND2X1_LVT csr_add_x_423_U176 ( .A1(csr_add_x_423_n161), .A2(
        io_ptw_pmp_3_addr[15]), .Y(csr_add_x_423_n191) );
  HADDX1_LVT csr_add_x_423_U175 ( .A0(csr_add_x_423_n191), .B0(
        io_ptw_pmp_3_addr[16]), .SO(csr_n_T_268[17]) );
  AND3X1_LVT csr_add_x_423_U174 ( .A1(io_ptw_pmp_3_addr[15]), .A2(
        io_ptw_pmp_3_addr[16]), .A3(csr_add_x_423_n161), .Y(csr_add_x_423_n190) );
  HADDX1_LVT csr_add_x_423_U173 ( .A0(io_ptw_pmp_3_addr[17]), .B0(
        csr_add_x_423_n190), .SO(csr_n_T_268[18]) );
  AND4X1_LVT csr_add_x_423_U172 ( .A1(io_ptw_pmp_3_addr[15]), .A2(
        io_ptw_pmp_3_addr[16]), .A3(io_ptw_pmp_3_addr[17]), .A4(
        csr_add_x_423_n161), .Y(csr_add_x_423_n189) );
  HADDX1_LVT csr_add_x_423_U171 ( .A0(io_ptw_pmp_3_addr[18]), .B0(
        csr_add_x_423_n189), .SO(csr_n_T_268[19]) );
  AND4X1_LVT csr_add_x_423_U170 ( .A1(io_ptw_pmp_3_addr[15]), .A2(
        io_ptw_pmp_3_addr[16]), .A3(io_ptw_pmp_3_addr[18]), .A4(
        io_ptw_pmp_3_addr[17]), .Y(csr_add_x_423_n188) );
  NAND2X0_LVT csr_add_x_423_U169 ( .A1(csr_add_x_423_n188), .A2(
        csr_add_x_423_n161), .Y(csr_add_x_423_n187) );
  AO22X1_LVT csr_add_x_423_U168 ( .A1(io_ptw_pmp_3_addr[19]), .A2(
        csr_add_x_423_n187), .A3(csr_add_x_423_n166), .A4(csr_add_x_423_n160), 
        .Y(csr_n_T_268[20]) );
  AND2X1_LVT csr_add_x_423_U167 ( .A1(csr_add_x_423_n160), .A2(
        io_ptw_pmp_3_addr[19]), .Y(csr_add_x_423_n186) );
  HADDX1_LVT csr_add_x_423_U166 ( .A0(csr_add_x_423_n186), .B0(
        io_ptw_pmp_3_addr[20]), .SO(csr_n_T_268[21]) );
  AND3X1_LVT csr_add_x_423_U165 ( .A1(io_ptw_pmp_3_addr[19]), .A2(
        io_ptw_pmp_3_addr[20]), .A3(csr_add_x_423_n160), .Y(csr_add_x_423_n184) );
  HADDX1_LVT csr_add_x_423_U164 ( .A0(io_ptw_pmp_3_addr[21]), .B0(
        csr_add_x_423_n184), .SO(csr_n_T_268[22]) );
  AND2X1_LVT csr_add_x_423_U163 ( .A1(csr_add_x_423_n184), .A2(
        io_ptw_pmp_3_addr[21]), .Y(csr_add_x_423_n185) );
  HADDX1_LVT csr_add_x_423_U162 ( .A0(csr_add_x_423_n185), .B0(
        io_ptw_pmp_3_addr[22]), .SO(csr_n_T_268[23]) );
  NAND3X0_LVT csr_add_x_423_U161 ( .A1(io_ptw_pmp_3_addr[22]), .A2(
        io_ptw_pmp_3_addr[21]), .A3(csr_add_x_423_n184), .Y(csr_add_x_423_n183) );
  AO22X1_LVT csr_add_x_423_U160 ( .A1(io_ptw_pmp_3_addr[23]), .A2(
        csr_add_x_423_n183), .A3(csr_add_x_423_n165), .A4(csr_add_x_423_n159), 
        .Y(csr_n_T_268[24]) );
  AND2X1_LVT csr_add_x_423_U159 ( .A1(csr_add_x_423_n159), .A2(
        io_ptw_pmp_3_addr[23]), .Y(csr_add_x_423_n182) );
  HADDX1_LVT csr_add_x_423_U158 ( .A0(csr_add_x_423_n182), .B0(
        io_ptw_pmp_3_addr[24]), .SO(csr_n_T_268[25]) );
  AND3X1_LVT csr_add_x_423_U157 ( .A1(io_ptw_pmp_3_addr[23]), .A2(
        io_ptw_pmp_3_addr[24]), .A3(csr_add_x_423_n159), .Y(csr_add_x_423_n181) );
  HADDX1_LVT csr_add_x_423_U156 ( .A0(io_ptw_pmp_3_addr[25]), .B0(
        csr_add_x_423_n181), .SO(csr_n_T_268[26]) );
  AND2X1_LVT csr_add_x_423_U155 ( .A1(io_ptw_pmp_3_addr[25]), .A2(
        csr_add_x_423_n181), .Y(csr_add_x_423_n179) );
  HADDX1_LVT csr_add_x_423_U154 ( .A0(io_ptw_pmp_3_addr[26]), .B0(
        csr_add_x_423_n179), .SO(csr_n_T_268[27]) );
  AND2X1_LVT csr_add_x_423_U153 ( .A1(io_ptw_pmp_3_addr[26]), .A2(
        csr_add_x_423_n179), .Y(csr_add_x_423_n180) );
  HADDX1_LVT csr_add_x_423_U152 ( .A0(csr_add_x_423_n180), .B0(
        io_ptw_pmp_3_addr[27]), .SO(csr_n_T_268[28]) );
  AND3X1_LVT csr_add_x_423_U151 ( .A1(csr_add_x_423_n179), .A2(
        io_ptw_pmp_3_addr[26]), .A3(io_ptw_pmp_3_addr[27]), .Y(
        csr_add_x_423_n178) );
  HADDX1_LVT csr_add_x_423_U150 ( .A0(csr_add_x_423_n178), .B0(
        io_ptw_pmp_3_addr[28]), .SO(csr_n_T_268[29]) );
  HADDX1_LVT csr_add_x_423_U149 ( .A0(csr_add_x_423_n93), .B0(
        io_ptw_pmp_3_addr[1]), .SO(csr_n_T_268[2]) );
  AND2X1_LVT csr_add_x_423_U148 ( .A1(csr_add_x_423_n93), .A2(
        io_ptw_pmp_3_addr[1]), .Y(csr_add_x_423_n177) );
  HADDX1_LVT csr_add_x_423_U147 ( .A0(io_ptw_pmp_3_addr[2]), .B0(
        csr_add_x_423_n177), .SO(csr_n_T_268[3]) );
  AO22X1_LVT csr_add_x_423_U146 ( .A1(io_ptw_pmp_3_addr[3]), .A2(
        csr_add_x_423_n176), .A3(csr_add_x_423_n170), .A4(csr_add_x_423_n164), 
        .Y(csr_n_T_268[4]) );
  AND2X1_LVT csr_add_x_423_U145 ( .A1(csr_add_x_423_n164), .A2(
        io_ptw_pmp_3_addr[3]), .Y(csr_add_x_423_n175) );
  HADDX1_LVT csr_add_x_423_U144 ( .A0(csr_add_x_423_n175), .B0(
        io_ptw_pmp_3_addr[4]), .SO(csr_n_T_268[5]) );
  HADDX1_LVT csr_add_x_423_U143 ( .A0(io_ptw_pmp_3_addr[5]), .B0(
        csr_add_x_423_n174), .SO(csr_n_T_268[6]) );
  AND2X1_LVT csr_add_x_423_U142 ( .A1(io_ptw_pmp_3_addr[5]), .A2(
        csr_add_x_423_n174), .Y(csr_add_x_423_n173) );
  HADDX1_LVT csr_add_x_423_U141 ( .A0(io_ptw_pmp_3_addr[6]), .B0(
        csr_add_x_423_n173), .SO(csr_n_T_268[7]) );
  AO22X1_LVT csr_add_x_423_U140 ( .A1(csr_add_x_423_n163), .A2(
        csr_add_x_423_n169), .A3(csr_add_x_423_n172), .A4(io_ptw_pmp_3_addr[7]), .Y(csr_n_T_268[8]) );
  AND2X1_LVT csr_add_x_423_U139 ( .A1(io_ptw_pmp_3_addr[7]), .A2(
        csr_add_x_423_n163), .Y(csr_add_x_423_n171) );
  HADDX1_LVT csr_add_x_423_U138 ( .A0(csr_add_x_423_n171), .B0(
        io_ptw_pmp_3_addr[8]), .SO(csr_n_T_268[9]) );
  INVX1_LVT csr_add_x_423_U137 ( .A(io_ptw_pmp_3_addr[3]), .Y(
        csr_add_x_423_n170) );
  INVX1_LVT csr_add_x_423_U136 ( .A(io_ptw_pmp_3_addr[7]), .Y(
        csr_add_x_423_n169) );
  INVX1_LVT csr_add_x_423_U135 ( .A(io_ptw_pmp_3_addr[11]), .Y(
        csr_add_x_423_n168) );
  INVX1_LVT csr_add_x_423_U134 ( .A(io_ptw_pmp_3_addr[15]), .Y(
        csr_add_x_423_n167) );
  INVX1_LVT csr_add_x_423_U133 ( .A(io_ptw_pmp_3_addr[19]), .Y(
        csr_add_x_423_n166) );
  INVX1_LVT csr_add_x_423_U132 ( .A(io_ptw_pmp_3_addr[23]), .Y(
        csr_add_x_423_n165) );
  INVX1_LVT csr_add_x_423_U131 ( .A(csr_add_x_423_n176), .Y(csr_add_x_423_n164) );
  INVX1_LVT csr_add_x_423_U130 ( .A(csr_add_x_423_n172), .Y(csr_add_x_423_n163) );
  INVX1_LVT csr_add_x_423_U129 ( .A(csr_add_x_423_n196), .Y(csr_add_x_423_n162) );
  INVX1_LVT csr_add_x_423_U128 ( .A(csr_add_x_423_n192), .Y(csr_add_x_423_n161) );
  INVX1_LVT csr_add_x_423_U127 ( .A(csr_add_x_423_n187), .Y(csr_add_x_423_n160) );
  INVX1_LVT csr_add_x_423_U126 ( .A(csr_add_x_423_n183), .Y(csr_add_x_423_n159) );
  HADDX1_LVT csr_add_x_423_U121 ( .A0(io_ptw_pmp_3_addr[0]), .B0(
        io_ptw_pmp_3_cfg_a[0]), .C1(csr_add_x_423_n93), .SO(csr_n_T_268[1]) );
  NAND3X0_LVT csr_add_x_422_U194 ( .A1(csr_add_x_422_n93), .A2(
        io_ptw_pmp_2_addr[1]), .A3(io_ptw_pmp_2_addr[2]), .Y(
        csr_add_x_422_n176) );
  AND3X1_LVT csr_add_x_422_U193 ( .A1(io_ptw_pmp_2_addr[3]), .A2(
        io_ptw_pmp_2_addr[4]), .A3(csr_add_x_422_n164), .Y(csr_add_x_422_n174)
         );
  NAND3X0_LVT csr_add_x_422_U192 ( .A1(io_ptw_pmp_2_addr[5]), .A2(
        io_ptw_pmp_2_addr[6]), .A3(csr_add_x_422_n174), .Y(csr_add_x_422_n172)
         );
  AND3X1_LVT csr_add_x_422_U191 ( .A1(csr_add_x_422_n163), .A2(
        io_ptw_pmp_2_addr[8]), .A3(io_ptw_pmp_2_addr[7]), .Y(
        csr_add_x_422_n199) );
  HADDX1_LVT csr_add_x_422_U190 ( .A0(io_ptw_pmp_2_addr[9]), .B0(
        csr_add_x_422_n199), .SO(csr_n_T_259[10]) );
  AND4X1_LVT csr_add_x_422_U189 ( .A1(csr_add_x_422_n163), .A2(
        io_ptw_pmp_2_addr[8]), .A3(io_ptw_pmp_2_addr[7]), .A4(
        io_ptw_pmp_2_addr[9]), .Y(csr_add_x_422_n198) );
  HADDX1_LVT csr_add_x_422_U188 ( .A0(io_ptw_pmp_2_addr[10]), .B0(
        csr_add_x_422_n198), .SO(csr_n_T_259[11]) );
  AND4X1_LVT csr_add_x_422_U187 ( .A1(io_ptw_pmp_2_addr[8]), .A2(
        io_ptw_pmp_2_addr[7]), .A3(io_ptw_pmp_2_addr[10]), .A4(
        io_ptw_pmp_2_addr[9]), .Y(csr_add_x_422_n197) );
  NAND2X0_LVT csr_add_x_422_U186 ( .A1(csr_add_x_422_n163), .A2(
        csr_add_x_422_n197), .Y(csr_add_x_422_n196) );
  AO22X1_LVT csr_add_x_422_U185 ( .A1(io_ptw_pmp_2_addr[11]), .A2(
        csr_add_x_422_n196), .A3(csr_add_x_422_n168), .A4(csr_add_x_422_n162), 
        .Y(csr_n_T_259[12]) );
  AND2X1_LVT csr_add_x_422_U184 ( .A1(csr_add_x_422_n162), .A2(
        io_ptw_pmp_2_addr[11]), .Y(csr_add_x_422_n195) );
  HADDX1_LVT csr_add_x_422_U183 ( .A0(csr_add_x_422_n195), .B0(
        io_ptw_pmp_2_addr[12]), .SO(csr_n_T_259[13]) );
  AND3X1_LVT csr_add_x_422_U182 ( .A1(io_ptw_pmp_2_addr[11]), .A2(
        io_ptw_pmp_2_addr[12]), .A3(csr_add_x_422_n162), .Y(csr_add_x_422_n193) );
  HADDX1_LVT csr_add_x_422_U181 ( .A0(io_ptw_pmp_2_addr[13]), .B0(
        csr_add_x_422_n193), .SO(csr_n_T_259[14]) );
  AND4X1_LVT csr_add_x_422_U180 ( .A1(io_ptw_pmp_2_addr[11]), .A2(
        io_ptw_pmp_2_addr[12]), .A3(io_ptw_pmp_2_addr[13]), .A4(
        csr_add_x_422_n162), .Y(csr_add_x_422_n194) );
  HADDX1_LVT csr_add_x_422_U179 ( .A0(io_ptw_pmp_2_addr[14]), .B0(
        csr_add_x_422_n194), .SO(csr_n_T_259[15]) );
  NAND3X0_LVT csr_add_x_422_U178 ( .A1(io_ptw_pmp_2_addr[13]), .A2(
        io_ptw_pmp_2_addr[14]), .A3(csr_add_x_422_n193), .Y(csr_add_x_422_n192) );
  AO22X1_LVT csr_add_x_422_U177 ( .A1(io_ptw_pmp_2_addr[15]), .A2(
        csr_add_x_422_n192), .A3(csr_add_x_422_n167), .A4(csr_add_x_422_n161), 
        .Y(csr_n_T_259[16]) );
  AND2X1_LVT csr_add_x_422_U176 ( .A1(csr_add_x_422_n161), .A2(
        io_ptw_pmp_2_addr[15]), .Y(csr_add_x_422_n191) );
  HADDX1_LVT csr_add_x_422_U175 ( .A0(csr_add_x_422_n191), .B0(
        io_ptw_pmp_2_addr[16]), .SO(csr_n_T_259[17]) );
  AND3X1_LVT csr_add_x_422_U174 ( .A1(io_ptw_pmp_2_addr[15]), .A2(
        io_ptw_pmp_2_addr[16]), .A3(csr_add_x_422_n161), .Y(csr_add_x_422_n190) );
  HADDX1_LVT csr_add_x_422_U173 ( .A0(io_ptw_pmp_2_addr[17]), .B0(
        csr_add_x_422_n190), .SO(csr_n_T_259[18]) );
  AND4X1_LVT csr_add_x_422_U172 ( .A1(io_ptw_pmp_2_addr[15]), .A2(
        io_ptw_pmp_2_addr[16]), .A3(io_ptw_pmp_2_addr[17]), .A4(
        csr_add_x_422_n161), .Y(csr_add_x_422_n189) );
  HADDX1_LVT csr_add_x_422_U171 ( .A0(io_ptw_pmp_2_addr[18]), .B0(
        csr_add_x_422_n189), .SO(csr_n_T_259[19]) );
  AND4X1_LVT csr_add_x_422_U170 ( .A1(io_ptw_pmp_2_addr[15]), .A2(
        io_ptw_pmp_2_addr[16]), .A3(io_ptw_pmp_2_addr[18]), .A4(
        io_ptw_pmp_2_addr[17]), .Y(csr_add_x_422_n188) );
  NAND2X0_LVT csr_add_x_422_U169 ( .A1(csr_add_x_422_n188), .A2(
        csr_add_x_422_n161), .Y(csr_add_x_422_n187) );
  AO22X1_LVT csr_add_x_422_U168 ( .A1(io_ptw_pmp_2_addr[19]), .A2(
        csr_add_x_422_n187), .A3(csr_add_x_422_n166), .A4(csr_add_x_422_n160), 
        .Y(csr_n_T_259[20]) );
  AND2X1_LVT csr_add_x_422_U167 ( .A1(csr_add_x_422_n160), .A2(
        io_ptw_pmp_2_addr[19]), .Y(csr_add_x_422_n186) );
  HADDX1_LVT csr_add_x_422_U166 ( .A0(csr_add_x_422_n186), .B0(
        io_ptw_pmp_2_addr[20]), .SO(csr_n_T_259[21]) );
  AND3X1_LVT csr_add_x_422_U165 ( .A1(io_ptw_pmp_2_addr[19]), .A2(
        io_ptw_pmp_2_addr[20]), .A3(csr_add_x_422_n160), .Y(csr_add_x_422_n184) );
  HADDX1_LVT csr_add_x_422_U164 ( .A0(io_ptw_pmp_2_addr[21]), .B0(
        csr_add_x_422_n184), .SO(csr_n_T_259[22]) );
  AND2X1_LVT csr_add_x_422_U163 ( .A1(csr_add_x_422_n184), .A2(
        io_ptw_pmp_2_addr[21]), .Y(csr_add_x_422_n185) );
  HADDX1_LVT csr_add_x_422_U162 ( .A0(csr_add_x_422_n185), .B0(
        io_ptw_pmp_2_addr[22]), .SO(csr_n_T_259[23]) );
  NAND3X0_LVT csr_add_x_422_U161 ( .A1(io_ptw_pmp_2_addr[22]), .A2(
        io_ptw_pmp_2_addr[21]), .A3(csr_add_x_422_n184), .Y(csr_add_x_422_n183) );
  AO22X1_LVT csr_add_x_422_U160 ( .A1(io_ptw_pmp_2_addr[23]), .A2(
        csr_add_x_422_n183), .A3(csr_add_x_422_n165), .A4(csr_add_x_422_n159), 
        .Y(csr_n_T_259[24]) );
  AND2X1_LVT csr_add_x_422_U159 ( .A1(csr_add_x_422_n159), .A2(
        io_ptw_pmp_2_addr[23]), .Y(csr_add_x_422_n182) );
  HADDX1_LVT csr_add_x_422_U158 ( .A0(csr_add_x_422_n182), .B0(
        io_ptw_pmp_2_addr[24]), .SO(csr_n_T_259[25]) );
  AND3X1_LVT csr_add_x_422_U157 ( .A1(io_ptw_pmp_2_addr[23]), .A2(
        io_ptw_pmp_2_addr[24]), .A3(csr_add_x_422_n159), .Y(csr_add_x_422_n181) );
  HADDX1_LVT csr_add_x_422_U156 ( .A0(io_ptw_pmp_2_addr[25]), .B0(
        csr_add_x_422_n181), .SO(csr_n_T_259[26]) );
  AND2X1_LVT csr_add_x_422_U155 ( .A1(io_ptw_pmp_2_addr[25]), .A2(
        csr_add_x_422_n181), .Y(csr_add_x_422_n179) );
  HADDX1_LVT csr_add_x_422_U154 ( .A0(io_ptw_pmp_2_addr[26]), .B0(
        csr_add_x_422_n179), .SO(csr_n_T_259[27]) );
  AND2X1_LVT csr_add_x_422_U153 ( .A1(io_ptw_pmp_2_addr[26]), .A2(
        csr_add_x_422_n179), .Y(csr_add_x_422_n180) );
  HADDX1_LVT csr_add_x_422_U152 ( .A0(csr_add_x_422_n180), .B0(
        io_ptw_pmp_2_addr[27]), .SO(csr_n_T_259[28]) );
  AND3X1_LVT csr_add_x_422_U151 ( .A1(csr_add_x_422_n179), .A2(
        io_ptw_pmp_2_addr[26]), .A3(io_ptw_pmp_2_addr[27]), .Y(
        csr_add_x_422_n178) );
  HADDX1_LVT csr_add_x_422_U150 ( .A0(csr_add_x_422_n178), .B0(
        io_ptw_pmp_2_addr[28]), .SO(csr_n_T_259[29]) );
  HADDX1_LVT csr_add_x_422_U149 ( .A0(csr_add_x_422_n93), .B0(
        io_ptw_pmp_2_addr[1]), .SO(csr_n_T_259[2]) );
  AND2X1_LVT csr_add_x_422_U148 ( .A1(csr_add_x_422_n93), .A2(
        io_ptw_pmp_2_addr[1]), .Y(csr_add_x_422_n177) );
  HADDX1_LVT csr_add_x_422_U147 ( .A0(io_ptw_pmp_2_addr[2]), .B0(
        csr_add_x_422_n177), .SO(csr_n_T_259[3]) );
  AO22X1_LVT csr_add_x_422_U146 ( .A1(io_ptw_pmp_2_addr[3]), .A2(
        csr_add_x_422_n176), .A3(csr_add_x_422_n170), .A4(csr_add_x_422_n164), 
        .Y(csr_n_T_259[4]) );
  AND2X1_LVT csr_add_x_422_U145 ( .A1(csr_add_x_422_n164), .A2(
        io_ptw_pmp_2_addr[3]), .Y(csr_add_x_422_n175) );
  HADDX1_LVT csr_add_x_422_U144 ( .A0(csr_add_x_422_n175), .B0(
        io_ptw_pmp_2_addr[4]), .SO(csr_n_T_259[5]) );
  HADDX1_LVT csr_add_x_422_U143 ( .A0(io_ptw_pmp_2_addr[5]), .B0(
        csr_add_x_422_n174), .SO(csr_n_T_259[6]) );
  AND2X1_LVT csr_add_x_422_U142 ( .A1(io_ptw_pmp_2_addr[5]), .A2(
        csr_add_x_422_n174), .Y(csr_add_x_422_n173) );
  HADDX1_LVT csr_add_x_422_U141 ( .A0(io_ptw_pmp_2_addr[6]), .B0(
        csr_add_x_422_n173), .SO(csr_n_T_259[7]) );
  AO22X1_LVT csr_add_x_422_U140 ( .A1(csr_add_x_422_n163), .A2(
        csr_add_x_422_n169), .A3(csr_add_x_422_n172), .A4(io_ptw_pmp_2_addr[7]), .Y(csr_n_T_259[8]) );
  AND2X1_LVT csr_add_x_422_U139 ( .A1(io_ptw_pmp_2_addr[7]), .A2(
        csr_add_x_422_n163), .Y(csr_add_x_422_n171) );
  HADDX1_LVT csr_add_x_422_U138 ( .A0(csr_add_x_422_n171), .B0(
        io_ptw_pmp_2_addr[8]), .SO(csr_n_T_259[9]) );
  INVX1_LVT csr_add_x_422_U137 ( .A(io_ptw_pmp_2_addr[3]), .Y(
        csr_add_x_422_n170) );
  INVX1_LVT csr_add_x_422_U136 ( .A(io_ptw_pmp_2_addr[7]), .Y(
        csr_add_x_422_n169) );
  INVX1_LVT csr_add_x_422_U135 ( .A(io_ptw_pmp_2_addr[11]), .Y(
        csr_add_x_422_n168) );
  INVX1_LVT csr_add_x_422_U134 ( .A(io_ptw_pmp_2_addr[15]), .Y(
        csr_add_x_422_n167) );
  INVX1_LVT csr_add_x_422_U133 ( .A(io_ptw_pmp_2_addr[19]), .Y(
        csr_add_x_422_n166) );
  INVX1_LVT csr_add_x_422_U132 ( .A(io_ptw_pmp_2_addr[23]), .Y(
        csr_add_x_422_n165) );
  INVX1_LVT csr_add_x_422_U131 ( .A(csr_add_x_422_n176), .Y(csr_add_x_422_n164) );
  INVX1_LVT csr_add_x_422_U130 ( .A(csr_add_x_422_n172), .Y(csr_add_x_422_n163) );
  INVX1_LVT csr_add_x_422_U129 ( .A(csr_add_x_422_n196), .Y(csr_add_x_422_n162) );
  INVX1_LVT csr_add_x_422_U128 ( .A(csr_add_x_422_n192), .Y(csr_add_x_422_n161) );
  INVX1_LVT csr_add_x_422_U127 ( .A(csr_add_x_422_n187), .Y(csr_add_x_422_n160) );
  INVX1_LVT csr_add_x_422_U126 ( .A(csr_add_x_422_n183), .Y(csr_add_x_422_n159) );
  HADDX1_LVT csr_add_x_422_U121 ( .A0(io_ptw_pmp_2_addr[0]), .B0(
        io_ptw_pmp_2_cfg_a[0]), .C1(csr_add_x_422_n93), .SO(csr_n_T_259[1]) );
  NAND3X0_LVT csr_add_x_421_U194 ( .A1(csr_add_x_421_n93), .A2(
        io_ptw_pmp_1_addr[1]), .A3(io_ptw_pmp_1_addr[2]), .Y(
        csr_add_x_421_n176) );
  AND3X1_LVT csr_add_x_421_U193 ( .A1(io_ptw_pmp_1_addr[3]), .A2(
        io_ptw_pmp_1_addr[4]), .A3(csr_add_x_421_n170), .Y(csr_add_x_421_n174)
         );
  NAND3X0_LVT csr_add_x_421_U192 ( .A1(io_ptw_pmp_1_addr[5]), .A2(
        io_ptw_pmp_1_addr[6]), .A3(csr_add_x_421_n174), .Y(csr_add_x_421_n172)
         );
  AND3X1_LVT csr_add_x_421_U191 ( .A1(csr_add_x_421_n168), .A2(
        io_ptw_pmp_1_addr[8]), .A3(io_ptw_pmp_1_addr[7]), .Y(
        csr_add_x_421_n199) );
  HADDX1_LVT csr_add_x_421_U190 ( .A0(io_ptw_pmp_1_addr[9]), .B0(
        csr_add_x_421_n199), .SO(csr_n_T_250[10]) );
  AND4X1_LVT csr_add_x_421_U189 ( .A1(csr_add_x_421_n168), .A2(
        io_ptw_pmp_1_addr[8]), .A3(io_ptw_pmp_1_addr[7]), .A4(
        io_ptw_pmp_1_addr[9]), .Y(csr_add_x_421_n198) );
  HADDX1_LVT csr_add_x_421_U188 ( .A0(io_ptw_pmp_1_addr[10]), .B0(
        csr_add_x_421_n198), .SO(csr_n_T_250[11]) );
  AND4X1_LVT csr_add_x_421_U187 ( .A1(io_ptw_pmp_1_addr[8]), .A2(
        io_ptw_pmp_1_addr[7]), .A3(io_ptw_pmp_1_addr[10]), .A4(
        io_ptw_pmp_1_addr[9]), .Y(csr_add_x_421_n197) );
  NAND2X0_LVT csr_add_x_421_U186 ( .A1(csr_add_x_421_n168), .A2(
        csr_add_x_421_n197), .Y(csr_add_x_421_n196) );
  AO22X1_LVT csr_add_x_421_U185 ( .A1(io_ptw_pmp_1_addr[11]), .A2(
        csr_add_x_421_n196), .A3(csr_add_x_421_n165), .A4(csr_add_x_421_n166), 
        .Y(csr_n_T_250[12]) );
  AND2X1_LVT csr_add_x_421_U184 ( .A1(csr_add_x_421_n166), .A2(
        io_ptw_pmp_1_addr[11]), .Y(csr_add_x_421_n195) );
  HADDX1_LVT csr_add_x_421_U183 ( .A0(csr_add_x_421_n195), .B0(
        io_ptw_pmp_1_addr[12]), .SO(csr_n_T_250[13]) );
  AND3X1_LVT csr_add_x_421_U182 ( .A1(io_ptw_pmp_1_addr[11]), .A2(
        io_ptw_pmp_1_addr[12]), .A3(csr_add_x_421_n166), .Y(csr_add_x_421_n193) );
  HADDX1_LVT csr_add_x_421_U181 ( .A0(io_ptw_pmp_1_addr[13]), .B0(
        csr_add_x_421_n193), .SO(csr_n_T_250[14]) );
  AND4X1_LVT csr_add_x_421_U180 ( .A1(io_ptw_pmp_1_addr[11]), .A2(
        io_ptw_pmp_1_addr[12]), .A3(io_ptw_pmp_1_addr[13]), .A4(
        csr_add_x_421_n166), .Y(csr_add_x_421_n194) );
  HADDX1_LVT csr_add_x_421_U179 ( .A0(io_ptw_pmp_1_addr[14]), .B0(
        csr_add_x_421_n194), .SO(csr_n_T_250[15]) );
  NAND3X0_LVT csr_add_x_421_U178 ( .A1(io_ptw_pmp_1_addr[13]), .A2(
        io_ptw_pmp_1_addr[14]), .A3(csr_add_x_421_n193), .Y(csr_add_x_421_n192) );
  AO22X1_LVT csr_add_x_421_U177 ( .A1(io_ptw_pmp_1_addr[15]), .A2(
        csr_add_x_421_n192), .A3(csr_add_x_421_n163), .A4(csr_add_x_421_n164), 
        .Y(csr_n_T_250[16]) );
  AND2X1_LVT csr_add_x_421_U176 ( .A1(csr_add_x_421_n164), .A2(
        io_ptw_pmp_1_addr[15]), .Y(csr_add_x_421_n191) );
  HADDX1_LVT csr_add_x_421_U175 ( .A0(csr_add_x_421_n191), .B0(
        io_ptw_pmp_1_addr[16]), .SO(csr_n_T_250[17]) );
  AND3X1_LVT csr_add_x_421_U174 ( .A1(io_ptw_pmp_1_addr[15]), .A2(
        io_ptw_pmp_1_addr[16]), .A3(csr_add_x_421_n164), .Y(csr_add_x_421_n190) );
  HADDX1_LVT csr_add_x_421_U173 ( .A0(io_ptw_pmp_1_addr[17]), .B0(
        csr_add_x_421_n190), .SO(csr_n_T_250[18]) );
  AND4X1_LVT csr_add_x_421_U172 ( .A1(io_ptw_pmp_1_addr[15]), .A2(
        io_ptw_pmp_1_addr[16]), .A3(io_ptw_pmp_1_addr[17]), .A4(
        csr_add_x_421_n164), .Y(csr_add_x_421_n189) );
  HADDX1_LVT csr_add_x_421_U171 ( .A0(io_ptw_pmp_1_addr[18]), .B0(
        csr_add_x_421_n189), .SO(csr_n_T_250[19]) );
  AND4X1_LVT csr_add_x_421_U170 ( .A1(io_ptw_pmp_1_addr[15]), .A2(
        io_ptw_pmp_1_addr[16]), .A3(io_ptw_pmp_1_addr[18]), .A4(
        io_ptw_pmp_1_addr[17]), .Y(csr_add_x_421_n188) );
  NAND2X0_LVT csr_add_x_421_U169 ( .A1(csr_add_x_421_n188), .A2(
        csr_add_x_421_n164), .Y(csr_add_x_421_n187) );
  AO22X1_LVT csr_add_x_421_U168 ( .A1(io_ptw_pmp_1_addr[19]), .A2(
        csr_add_x_421_n187), .A3(csr_add_x_421_n161), .A4(csr_add_x_421_n162), 
        .Y(csr_n_T_250[20]) );
  AND2X1_LVT csr_add_x_421_U167 ( .A1(csr_add_x_421_n162), .A2(
        io_ptw_pmp_1_addr[19]), .Y(csr_add_x_421_n186) );
  HADDX1_LVT csr_add_x_421_U166 ( .A0(csr_add_x_421_n186), .B0(
        io_ptw_pmp_1_addr[20]), .SO(csr_n_T_250[21]) );
  AND3X1_LVT csr_add_x_421_U165 ( .A1(io_ptw_pmp_1_addr[19]), .A2(
        io_ptw_pmp_1_addr[20]), .A3(csr_add_x_421_n162), .Y(csr_add_x_421_n184) );
  HADDX1_LVT csr_add_x_421_U164 ( .A0(io_ptw_pmp_1_addr[21]), .B0(
        csr_add_x_421_n184), .SO(csr_n_T_250[22]) );
  AND2X1_LVT csr_add_x_421_U163 ( .A1(csr_add_x_421_n184), .A2(
        io_ptw_pmp_1_addr[21]), .Y(csr_add_x_421_n185) );
  HADDX1_LVT csr_add_x_421_U162 ( .A0(csr_add_x_421_n185), .B0(
        io_ptw_pmp_1_addr[22]), .SO(csr_n_T_250[23]) );
  NAND3X0_LVT csr_add_x_421_U161 ( .A1(io_ptw_pmp_1_addr[22]), .A2(
        io_ptw_pmp_1_addr[21]), .A3(csr_add_x_421_n184), .Y(csr_add_x_421_n183) );
  AO22X1_LVT csr_add_x_421_U160 ( .A1(io_ptw_pmp_1_addr[23]), .A2(
        csr_add_x_421_n183), .A3(csr_add_x_421_n159), .A4(csr_add_x_421_n160), 
        .Y(csr_n_T_250[24]) );
  AND2X1_LVT csr_add_x_421_U159 ( .A1(csr_add_x_421_n160), .A2(
        io_ptw_pmp_1_addr[23]), .Y(csr_add_x_421_n182) );
  HADDX1_LVT csr_add_x_421_U158 ( .A0(csr_add_x_421_n182), .B0(
        io_ptw_pmp_1_addr[24]), .SO(csr_n_T_250[25]) );
  AND3X1_LVT csr_add_x_421_U157 ( .A1(io_ptw_pmp_1_addr[23]), .A2(
        io_ptw_pmp_1_addr[24]), .A3(csr_add_x_421_n160), .Y(csr_add_x_421_n181) );
  HADDX1_LVT csr_add_x_421_U156 ( .A0(io_ptw_pmp_1_addr[25]), .B0(
        csr_add_x_421_n181), .SO(csr_n_T_250[26]) );
  AND2X1_LVT csr_add_x_421_U155 ( .A1(io_ptw_pmp_1_addr[25]), .A2(
        csr_add_x_421_n181), .Y(csr_add_x_421_n179) );
  HADDX1_LVT csr_add_x_421_U154 ( .A0(io_ptw_pmp_1_addr[26]), .B0(
        csr_add_x_421_n179), .SO(csr_n_T_250[27]) );
  AND2X1_LVT csr_add_x_421_U153 ( .A1(io_ptw_pmp_1_addr[26]), .A2(
        csr_add_x_421_n179), .Y(csr_add_x_421_n180) );
  HADDX1_LVT csr_add_x_421_U152 ( .A0(csr_add_x_421_n180), .B0(
        io_ptw_pmp_1_addr[27]), .SO(csr_n_T_250[28]) );
  AND3X1_LVT csr_add_x_421_U151 ( .A1(csr_add_x_421_n179), .A2(
        io_ptw_pmp_1_addr[26]), .A3(io_ptw_pmp_1_addr[27]), .Y(
        csr_add_x_421_n178) );
  HADDX1_LVT csr_add_x_421_U150 ( .A0(csr_add_x_421_n178), .B0(
        io_ptw_pmp_1_addr[28]), .SO(csr_n_T_250[29]) );
  HADDX1_LVT csr_add_x_421_U149 ( .A0(csr_add_x_421_n93), .B0(
        io_ptw_pmp_1_addr[1]), .SO(csr_n_T_250[2]) );
  AND2X1_LVT csr_add_x_421_U148 ( .A1(csr_add_x_421_n93), .A2(
        io_ptw_pmp_1_addr[1]), .Y(csr_add_x_421_n177) );
  HADDX1_LVT csr_add_x_421_U147 ( .A0(io_ptw_pmp_1_addr[2]), .B0(
        csr_add_x_421_n177), .SO(csr_n_T_250[3]) );
  AO22X1_LVT csr_add_x_421_U146 ( .A1(io_ptw_pmp_1_addr[3]), .A2(
        csr_add_x_421_n176), .A3(csr_add_x_421_n169), .A4(csr_add_x_421_n170), 
        .Y(csr_n_T_250[4]) );
  AND2X1_LVT csr_add_x_421_U145 ( .A1(csr_add_x_421_n170), .A2(
        io_ptw_pmp_1_addr[3]), .Y(csr_add_x_421_n175) );
  HADDX1_LVT csr_add_x_421_U144 ( .A0(csr_add_x_421_n175), .B0(
        io_ptw_pmp_1_addr[4]), .SO(csr_n_T_250[5]) );
  HADDX1_LVT csr_add_x_421_U143 ( .A0(io_ptw_pmp_1_addr[5]), .B0(
        csr_add_x_421_n174), .SO(csr_n_T_250[6]) );
  AND2X1_LVT csr_add_x_421_U142 ( .A1(io_ptw_pmp_1_addr[5]), .A2(
        csr_add_x_421_n174), .Y(csr_add_x_421_n173) );
  HADDX1_LVT csr_add_x_421_U141 ( .A0(io_ptw_pmp_1_addr[6]), .B0(
        csr_add_x_421_n173), .SO(csr_n_T_250[7]) );
  AO22X1_LVT csr_add_x_421_U140 ( .A1(csr_add_x_421_n168), .A2(
        csr_add_x_421_n167), .A3(csr_add_x_421_n172), .A4(io_ptw_pmp_1_addr[7]), .Y(csr_n_T_250[8]) );
  AND2X1_LVT csr_add_x_421_U139 ( .A1(io_ptw_pmp_1_addr[7]), .A2(
        csr_add_x_421_n168), .Y(csr_add_x_421_n171) );
  HADDX1_LVT csr_add_x_421_U138 ( .A0(csr_add_x_421_n171), .B0(
        io_ptw_pmp_1_addr[8]), .SO(csr_n_T_250[9]) );
  INVX1_LVT csr_add_x_421_U137 ( .A(csr_add_x_421_n176), .Y(csr_add_x_421_n170) );
  INVX1_LVT csr_add_x_421_U136 ( .A(io_ptw_pmp_1_addr[3]), .Y(
        csr_add_x_421_n169) );
  INVX1_LVT csr_add_x_421_U135 ( .A(csr_add_x_421_n172), .Y(csr_add_x_421_n168) );
  INVX1_LVT csr_add_x_421_U134 ( .A(io_ptw_pmp_1_addr[7]), .Y(
        csr_add_x_421_n167) );
  INVX1_LVT csr_add_x_421_U133 ( .A(csr_add_x_421_n196), .Y(csr_add_x_421_n166) );
  INVX1_LVT csr_add_x_421_U132 ( .A(io_ptw_pmp_1_addr[11]), .Y(
        csr_add_x_421_n165) );
  INVX1_LVT csr_add_x_421_U131 ( .A(csr_add_x_421_n192), .Y(csr_add_x_421_n164) );
  INVX1_LVT csr_add_x_421_U130 ( .A(io_ptw_pmp_1_addr[15]), .Y(
        csr_add_x_421_n163) );
  INVX1_LVT csr_add_x_421_U129 ( .A(csr_add_x_421_n187), .Y(csr_add_x_421_n162) );
  INVX1_LVT csr_add_x_421_U128 ( .A(io_ptw_pmp_1_addr[19]), .Y(
        csr_add_x_421_n161) );
  INVX1_LVT csr_add_x_421_U127 ( .A(csr_add_x_421_n183), .Y(csr_add_x_421_n160) );
  INVX1_LVT csr_add_x_421_U126 ( .A(io_ptw_pmp_1_addr[23]), .Y(
        csr_add_x_421_n159) );
  HADDX1_LVT csr_add_x_421_U121 ( .A0(io_ptw_pmp_1_addr[0]), .B0(
        io_ptw_pmp_1_cfg_a[0]), .C1(csr_add_x_421_n93), .SO(csr_n_T_250[1]) );
  NAND3X0_LVT csr_add_x_420_U194 ( .A1(csr_add_x_420_n93), .A2(
        io_ptw_pmp_0_addr[1]), .A3(io_ptw_pmp_0_addr[2]), .Y(
        csr_add_x_420_n176) );
  AND3X1_LVT csr_add_x_420_U193 ( .A1(io_ptw_pmp_0_addr[3]), .A2(
        io_ptw_pmp_0_addr[4]), .A3(csr_add_x_420_n164), .Y(csr_add_x_420_n174)
         );
  NAND3X0_LVT csr_add_x_420_U192 ( .A1(io_ptw_pmp_0_addr[5]), .A2(
        io_ptw_pmp_0_addr[6]), .A3(csr_add_x_420_n174), .Y(csr_add_x_420_n172)
         );
  AND3X1_LVT csr_add_x_420_U191 ( .A1(csr_add_x_420_n163), .A2(
        io_ptw_pmp_0_addr[8]), .A3(io_ptw_pmp_0_addr[7]), .Y(
        csr_add_x_420_n199) );
  HADDX1_LVT csr_add_x_420_U190 ( .A0(io_ptw_pmp_0_addr[9]), .B0(
        csr_add_x_420_n199), .SO(csr_n_T_241[10]) );
  AND4X1_LVT csr_add_x_420_U189 ( .A1(csr_add_x_420_n163), .A2(
        io_ptw_pmp_0_addr[8]), .A3(io_ptw_pmp_0_addr[7]), .A4(
        io_ptw_pmp_0_addr[9]), .Y(csr_add_x_420_n198) );
  HADDX1_LVT csr_add_x_420_U188 ( .A0(io_ptw_pmp_0_addr[10]), .B0(
        csr_add_x_420_n198), .SO(csr_n_T_241[11]) );
  AND4X1_LVT csr_add_x_420_U187 ( .A1(io_ptw_pmp_0_addr[8]), .A2(
        io_ptw_pmp_0_addr[7]), .A3(io_ptw_pmp_0_addr[10]), .A4(
        io_ptw_pmp_0_addr[9]), .Y(csr_add_x_420_n197) );
  NAND2X0_LVT csr_add_x_420_U186 ( .A1(csr_add_x_420_n163), .A2(
        csr_add_x_420_n197), .Y(csr_add_x_420_n196) );
  AO22X1_LVT csr_add_x_420_U185 ( .A1(io_ptw_pmp_0_addr[11]), .A2(
        csr_add_x_420_n196), .A3(csr_add_x_420_n168), .A4(csr_add_x_420_n162), 
        .Y(csr_n_T_241[12]) );
  AND2X1_LVT csr_add_x_420_U184 ( .A1(csr_add_x_420_n162), .A2(
        io_ptw_pmp_0_addr[11]), .Y(csr_add_x_420_n195) );
  HADDX1_LVT csr_add_x_420_U183 ( .A0(csr_add_x_420_n195), .B0(
        io_ptw_pmp_0_addr[12]), .SO(csr_n_T_241[13]) );
  AND3X1_LVT csr_add_x_420_U182 ( .A1(io_ptw_pmp_0_addr[11]), .A2(
        io_ptw_pmp_0_addr[12]), .A3(csr_add_x_420_n162), .Y(csr_add_x_420_n193) );
  HADDX1_LVT csr_add_x_420_U181 ( .A0(io_ptw_pmp_0_addr[13]), .B0(
        csr_add_x_420_n193), .SO(csr_n_T_241[14]) );
  AND4X1_LVT csr_add_x_420_U180 ( .A1(io_ptw_pmp_0_addr[11]), .A2(
        io_ptw_pmp_0_addr[12]), .A3(io_ptw_pmp_0_addr[13]), .A4(
        csr_add_x_420_n162), .Y(csr_add_x_420_n194) );
  HADDX1_LVT csr_add_x_420_U179 ( .A0(io_ptw_pmp_0_addr[14]), .B0(
        csr_add_x_420_n194), .SO(csr_n_T_241[15]) );
  NAND3X0_LVT csr_add_x_420_U178 ( .A1(io_ptw_pmp_0_addr[13]), .A2(
        io_ptw_pmp_0_addr[14]), .A3(csr_add_x_420_n193), .Y(csr_add_x_420_n192) );
  AO22X1_LVT csr_add_x_420_U177 ( .A1(io_ptw_pmp_0_addr[15]), .A2(
        csr_add_x_420_n192), .A3(csr_add_x_420_n167), .A4(csr_add_x_420_n161), 
        .Y(csr_n_T_241[16]) );
  AND2X1_LVT csr_add_x_420_U176 ( .A1(csr_add_x_420_n161), .A2(
        io_ptw_pmp_0_addr[15]), .Y(csr_add_x_420_n191) );
  HADDX1_LVT csr_add_x_420_U175 ( .A0(csr_add_x_420_n191), .B0(
        io_ptw_pmp_0_addr[16]), .SO(csr_n_T_241[17]) );
  AND3X1_LVT csr_add_x_420_U174 ( .A1(io_ptw_pmp_0_addr[15]), .A2(
        io_ptw_pmp_0_addr[16]), .A3(csr_add_x_420_n161), .Y(csr_add_x_420_n190) );
  HADDX1_LVT csr_add_x_420_U173 ( .A0(io_ptw_pmp_0_addr[17]), .B0(
        csr_add_x_420_n190), .SO(csr_n_T_241[18]) );
  AND4X1_LVT csr_add_x_420_U172 ( .A1(io_ptw_pmp_0_addr[15]), .A2(
        io_ptw_pmp_0_addr[16]), .A3(io_ptw_pmp_0_addr[17]), .A4(
        csr_add_x_420_n161), .Y(csr_add_x_420_n189) );
  HADDX1_LVT csr_add_x_420_U171 ( .A0(io_ptw_pmp_0_addr[18]), .B0(
        csr_add_x_420_n189), .SO(csr_n_T_241[19]) );
  AND4X1_LVT csr_add_x_420_U170 ( .A1(io_ptw_pmp_0_addr[15]), .A2(
        io_ptw_pmp_0_addr[16]), .A3(io_ptw_pmp_0_addr[18]), .A4(
        io_ptw_pmp_0_addr[17]), .Y(csr_add_x_420_n188) );
  NAND2X0_LVT csr_add_x_420_U169 ( .A1(csr_add_x_420_n188), .A2(
        csr_add_x_420_n161), .Y(csr_add_x_420_n187) );
  AO22X1_LVT csr_add_x_420_U168 ( .A1(io_ptw_pmp_0_addr[19]), .A2(
        csr_add_x_420_n187), .A3(csr_add_x_420_n166), .A4(csr_add_x_420_n160), 
        .Y(csr_n_T_241[20]) );
  AND2X1_LVT csr_add_x_420_U167 ( .A1(csr_add_x_420_n160), .A2(
        io_ptw_pmp_0_addr[19]), .Y(csr_add_x_420_n186) );
  HADDX1_LVT csr_add_x_420_U166 ( .A0(csr_add_x_420_n186), .B0(
        io_ptw_pmp_0_addr[20]), .SO(csr_n_T_241[21]) );
  AND3X1_LVT csr_add_x_420_U165 ( .A1(io_ptw_pmp_0_addr[19]), .A2(
        io_ptw_pmp_0_addr[20]), .A3(csr_add_x_420_n160), .Y(csr_add_x_420_n184) );
  HADDX1_LVT csr_add_x_420_U164 ( .A0(io_ptw_pmp_0_addr[21]), .B0(
        csr_add_x_420_n184), .SO(csr_n_T_241[22]) );
  AND2X1_LVT csr_add_x_420_U163 ( .A1(csr_add_x_420_n184), .A2(
        io_ptw_pmp_0_addr[21]), .Y(csr_add_x_420_n185) );
  HADDX1_LVT csr_add_x_420_U162 ( .A0(csr_add_x_420_n185), .B0(
        io_ptw_pmp_0_addr[22]), .SO(csr_n_T_241[23]) );
  NAND3X0_LVT csr_add_x_420_U161 ( .A1(io_ptw_pmp_0_addr[22]), .A2(
        io_ptw_pmp_0_addr[21]), .A3(csr_add_x_420_n184), .Y(csr_add_x_420_n183) );
  AO22X1_LVT csr_add_x_420_U160 ( .A1(io_ptw_pmp_0_addr[23]), .A2(
        csr_add_x_420_n183), .A3(csr_add_x_420_n165), .A4(csr_add_x_420_n159), 
        .Y(csr_n_T_241[24]) );
  AND2X1_LVT csr_add_x_420_U159 ( .A1(csr_add_x_420_n159), .A2(
        io_ptw_pmp_0_addr[23]), .Y(csr_add_x_420_n182) );
  HADDX1_LVT csr_add_x_420_U158 ( .A0(csr_add_x_420_n182), .B0(
        io_ptw_pmp_0_addr[24]), .SO(csr_n_T_241[25]) );
  AND3X1_LVT csr_add_x_420_U157 ( .A1(io_ptw_pmp_0_addr[23]), .A2(
        io_ptw_pmp_0_addr[24]), .A3(csr_add_x_420_n159), .Y(csr_add_x_420_n181) );
  HADDX1_LVT csr_add_x_420_U156 ( .A0(io_ptw_pmp_0_addr[25]), .B0(
        csr_add_x_420_n181), .SO(csr_n_T_241[26]) );
  AND2X1_LVT csr_add_x_420_U155 ( .A1(io_ptw_pmp_0_addr[25]), .A2(
        csr_add_x_420_n181), .Y(csr_add_x_420_n179) );
  HADDX1_LVT csr_add_x_420_U154 ( .A0(io_ptw_pmp_0_addr[26]), .B0(
        csr_add_x_420_n179), .SO(csr_n_T_241[27]) );
  AND2X1_LVT csr_add_x_420_U153 ( .A1(io_ptw_pmp_0_addr[26]), .A2(
        csr_add_x_420_n179), .Y(csr_add_x_420_n180) );
  HADDX1_LVT csr_add_x_420_U152 ( .A0(csr_add_x_420_n180), .B0(
        io_ptw_pmp_0_addr[27]), .SO(csr_n_T_241[28]) );
  AND3X1_LVT csr_add_x_420_U151 ( .A1(csr_add_x_420_n179), .A2(
        io_ptw_pmp_0_addr[26]), .A3(io_ptw_pmp_0_addr[27]), .Y(
        csr_add_x_420_n178) );
  HADDX1_LVT csr_add_x_420_U150 ( .A0(csr_add_x_420_n178), .B0(
        io_ptw_pmp_0_addr[28]), .SO(csr_n_T_241[29]) );
  HADDX1_LVT csr_add_x_420_U149 ( .A0(csr_add_x_420_n93), .B0(
        io_ptw_pmp_0_addr[1]), .SO(csr_n_T_241[2]) );
  AND2X1_LVT csr_add_x_420_U148 ( .A1(csr_add_x_420_n93), .A2(
        io_ptw_pmp_0_addr[1]), .Y(csr_add_x_420_n177) );
  HADDX1_LVT csr_add_x_420_U147 ( .A0(io_ptw_pmp_0_addr[2]), .B0(
        csr_add_x_420_n177), .SO(csr_n_T_241[3]) );
  AO22X1_LVT csr_add_x_420_U146 ( .A1(io_ptw_pmp_0_addr[3]), .A2(
        csr_add_x_420_n176), .A3(csr_add_x_420_n170), .A4(csr_add_x_420_n164), 
        .Y(csr_n_T_241[4]) );
  AND2X1_LVT csr_add_x_420_U145 ( .A1(csr_add_x_420_n164), .A2(
        io_ptw_pmp_0_addr[3]), .Y(csr_add_x_420_n175) );
  HADDX1_LVT csr_add_x_420_U144 ( .A0(csr_add_x_420_n175), .B0(
        io_ptw_pmp_0_addr[4]), .SO(csr_n_T_241[5]) );
  HADDX1_LVT csr_add_x_420_U143 ( .A0(io_ptw_pmp_0_addr[5]), .B0(
        csr_add_x_420_n174), .SO(csr_n_T_241[6]) );
  AND2X1_LVT csr_add_x_420_U142 ( .A1(io_ptw_pmp_0_addr[5]), .A2(
        csr_add_x_420_n174), .Y(csr_add_x_420_n173) );
  HADDX1_LVT csr_add_x_420_U141 ( .A0(io_ptw_pmp_0_addr[6]), .B0(
        csr_add_x_420_n173), .SO(csr_n_T_241[7]) );
  AO22X1_LVT csr_add_x_420_U140 ( .A1(csr_add_x_420_n163), .A2(
        csr_add_x_420_n169), .A3(csr_add_x_420_n172), .A4(io_ptw_pmp_0_addr[7]), .Y(csr_n_T_241[8]) );
  AND2X1_LVT csr_add_x_420_U139 ( .A1(io_ptw_pmp_0_addr[7]), .A2(
        csr_add_x_420_n163), .Y(csr_add_x_420_n171) );
  HADDX1_LVT csr_add_x_420_U138 ( .A0(csr_add_x_420_n171), .B0(
        io_ptw_pmp_0_addr[8]), .SO(csr_n_T_241[9]) );
  INVX1_LVT csr_add_x_420_U137 ( .A(io_ptw_pmp_0_addr[3]), .Y(
        csr_add_x_420_n170) );
  INVX1_LVT csr_add_x_420_U136 ( .A(io_ptw_pmp_0_addr[7]), .Y(
        csr_add_x_420_n169) );
  INVX1_LVT csr_add_x_420_U135 ( .A(io_ptw_pmp_0_addr[11]), .Y(
        csr_add_x_420_n168) );
  INVX1_LVT csr_add_x_420_U134 ( .A(io_ptw_pmp_0_addr[15]), .Y(
        csr_add_x_420_n167) );
  INVX1_LVT csr_add_x_420_U133 ( .A(io_ptw_pmp_0_addr[19]), .Y(
        csr_add_x_420_n166) );
  INVX1_LVT csr_add_x_420_U132 ( .A(io_ptw_pmp_0_addr[23]), .Y(
        csr_add_x_420_n165) );
  INVX1_LVT csr_add_x_420_U131 ( .A(csr_add_x_420_n176), .Y(csr_add_x_420_n164) );
  INVX1_LVT csr_add_x_420_U130 ( .A(csr_add_x_420_n172), .Y(csr_add_x_420_n163) );
  INVX1_LVT csr_add_x_420_U129 ( .A(csr_add_x_420_n196), .Y(csr_add_x_420_n162) );
  INVX1_LVT csr_add_x_420_U128 ( .A(csr_add_x_420_n192), .Y(csr_add_x_420_n161) );
  INVX1_LVT csr_add_x_420_U127 ( .A(csr_add_x_420_n187), .Y(csr_add_x_420_n160) );
  INVX1_LVT csr_add_x_420_U126 ( .A(csr_add_x_420_n183), .Y(csr_add_x_420_n159) );
  HADDX1_LVT csr_add_x_420_U121 ( .A0(io_ptw_pmp_0_addr[0]), .B0(
        io_ptw_pmp_0_cfg_a[0]), .C1(csr_add_x_420_n93), .SO(csr_n_T_241[1]) );
  NAND3X0_LVT csr_add_x_381_U406 ( .A1(csr_add_x_381_n203), .A2(csr_io_time[8]), .A3(csr_io_time[9]), .Y(csr_add_x_381_n359) );
  AND3X1_LVT csr_add_x_381_U405 ( .A1(csr_io_time[10]), .A2(csr_io_time[11]), 
        .A3(csr_add_x_381_n344), .Y(csr_add_x_381_n348) );
  NAND3X0_LVT csr_add_x_381_U404 ( .A1(csr_io_time[12]), .A2(csr_io_time[13]), 
        .A3(csr_add_x_381_n348), .Y(csr_add_x_381_n346) );
  AND3X1_LVT csr_add_x_381_U403 ( .A1(csr_add_x_381_n342), .A2(csr_io_time[15]), .A3(csr_io_time[14]), .Y(csr_add_x_381_n411) );
  HADDX1_LVT csr_add_x_381_U402 ( .A0(csr_io_time[16]), .B0(csr_add_x_381_n411), .SO(csr_n_T_52[10]) );
  AND4X1_LVT csr_add_x_381_U401 ( .A1(csr_add_x_381_n342), .A2(csr_io_time[15]), .A3(csr_io_time[14]), .A4(csr_io_time[16]), .Y(csr_add_x_381_n410) );
  HADDX1_LVT csr_add_x_381_U400 ( .A0(csr_io_time[17]), .B0(csr_add_x_381_n410), .SO(csr_n_T_52[11]) );
  AND4X1_LVT csr_add_x_381_U399 ( .A1(csr_io_time[15]), .A2(csr_io_time[14]), 
        .A3(csr_io_time[17]), .A4(csr_io_time[16]), .Y(csr_add_x_381_n409) );
  NAND2X0_LVT csr_add_x_381_U398 ( .A1(csr_add_x_381_n342), .A2(
        csr_add_x_381_n409), .Y(csr_add_x_381_n408) );
  AO22X1_LVT csr_add_x_381_U397 ( .A1(csr_io_time[18]), .A2(csr_add_x_381_n408), .A3(csr_add_x_381_n339), .A4(csr_add_x_381_n340), .Y(csr_n_T_52[12]) );
  AND2X1_LVT csr_add_x_381_U396 ( .A1(csr_add_x_381_n340), .A2(csr_io_time[18]), .Y(csr_add_x_381_n407) );
  HADDX1_LVT csr_add_x_381_U395 ( .A0(csr_add_x_381_n407), .B0(csr_io_time[19]), .SO(csr_n_T_52[13]) );
  AND3X1_LVT csr_add_x_381_U394 ( .A1(csr_io_time[18]), .A2(csr_io_time[19]), 
        .A3(csr_add_x_381_n340), .Y(csr_add_x_381_n405) );
  HADDX1_LVT csr_add_x_381_U393 ( .A0(csr_io_time[20]), .B0(csr_add_x_381_n405), .SO(csr_n_T_52[14]) );
  AND4X1_LVT csr_add_x_381_U392 ( .A1(csr_io_time[18]), .A2(csr_io_time[19]), 
        .A3(csr_io_time[20]), .A4(csr_add_x_381_n340), .Y(csr_add_x_381_n406)
         );
  HADDX1_LVT csr_add_x_381_U391 ( .A0(csr_io_time[21]), .B0(csr_add_x_381_n406), .SO(csr_n_T_52[15]) );
  NAND3X0_LVT csr_add_x_381_U390 ( .A1(csr_io_time[20]), .A2(csr_io_time[21]), 
        .A3(csr_add_x_381_n405), .Y(csr_add_x_381_n404) );
  AO22X1_LVT csr_add_x_381_U389 ( .A1(csr_io_time[22]), .A2(csr_add_x_381_n404), .A3(csr_add_x_381_n337), .A4(csr_add_x_381_n338), .Y(csr_n_T_52[16]) );
  AND2X1_LVT csr_add_x_381_U388 ( .A1(csr_add_x_381_n338), .A2(csr_io_time[22]), .Y(csr_add_x_381_n403) );
  HADDX1_LVT csr_add_x_381_U387 ( .A0(csr_add_x_381_n403), .B0(csr_io_time[23]), .SO(csr_n_T_52[17]) );
  AND3X1_LVT csr_add_x_381_U386 ( .A1(csr_io_time[22]), .A2(csr_io_time[23]), 
        .A3(csr_add_x_381_n338), .Y(csr_add_x_381_n402) );
  HADDX1_LVT csr_add_x_381_U385 ( .A0(csr_io_time[24]), .B0(csr_add_x_381_n402), .SO(csr_n_T_52[18]) );
  AND4X1_LVT csr_add_x_381_U384 ( .A1(csr_io_time[22]), .A2(csr_io_time[23]), 
        .A3(csr_io_time[24]), .A4(csr_add_x_381_n338), .Y(csr_add_x_381_n401)
         );
  HADDX1_LVT csr_add_x_381_U383 ( .A0(csr_io_time[25]), .B0(csr_add_x_381_n401), .SO(csr_n_T_52[19]) );
  AND4X1_LVT csr_add_x_381_U382 ( .A1(csr_io_time[22]), .A2(csr_io_time[23]), 
        .A3(csr_io_time[25]), .A4(csr_io_time[24]), .Y(csr_add_x_381_n396) );
  AND2X1_LVT csr_add_x_381_U381 ( .A1(csr_add_x_381_n396), .A2(
        csr_add_x_381_n338), .Y(csr_add_x_381_n400) );
  HADDX1_LVT csr_add_x_381_U380 ( .A0(csr_io_time[26]), .B0(csr_add_x_381_n400), .SO(csr_n_T_52[20]) );
  AND3X1_LVT csr_add_x_381_U379 ( .A1(csr_add_x_381_n396), .A2(csr_io_time[26]), .A3(csr_add_x_381_n338), .Y(csr_add_x_381_n399) );
  HADDX1_LVT csr_add_x_381_U378 ( .A0(csr_add_x_381_n399), .B0(csr_io_time[27]), .SO(csr_n_T_52[21]) );
  AND2X1_LVT csr_add_x_381_U377 ( .A1(csr_io_time[26]), .A2(csr_io_time[27]), 
        .Y(csr_add_x_381_n395) );
  AND3X1_LVT csr_add_x_381_U376 ( .A1(csr_add_x_381_n395), .A2(
        csr_add_x_381_n396), .A3(csr_add_x_381_n338), .Y(csr_add_x_381_n398)
         );
  HADDX1_LVT csr_add_x_381_U375 ( .A0(csr_io_time[28]), .B0(csr_add_x_381_n398), .SO(csr_n_T_52[22]) );
  AND4X1_LVT csr_add_x_381_U374 ( .A1(csr_io_time[28]), .A2(csr_add_x_381_n395), .A3(csr_add_x_381_n396), .A4(csr_add_x_381_n338), .Y(csr_add_x_381_n397) );
  HADDX1_LVT csr_add_x_381_U373 ( .A0(csr_io_time[29]), .B0(csr_add_x_381_n397), .SO(csr_n_T_52[23]) );
  AND4X1_LVT csr_add_x_381_U372 ( .A1(csr_io_time[28]), .A2(csr_io_time[29]), 
        .A3(csr_add_x_381_n395), .A4(csr_add_x_381_n396), .Y(
        csr_add_x_381_n394) );
  NAND2X0_LVT csr_add_x_381_U371 ( .A1(csr_add_x_381_n394), .A2(
        csr_add_x_381_n338), .Y(csr_add_x_381_n393) );
  AO22X1_LVT csr_add_x_381_U370 ( .A1(csr_io_time[30]), .A2(csr_add_x_381_n393), .A3(csr_add_x_381_n335), .A4(csr_add_x_381_n336), .Y(csr_n_T_52[24]) );
  AND2X1_LVT csr_add_x_381_U369 ( .A1(csr_add_x_381_n336), .A2(csr_io_time[30]), .Y(csr_add_x_381_n392) );
  HADDX1_LVT csr_add_x_381_U368 ( .A0(csr_add_x_381_n392), .B0(csr_io_time[31]), .SO(csr_n_T_52[25]) );
  AND3X1_LVT csr_add_x_381_U367 ( .A1(csr_io_time[30]), .A2(csr_io_time[31]), 
        .A3(csr_add_x_381_n336), .Y(csr_add_x_381_n391) );
  HADDX1_LVT csr_add_x_381_U366 ( .A0(csr_n1967), .B0(csr_add_x_381_n391), 
        .SO(csr_n_T_52[26]) );
  AND4X1_LVT csr_add_x_381_U365 ( .A1(csr_io_time[30]), .A2(csr_io_time[31]), 
        .A3(csr_n1967), .A4(csr_add_x_381_n336), .Y(csr_add_x_381_n390) );
  HADDX1_LVT csr_add_x_381_U364 ( .A0(csr_n1966), .B0(csr_add_x_381_n390), 
        .SO(csr_n_T_52[27]) );
  AND4X1_LVT csr_add_x_381_U363 ( .A1(csr_io_time[30]), .A2(csr_io_time[31]), 
        .A3(csr_n1966), .A4(csr_n1967), .Y(csr_add_x_381_n387) );
  AND2X1_LVT csr_add_x_381_U362 ( .A1(csr_add_x_381_n387), .A2(
        csr_add_x_381_n336), .Y(csr_add_x_381_n385) );
  HADDX1_LVT csr_add_x_381_U361 ( .A0(csr_n1965), .B0(csr_add_x_381_n385), 
        .SO(csr_n_T_52[28]) );
  AND3X1_LVT csr_add_x_381_U360 ( .A1(csr_n1965), .A2(csr_add_x_381_n387), 
        .A3(csr_add_x_381_n336), .Y(csr_add_x_381_n389) );
  HADDX1_LVT csr_add_x_381_U359 ( .A0(csr_add_x_381_n389), .B0(csr_n1964), 
        .SO(csr_n_T_52[29]) );
  HADDX1_LVT csr_add_x_381_U358 ( .A0(csr_add_x_381_n203), .B0(csr_io_time[8]), 
        .SO(csr_n_T_52[2]) );
  AND2X1_LVT csr_add_x_381_U357 ( .A1(csr_n1965), .A2(csr_n1964), .Y(
        csr_add_x_381_n384) );
  AND3X1_LVT csr_add_x_381_U356 ( .A1(csr_add_x_381_n387), .A2(
        csr_add_x_381_n384), .A3(csr_add_x_381_n336), .Y(csr_add_x_381_n388)
         );
  HADDX1_LVT csr_add_x_381_U355 ( .A0(csr_n1963), .B0(csr_add_x_381_n388), 
        .SO(csr_n_T_52[30]) );
  AND4X1_LVT csr_add_x_381_U354 ( .A1(csr_add_x_381_n387), .A2(csr_n1963), 
        .A3(csr_add_x_381_n384), .A4(csr_add_x_381_n336), .Y(
        csr_add_x_381_n386) );
  HADDX1_LVT csr_add_x_381_U353 ( .A0(csr_n1962), .B0(csr_add_x_381_n386), 
        .SO(csr_n_T_52[31]) );
  NAND4X0_LVT csr_add_x_381_U352 ( .A1(csr_n1962), .A2(csr_n1963), .A3(
        csr_add_x_381_n384), .A4(csr_add_x_381_n385), .Y(csr_add_x_381_n383)
         );
  AND2X1_LVT csr_add_x_381_U351 ( .A1(csr_n1961), .A2(csr_add_x_381_n334), .Y(
        csr_add_x_381_n382) );
  HADDX1_LVT csr_add_x_381_U350 ( .A0(csr_add_x_381_n382), .B0(csr_n1960), 
        .SO(csr_n_T_52[33]) );
  AND3X1_LVT csr_add_x_381_U349 ( .A1(csr_add_x_381_n334), .A2(csr_n1961), 
        .A3(csr_n1960), .Y(csr_add_x_381_n381) );
  HADDX1_LVT csr_add_x_381_U348 ( .A0(csr_n1959), .B0(csr_add_x_381_n381), 
        .SO(csr_n_T_52[34]) );
  AND4X1_LVT csr_add_x_381_U347 ( .A1(csr_add_x_381_n334), .A2(csr_n1961), 
        .A3(csr_n1960), .A4(csr_n1959), .Y(csr_add_x_381_n380) );
  HADDX1_LVT csr_add_x_381_U346 ( .A0(csr_n1958), .B0(csr_add_x_381_n380), 
        .SO(csr_n_T_52[35]) );
  AND4X1_LVT csr_add_x_381_U345 ( .A1(csr_n1961), .A2(csr_n1960), .A3(
        csr_n1958), .A4(csr_n1959), .Y(csr_add_x_381_n374) );
  AND2X1_LVT csr_add_x_381_U344 ( .A1(csr_add_x_381_n334), .A2(
        csr_add_x_381_n374), .Y(csr_add_x_381_n379) );
  HADDX1_LVT csr_add_x_381_U343 ( .A0(csr_n1957), .B0(csr_add_x_381_n379), 
        .SO(csr_n_T_52[36]) );
  AND3X1_LVT csr_add_x_381_U342 ( .A1(csr_n1957), .A2(csr_add_x_381_n334), 
        .A3(csr_add_x_381_n374), .Y(csr_add_x_381_n378) );
  HADDX1_LVT csr_add_x_381_U341 ( .A0(csr_add_x_381_n378), .B0(csr_n1956), 
        .SO(csr_n_T_52[37]) );
  AND2X1_LVT csr_add_x_381_U340 ( .A1(csr_n1957), .A2(csr_n1956), .Y(
        csr_add_x_381_n373) );
  AND3X1_LVT csr_add_x_381_U339 ( .A1(csr_add_x_381_n334), .A2(
        csr_add_x_381_n373), .A3(csr_add_x_381_n374), .Y(csr_add_x_381_n377)
         );
  HADDX1_LVT csr_add_x_381_U338 ( .A0(csr_n1955), .B0(csr_add_x_381_n377), 
        .SO(csr_n_T_52[38]) );
  AND4X1_LVT csr_add_x_381_U337 ( .A1(csr_add_x_381_n334), .A2(csr_n1955), 
        .A3(csr_add_x_381_n373), .A4(csr_add_x_381_n374), .Y(
        csr_add_x_381_n376) );
  HADDX1_LVT csr_add_x_381_U336 ( .A0(csr_n1954), .B0(csr_add_x_381_n376), 
        .SO(csr_n_T_52[39]) );
  AND2X1_LVT csr_add_x_381_U335 ( .A1(csr_add_x_381_n203), .A2(csr_io_time[8]), 
        .Y(csr_add_x_381_n375) );
  HADDX1_LVT csr_add_x_381_U334 ( .A0(csr_io_time[9]), .B0(csr_add_x_381_n375), 
        .SO(csr_n_T_52[3]) );
  AND4X1_LVT csr_add_x_381_U333 ( .A1(csr_n1955), .A2(csr_n1954), .A3(
        csr_add_x_381_n373), .A4(csr_add_x_381_n374), .Y(csr_add_x_381_n372)
         );
  NAND2X0_LVT csr_add_x_381_U332 ( .A1(csr_add_x_381_n334), .A2(
        csr_add_x_381_n372), .Y(csr_add_x_381_n371) );
  AO22X1_LVT csr_add_x_381_U331 ( .A1(csr_n1953), .A2(csr_add_x_381_n371), 
        .A3(csr_add_x_381_n332), .A4(csr_add_x_381_n333), .Y(csr_n_T_52[40])
         );
  AND2X1_LVT csr_add_x_381_U330 ( .A1(csr_add_x_381_n333), .A2(csr_n1953), .Y(
        csr_add_x_381_n370) );
  HADDX1_LVT csr_add_x_381_U329 ( .A0(csr_add_x_381_n370), .B0(csr_n1952), 
        .SO(csr_n_T_52[41]) );
  AND3X1_LVT csr_add_x_381_U328 ( .A1(csr_n1953), .A2(csr_n1952), .A3(
        csr_add_x_381_n333), .Y(csr_add_x_381_n369) );
  HADDX1_LVT csr_add_x_381_U327 ( .A0(csr_n1951), .B0(csr_add_x_381_n369), 
        .SO(csr_n_T_52[42]) );
  AND4X1_LVT csr_add_x_381_U326 ( .A1(csr_n1953), .A2(csr_n1952), .A3(
        csr_n1951), .A4(csr_add_x_381_n333), .Y(csr_add_x_381_n368) );
  HADDX1_LVT csr_add_x_381_U325 ( .A0(csr_n1950), .B0(csr_add_x_381_n368), 
        .SO(csr_n_T_52[43]) );
  AND4X1_LVT csr_add_x_381_U324 ( .A1(csr_n1953), .A2(csr_n1952), .A3(
        csr_n1950), .A4(csr_n1951), .Y(csr_add_x_381_n363) );
  NAND2X0_LVT csr_add_x_381_U323 ( .A1(csr_add_x_381_n363), .A2(
        csr_add_x_381_n333), .Y(csr_add_x_381_n367) );
  AND2X1_LVT csr_add_x_381_U322 ( .A1(csr_add_x_381_n331), .A2(csr_n1949), .Y(
        csr_add_x_381_n366) );
  HADDX1_LVT csr_add_x_381_U321 ( .A0(csr_add_x_381_n366), .B0(csr_n1948), 
        .SO(csr_n_T_52[45]) );
  AND3X1_LVT csr_add_x_381_U320 ( .A1(csr_n1949), .A2(csr_n1948), .A3(
        csr_add_x_381_n331), .Y(csr_add_x_381_n365) );
  HADDX1_LVT csr_add_x_381_U319 ( .A0(csr_n1947), .B0(csr_add_x_381_n365), 
        .SO(csr_n_T_52[46]) );
  AND4X1_LVT csr_add_x_381_U318 ( .A1(csr_n1947), .A2(csr_n1949), .A3(
        csr_n1948), .A4(csr_add_x_381_n331), .Y(csr_add_x_381_n364) );
  HADDX1_LVT csr_add_x_381_U317 ( .A0(csr_n1946), .B0(csr_add_x_381_n364), 
        .SO(csr_n_T_52[47]) );
  AND4X1_LVT csr_add_x_381_U316 ( .A1(csr_n1949), .A2(csr_n1948), .A3(
        csr_add_x_381_n363), .A4(csr_add_x_381_n333), .Y(csr_add_x_381_n362)
         );
  NAND3X0_LVT csr_add_x_381_U315 ( .A1(csr_n1946), .A2(csr_n1947), .A3(
        csr_add_x_381_n362), .Y(csr_add_x_381_n361) );
  AND2X1_LVT csr_add_x_381_U314 ( .A1(csr_add_x_381_n330), .A2(csr_n1945), .Y(
        csr_add_x_381_n360) );
  HADDX1_LVT csr_add_x_381_U313 ( .A0(csr_add_x_381_n360), .B0(csr_n1944), 
        .SO(csr_n_T_52[49]) );
  AO22X1_LVT csr_add_x_381_U312 ( .A1(csr_io_time[10]), .A2(csr_add_x_381_n359), .A3(csr_add_x_381_n343), .A4(csr_add_x_381_n344), .Y(csr_n_T_52[4]) );
  AND3X1_LVT csr_add_x_381_U311 ( .A1(csr_n1945), .A2(csr_n1944), .A3(
        csr_add_x_381_n330), .Y(csr_add_x_381_n358) );
  HADDX1_LVT csr_add_x_381_U310 ( .A0(csr_n1943), .B0(csr_add_x_381_n358), 
        .SO(csr_n_T_52[50]) );
  AND4X1_LVT csr_add_x_381_U309 ( .A1(csr_n1945), .A2(csr_n1944), .A3(
        csr_n1943), .A4(csr_add_x_381_n330), .Y(csr_add_x_381_n357) );
  HADDX1_LVT csr_add_x_381_U308 ( .A0(csr_n1942), .B0(csr_add_x_381_n357), 
        .SO(csr_n_T_52[51]) );
  AND4X1_LVT csr_add_x_381_U307 ( .A1(csr_n1945), .A2(csr_n1944), .A3(
        csr_n1942), .A4(csr_n1943), .Y(csr_add_x_381_n356) );
  NAND2X0_LVT csr_add_x_381_U306 ( .A1(csr_add_x_381_n356), .A2(
        csr_add_x_381_n330), .Y(csr_add_x_381_n355) );
  AND2X1_LVT csr_add_x_381_U305 ( .A1(csr_add_x_381_n329), .A2(csr_n1941), .Y(
        csr_add_x_381_n354) );
  HADDX1_LVT csr_add_x_381_U304 ( .A0(csr_add_x_381_n354), .B0(csr_n1940), 
        .SO(csr_n_T_52[53]) );
  AND3X1_LVT csr_add_x_381_U303 ( .A1(csr_n1941), .A2(csr_n1940), .A3(
        csr_add_x_381_n329), .Y(csr_add_x_381_n351) );
  HADDX1_LVT csr_add_x_381_U302 ( .A0(csr_n1939), .B0(csr_add_x_381_n351), 
        .SO(csr_n_T_52[54]) );
  AND2X1_LVT csr_add_x_381_U301 ( .A1(csr_add_x_381_n351), .A2(csr_n1939), .Y(
        csr_add_x_381_n353) );
  HADDX1_LVT csr_add_x_381_U300 ( .A0(csr_add_x_381_n353), .B0(csr_n1938), 
        .SO(csr_n_T_52[55]) );
  AND3X1_LVT csr_add_x_381_U299 ( .A1(csr_n1938), .A2(csr_n1939), .A3(
        csr_add_x_381_n351), .Y(csr_add_x_381_n352) );
  HADDX1_LVT csr_add_x_381_U298 ( .A0(csr_add_x_381_n352), .B0(csr_n1937), 
        .SO(csr_n_T_52[56]) );
  AND4X1_LVT csr_add_x_381_U297 ( .A1(csr_n1938), .A2(csr_n1939), .A3(
        csr_add_x_381_n351), .A4(csr_n1937), .Y(csr_add_x_381_n350) );
  HADDX1_LVT csr_add_x_381_U296 ( .A0(csr_n1936), .B0(csr_add_x_381_n350), 
        .SO(csr_n_T_52[57]) );
  AND2X1_LVT csr_add_x_381_U295 ( .A1(csr_add_x_381_n344), .A2(csr_io_time[10]), .Y(csr_add_x_381_n349) );
  HADDX1_LVT csr_add_x_381_U294 ( .A0(csr_add_x_381_n349), .B0(csr_io_time[11]), .SO(csr_n_T_52[5]) );
  HADDX1_LVT csr_add_x_381_U293 ( .A0(csr_io_time[12]), .B0(csr_add_x_381_n348), .SO(csr_n_T_52[6]) );
  AND2X1_LVT csr_add_x_381_U292 ( .A1(csr_io_time[12]), .A2(csr_add_x_381_n348), .Y(csr_add_x_381_n347) );
  HADDX1_LVT csr_add_x_381_U291 ( .A0(csr_io_time[13]), .B0(csr_add_x_381_n347), .SO(csr_n_T_52[7]) );
  AO22X1_LVT csr_add_x_381_U290 ( .A1(csr_add_x_381_n342), .A2(
        csr_add_x_381_n341), .A3(csr_add_x_381_n346), .A4(csr_io_time[14]), 
        .Y(csr_n_T_52[8]) );
  AND2X1_LVT csr_add_x_381_U289 ( .A1(csr_io_time[14]), .A2(csr_add_x_381_n342), .Y(csr_add_x_381_n345) );
  HADDX1_LVT csr_add_x_381_U288 ( .A0(csr_add_x_381_n345), .B0(csr_io_time[15]), .SO(csr_n_T_52[9]) );
  INVX1_LVT csr_add_x_381_U287 ( .A(csr_add_x_381_n359), .Y(csr_add_x_381_n344) );
  INVX1_LVT csr_add_x_381_U286 ( .A(csr_add_x_381_n346), .Y(csr_add_x_381_n342) );
  INVX1_LVT csr_add_x_381_U285 ( .A(csr_add_x_381_n408), .Y(csr_add_x_381_n340) );
  INVX1_LVT csr_add_x_381_U284 ( .A(csr_add_x_381_n371), .Y(csr_add_x_381_n333) );
  INVX1_LVT csr_add_x_381_U283 ( .A(csr_add_x_381_n367), .Y(csr_add_x_381_n331) );
  INVX1_LVT csr_add_x_381_U282 ( .A(csr_add_x_381_n361), .Y(csr_add_x_381_n330) );
  INVX1_LVT csr_add_x_381_U281 ( .A(csr_add_x_381_n355), .Y(csr_add_x_381_n329) );
  INVX1_LVT csr_add_x_381_U280 ( .A(csr_add_x_381_n404), .Y(csr_add_x_381_n338) );
  INVX1_LVT csr_add_x_381_U279 ( .A(csr_add_x_381_n393), .Y(csr_add_x_381_n336) );
  INVX1_LVT csr_add_x_381_U278 ( .A(csr_add_x_381_n383), .Y(csr_add_x_381_n334) );
  INVX0_LVT csr_add_x_381_U277 ( .A(csr_n1953), .Y(csr_add_x_381_n332) );
  INVX1_LVT csr_add_x_381_U276 ( .A(csr_io_time[22]), .Y(csr_add_x_381_n337)
         );
  INVX1_LVT csr_add_x_381_U275 ( .A(csr_io_time[18]), .Y(csr_add_x_381_n339)
         );
  INVX1_LVT csr_add_x_381_U274 ( .A(csr_io_time[10]), .Y(csr_add_x_381_n343)
         );
  INVX1_LVT csr_add_x_381_U273 ( .A(csr_io_time[14]), .Y(csr_add_x_381_n341)
         );
  INVX1_LVT csr_add_x_381_U272 ( .A(csr_io_time[30]), .Y(csr_add_x_381_n335)
         );
  AO22X1_LVT csr_add_x_381_U271 ( .A1(csr_n1945), .A2(csr_add_x_381_n361), 
        .A3(csr_add_x_381_n328), .A4(csr_add_x_381_n330), .Y(csr_n_T_52[48])
         );
  INVX0_LVT csr_add_x_381_U270 ( .A(csr_n1945), .Y(csr_add_x_381_n328) );
  AO22X1_LVT csr_add_x_381_U269 ( .A1(csr_n1941), .A2(csr_add_x_381_n355), 
        .A3(csr_add_x_381_n327), .A4(csr_add_x_381_n329), .Y(csr_n_T_52[52])
         );
  INVX0_LVT csr_add_x_381_U268 ( .A(csr_n1941), .Y(csr_add_x_381_n327) );
  AO22X1_LVT csr_add_x_381_U267 ( .A1(csr_n1949), .A2(csr_add_x_381_n367), 
        .A3(csr_add_x_381_n326), .A4(csr_add_x_381_n331), .Y(csr_n_T_52[44])
         );
  INVX0_LVT csr_add_x_381_U266 ( .A(csr_n1949), .Y(csr_add_x_381_n326) );
  AO22X1_LVT csr_add_x_381_U265 ( .A1(csr_n1961), .A2(csr_add_x_381_n383), 
        .A3(csr_add_x_381_n325), .A4(csr_add_x_381_n334), .Y(csr_n_T_52[32])
         );
  INVX0_LVT csr_add_x_381_U264 ( .A(csr_n1961), .Y(csr_add_x_381_n325) );
  HADDX1_LVT csr_add_x_381_U259 ( .A0(csr_io_time[7]), .B0(csr_io_time[6]), 
        .C1(csr_add_x_381_n203), .SO(csr_n_T_52[1]) );
  NAND3X0_LVT csr_add_x_379_U406 ( .A1(csr_add_x_379_n203), .A2(csr_n_T_45_8_), 
        .A3(csr_n_T_45_9_), .Y(csr_add_x_379_n359) );
  AND3X1_LVT csr_add_x_379_U405 ( .A1(csr_n_T_45_10_), .A2(csr_n_T_45_11_), 
        .A3(csr_add_x_379_n344), .Y(csr_add_x_379_n348) );
  NAND3X0_LVT csr_add_x_379_U404 ( .A1(csr_n_T_45_12_), .A2(csr_n_T_45_13_), 
        .A3(csr_add_x_379_n348), .Y(csr_add_x_379_n346) );
  AND3X1_LVT csr_add_x_379_U403 ( .A1(csr_add_x_379_n342), .A2(csr_n_T_45_15_), 
        .A3(csr_n_T_45_14_), .Y(csr_add_x_379_n411) );
  HADDX1_LVT csr_add_x_379_U402 ( .A0(csr_n_T_45_16_), .B0(csr_add_x_379_n411), 
        .SO(csr_n_T_44[10]) );
  AND4X1_LVT csr_add_x_379_U401 ( .A1(csr_add_x_379_n342), .A2(csr_n_T_45_15_), 
        .A3(csr_n_T_45_14_), .A4(csr_n_T_45_16_), .Y(csr_add_x_379_n410) );
  HADDX1_LVT csr_add_x_379_U400 ( .A0(csr_n_T_45_17_), .B0(csr_add_x_379_n410), 
        .SO(csr_n_T_44[11]) );
  AND4X1_LVT csr_add_x_379_U399 ( .A1(csr_n_T_45_15_), .A2(csr_n_T_45_14_), 
        .A3(csr_n_T_45_17_), .A4(csr_n_T_45_16_), .Y(csr_add_x_379_n409) );
  NAND2X0_LVT csr_add_x_379_U398 ( .A1(csr_add_x_379_n342), .A2(
        csr_add_x_379_n409), .Y(csr_add_x_379_n408) );
  AO22X1_LVT csr_add_x_379_U397 ( .A1(csr_n_T_45_18_), .A2(csr_add_x_379_n408), 
        .A3(csr_add_x_379_n339), .A4(csr_add_x_379_n340), .Y(csr_n_T_44[12])
         );
  AND2X1_LVT csr_add_x_379_U396 ( .A1(csr_add_x_379_n340), .A2(csr_n_T_45_18_), 
        .Y(csr_add_x_379_n407) );
  HADDX1_LVT csr_add_x_379_U395 ( .A0(csr_add_x_379_n407), .B0(csr_n_T_45_19_), 
        .SO(csr_n_T_44[13]) );
  AND3X1_LVT csr_add_x_379_U394 ( .A1(csr_n_T_45_18_), .A2(csr_n_T_45_19_), 
        .A3(csr_add_x_379_n340), .Y(csr_add_x_379_n405) );
  HADDX1_LVT csr_add_x_379_U393 ( .A0(csr_n_T_45_20_), .B0(csr_add_x_379_n405), 
        .SO(csr_n_T_44[14]) );
  AND4X1_LVT csr_add_x_379_U392 ( .A1(csr_n_T_45_18_), .A2(csr_n_T_45_19_), 
        .A3(csr_n_T_45_20_), .A4(csr_add_x_379_n340), .Y(csr_add_x_379_n406)
         );
  HADDX1_LVT csr_add_x_379_U391 ( .A0(csr_n_T_45_21_), .B0(csr_add_x_379_n406), 
        .SO(csr_n_T_44[15]) );
  NAND3X0_LVT csr_add_x_379_U390 ( .A1(csr_n_T_45_20_), .A2(csr_n_T_45_21_), 
        .A3(csr_add_x_379_n405), .Y(csr_add_x_379_n404) );
  AO22X1_LVT csr_add_x_379_U389 ( .A1(csr_n_T_45_22_), .A2(csr_add_x_379_n404), 
        .A3(csr_add_x_379_n337), .A4(csr_add_x_379_n338), .Y(csr_n_T_44[16])
         );
  AND2X1_LVT csr_add_x_379_U388 ( .A1(csr_add_x_379_n338), .A2(csr_n_T_45_22_), 
        .Y(csr_add_x_379_n403) );
  HADDX1_LVT csr_add_x_379_U387 ( .A0(csr_add_x_379_n403), .B0(csr_n_T_45_23_), 
        .SO(csr_n_T_44[17]) );
  AND3X1_LVT csr_add_x_379_U386 ( .A1(csr_n_T_45_22_), .A2(csr_n_T_45_23_), 
        .A3(csr_add_x_379_n338), .Y(csr_add_x_379_n402) );
  HADDX1_LVT csr_add_x_379_U385 ( .A0(csr_n_T_45_24_), .B0(csr_add_x_379_n402), 
        .SO(csr_n_T_44[18]) );
  AND4X1_LVT csr_add_x_379_U384 ( .A1(csr_n_T_45_22_), .A2(csr_n_T_45_23_), 
        .A3(csr_n_T_45_24_), .A4(csr_add_x_379_n338), .Y(csr_add_x_379_n401)
         );
  HADDX1_LVT csr_add_x_379_U383 ( .A0(csr_n_T_45_25_), .B0(csr_add_x_379_n401), 
        .SO(csr_n_T_44[19]) );
  AND4X1_LVT csr_add_x_379_U382 ( .A1(csr_n_T_45_22_), .A2(csr_n_T_45_23_), 
        .A3(csr_n_T_45_25_), .A4(csr_n_T_45_24_), .Y(csr_add_x_379_n396) );
  AND2X1_LVT csr_add_x_379_U381 ( .A1(csr_add_x_379_n396), .A2(
        csr_add_x_379_n338), .Y(csr_add_x_379_n400) );
  HADDX1_LVT csr_add_x_379_U380 ( .A0(csr_n_T_45_26_), .B0(csr_add_x_379_n400), 
        .SO(csr_n_T_44[20]) );
  AND3X1_LVT csr_add_x_379_U379 ( .A1(csr_add_x_379_n396), .A2(csr_n_T_45_26_), 
        .A3(csr_add_x_379_n338), .Y(csr_add_x_379_n399) );
  HADDX1_LVT csr_add_x_379_U378 ( .A0(csr_add_x_379_n399), .B0(csr_n_T_45_27_), 
        .SO(csr_n_T_44[21]) );
  AND2X1_LVT csr_add_x_379_U377 ( .A1(csr_n_T_45_26_), .A2(csr_n_T_45_27_), 
        .Y(csr_add_x_379_n395) );
  AND3X1_LVT csr_add_x_379_U376 ( .A1(csr_add_x_379_n395), .A2(
        csr_add_x_379_n396), .A3(csr_add_x_379_n338), .Y(csr_add_x_379_n398)
         );
  HADDX1_LVT csr_add_x_379_U375 ( .A0(csr_n_T_45_28_), .B0(csr_add_x_379_n398), 
        .SO(csr_n_T_44[22]) );
  AND4X1_LVT csr_add_x_379_U374 ( .A1(csr_n_T_45_28_), .A2(csr_add_x_379_n395), 
        .A3(csr_add_x_379_n396), .A4(csr_add_x_379_n338), .Y(
        csr_add_x_379_n397) );
  HADDX1_LVT csr_add_x_379_U373 ( .A0(csr_n_T_45_29_), .B0(csr_add_x_379_n397), 
        .SO(csr_n_T_44[23]) );
  AND4X1_LVT csr_add_x_379_U372 ( .A1(csr_n_T_45_28_), .A2(csr_n_T_45_29_), 
        .A3(csr_add_x_379_n395), .A4(csr_add_x_379_n396), .Y(
        csr_add_x_379_n394) );
  NAND2X0_LVT csr_add_x_379_U371 ( .A1(csr_add_x_379_n394), .A2(
        csr_add_x_379_n338), .Y(csr_add_x_379_n393) );
  AO22X1_LVT csr_add_x_379_U370 ( .A1(csr_n_T_45_30_), .A2(csr_add_x_379_n393), 
        .A3(csr_add_x_379_n335), .A4(csr_add_x_379_n336), .Y(csr_n_T_44[24])
         );
  AND2X1_LVT csr_add_x_379_U369 ( .A1(csr_add_x_379_n336), .A2(csr_n_T_45_30_), 
        .Y(csr_add_x_379_n392) );
  HADDX1_LVT csr_add_x_379_U368 ( .A0(csr_add_x_379_n392), .B0(csr_n_T_45_31_), 
        .SO(csr_n_T_44[25]) );
  AND3X1_LVT csr_add_x_379_U367 ( .A1(csr_n_T_45_30_), .A2(csr_n_T_45_31_), 
        .A3(csr_add_x_379_n336), .Y(csr_add_x_379_n391) );
  HADDX1_LVT csr_add_x_379_U366 ( .A0(csr_n_T_45_32_), .B0(csr_add_x_379_n391), 
        .SO(csr_n_T_44[26]) );
  AND4X1_LVT csr_add_x_379_U365 ( .A1(csr_n_T_45_30_), .A2(csr_n_T_45_31_), 
        .A3(csr_n_T_45_32_), .A4(csr_add_x_379_n336), .Y(csr_add_x_379_n390)
         );
  HADDX1_LVT csr_add_x_379_U364 ( .A0(csr_n_T_45_33_), .B0(csr_add_x_379_n390), 
        .SO(csr_n_T_44[27]) );
  AND4X1_LVT csr_add_x_379_U363 ( .A1(csr_n_T_45_30_), .A2(csr_n_T_45_31_), 
        .A3(csr_n_T_45_33_), .A4(csr_n_T_45_32_), .Y(csr_add_x_379_n387) );
  AND2X1_LVT csr_add_x_379_U362 ( .A1(csr_add_x_379_n387), .A2(
        csr_add_x_379_n336), .Y(csr_add_x_379_n385) );
  HADDX1_LVT csr_add_x_379_U361 ( .A0(csr_n_T_45_34_), .B0(csr_add_x_379_n385), 
        .SO(csr_n_T_44[28]) );
  AND3X1_LVT csr_add_x_379_U360 ( .A1(csr_n_T_45_34_), .A2(csr_add_x_379_n387), 
        .A3(csr_add_x_379_n336), .Y(csr_add_x_379_n389) );
  HADDX1_LVT csr_add_x_379_U359 ( .A0(csr_add_x_379_n389), .B0(csr_n_T_45_35_), 
        .SO(csr_n_T_44[29]) );
  HADDX1_LVT csr_add_x_379_U358 ( .A0(csr_add_x_379_n203), .B0(csr_n_T_45_8_), 
        .SO(csr_n_T_44[2]) );
  AND2X1_LVT csr_add_x_379_U357 ( .A1(csr_n_T_45_34_), .A2(csr_n_T_45_35_), 
        .Y(csr_add_x_379_n384) );
  AND3X1_LVT csr_add_x_379_U356 ( .A1(csr_add_x_379_n387), .A2(
        csr_add_x_379_n384), .A3(csr_add_x_379_n336), .Y(csr_add_x_379_n388)
         );
  HADDX1_LVT csr_add_x_379_U355 ( .A0(csr_n_T_45_36_), .B0(csr_add_x_379_n388), 
        .SO(csr_n_T_44[30]) );
  AND4X1_LVT csr_add_x_379_U354 ( .A1(csr_add_x_379_n387), .A2(csr_n_T_45_36_), 
        .A3(csr_add_x_379_n384), .A4(csr_add_x_379_n336), .Y(
        csr_add_x_379_n386) );
  HADDX1_LVT csr_add_x_379_U353 ( .A0(csr_n_T_45_37_), .B0(csr_add_x_379_n386), 
        .SO(csr_n_T_44[31]) );
  NAND4X0_LVT csr_add_x_379_U352 ( .A1(csr_n_T_45_37_), .A2(csr_n_T_45_36_), 
        .A3(csr_add_x_379_n384), .A4(csr_add_x_379_n385), .Y(
        csr_add_x_379_n383) );
  AND2X1_LVT csr_add_x_379_U351 ( .A1(csr_n_T_45_38_), .A2(csr_add_x_379_n334), 
        .Y(csr_add_x_379_n382) );
  HADDX1_LVT csr_add_x_379_U350 ( .A0(csr_add_x_379_n382), .B0(csr_n_T_45_39_), 
        .SO(csr_n_T_44[33]) );
  AND3X1_LVT csr_add_x_379_U349 ( .A1(csr_add_x_379_n334), .A2(csr_n_T_45_38_), 
        .A3(csr_n_T_45_39_), .Y(csr_add_x_379_n381) );
  HADDX1_LVT csr_add_x_379_U348 ( .A0(csr_n_T_45_40_), .B0(csr_add_x_379_n381), 
        .SO(csr_n_T_44[34]) );
  AND4X1_LVT csr_add_x_379_U347 ( .A1(csr_add_x_379_n334), .A2(csr_n_T_45_38_), 
        .A3(csr_n_T_45_39_), .A4(csr_n_T_45_40_), .Y(csr_add_x_379_n380) );
  HADDX1_LVT csr_add_x_379_U346 ( .A0(csr_n_T_45_41_), .B0(csr_add_x_379_n380), 
        .SO(csr_n_T_44[35]) );
  AND4X1_LVT csr_add_x_379_U345 ( .A1(csr_n_T_45_38_), .A2(csr_n_T_45_39_), 
        .A3(csr_n_T_45_41_), .A4(csr_n_T_45_40_), .Y(csr_add_x_379_n374) );
  AND2X1_LVT csr_add_x_379_U344 ( .A1(csr_add_x_379_n334), .A2(
        csr_add_x_379_n374), .Y(csr_add_x_379_n379) );
  HADDX1_LVT csr_add_x_379_U343 ( .A0(csr_n_T_45_42_), .B0(csr_add_x_379_n379), 
        .SO(csr_n_T_44[36]) );
  AND3X1_LVT csr_add_x_379_U342 ( .A1(csr_n_T_45_42_), .A2(csr_add_x_379_n334), 
        .A3(csr_add_x_379_n374), .Y(csr_add_x_379_n378) );
  HADDX1_LVT csr_add_x_379_U341 ( .A0(csr_add_x_379_n378), .B0(csr_n_T_45_43_), 
        .SO(csr_n_T_44[37]) );
  AND2X1_LVT csr_add_x_379_U340 ( .A1(csr_n_T_45_42_), .A2(csr_n_T_45_43_), 
        .Y(csr_add_x_379_n373) );
  AND3X1_LVT csr_add_x_379_U339 ( .A1(csr_add_x_379_n334), .A2(
        csr_add_x_379_n373), .A3(csr_add_x_379_n374), .Y(csr_add_x_379_n377)
         );
  HADDX1_LVT csr_add_x_379_U338 ( .A0(csr_n_T_45_44_), .B0(csr_add_x_379_n377), 
        .SO(csr_n_T_44[38]) );
  AND4X1_LVT csr_add_x_379_U337 ( .A1(csr_add_x_379_n334), .A2(csr_n_T_45_44_), 
        .A3(csr_add_x_379_n373), .A4(csr_add_x_379_n374), .Y(
        csr_add_x_379_n376) );
  HADDX1_LVT csr_add_x_379_U336 ( .A0(csr_n_T_45_45_), .B0(csr_add_x_379_n376), 
        .SO(csr_n_T_44[39]) );
  AND2X1_LVT csr_add_x_379_U335 ( .A1(csr_add_x_379_n203), .A2(csr_n_T_45_8_), 
        .Y(csr_add_x_379_n375) );
  HADDX1_LVT csr_add_x_379_U334 ( .A0(csr_n_T_45_9_), .B0(csr_add_x_379_n375), 
        .SO(csr_n_T_44[3]) );
  AND4X1_LVT csr_add_x_379_U333 ( .A1(csr_n_T_45_44_), .A2(csr_n_T_45_45_), 
        .A3(csr_add_x_379_n373), .A4(csr_add_x_379_n374), .Y(
        csr_add_x_379_n372) );
  NAND2X0_LVT csr_add_x_379_U332 ( .A1(csr_add_x_379_n334), .A2(
        csr_add_x_379_n372), .Y(csr_add_x_379_n371) );
  AO22X1_LVT csr_add_x_379_U331 ( .A1(csr_n_T_45_46_), .A2(csr_add_x_379_n371), 
        .A3(csr_add_x_379_n332), .A4(csr_add_x_379_n333), .Y(csr_n_T_44[40])
         );
  AND2X1_LVT csr_add_x_379_U330 ( .A1(csr_add_x_379_n333), .A2(csr_n_T_45_46_), 
        .Y(csr_add_x_379_n370) );
  HADDX1_LVT csr_add_x_379_U329 ( .A0(csr_add_x_379_n370), .B0(csr_n_T_45_47_), 
        .SO(csr_n_T_44[41]) );
  AND3X1_LVT csr_add_x_379_U328 ( .A1(csr_n_T_45_46_), .A2(csr_n_T_45_47_), 
        .A3(csr_add_x_379_n333), .Y(csr_add_x_379_n369) );
  HADDX1_LVT csr_add_x_379_U327 ( .A0(csr_n_T_45_48_), .B0(csr_add_x_379_n369), 
        .SO(csr_n_T_44[42]) );
  AND4X1_LVT csr_add_x_379_U326 ( .A1(csr_n_T_45_46_), .A2(csr_n_T_45_47_), 
        .A3(csr_n_T_45_48_), .A4(csr_add_x_379_n333), .Y(csr_add_x_379_n368)
         );
  HADDX1_LVT csr_add_x_379_U325 ( .A0(csr_n_T_45_49_), .B0(csr_add_x_379_n368), 
        .SO(csr_n_T_44[43]) );
  AND4X1_LVT csr_add_x_379_U324 ( .A1(csr_n_T_45_46_), .A2(csr_n_T_45_47_), 
        .A3(csr_n_T_45_49_), .A4(csr_n_T_45_48_), .Y(csr_add_x_379_n363) );
  NAND2X0_LVT csr_add_x_379_U323 ( .A1(csr_add_x_379_n363), .A2(
        csr_add_x_379_n333), .Y(csr_add_x_379_n367) );
  AND2X1_LVT csr_add_x_379_U322 ( .A1(csr_add_x_379_n331), .A2(csr_n_T_45_50_), 
        .Y(csr_add_x_379_n366) );
  HADDX1_LVT csr_add_x_379_U321 ( .A0(csr_add_x_379_n366), .B0(csr_n_T_45_51_), 
        .SO(csr_n_T_44[45]) );
  AND3X1_LVT csr_add_x_379_U320 ( .A1(csr_n_T_45_50_), .A2(csr_n_T_45_51_), 
        .A3(csr_add_x_379_n331), .Y(csr_add_x_379_n365) );
  HADDX1_LVT csr_add_x_379_U319 ( .A0(csr_n_T_45_52_), .B0(csr_add_x_379_n365), 
        .SO(csr_n_T_44[46]) );
  AND4X1_LVT csr_add_x_379_U318 ( .A1(csr_n_T_45_52_), .A2(csr_n_T_45_50_), 
        .A3(csr_n_T_45_51_), .A4(csr_add_x_379_n331), .Y(csr_add_x_379_n364)
         );
  HADDX1_LVT csr_add_x_379_U317 ( .A0(csr_n_T_45_53_), .B0(csr_add_x_379_n364), 
        .SO(csr_n_T_44[47]) );
  AND4X1_LVT csr_add_x_379_U316 ( .A1(csr_n_T_45_50_), .A2(csr_n_T_45_51_), 
        .A3(csr_add_x_379_n363), .A4(csr_add_x_379_n333), .Y(
        csr_add_x_379_n362) );
  NAND3X0_LVT csr_add_x_379_U315 ( .A1(csr_n_T_45_53_), .A2(csr_n_T_45_52_), 
        .A3(csr_add_x_379_n362), .Y(csr_add_x_379_n361) );
  AO22X1_LVT csr_add_x_379_U314 ( .A1(csr_n_T_45_54_), .A2(csr_add_x_379_n361), 
        .A3(csr_add_x_379_n329), .A4(csr_add_x_379_n330), .Y(csr_n_T_44[48])
         );
  AND2X1_LVT csr_add_x_379_U313 ( .A1(csr_add_x_379_n330), .A2(csr_n_T_45_54_), 
        .Y(csr_add_x_379_n360) );
  HADDX1_LVT csr_add_x_379_U312 ( .A0(csr_add_x_379_n360), .B0(csr_n_T_45_55_), 
        .SO(csr_n_T_44[49]) );
  AO22X1_LVT csr_add_x_379_U311 ( .A1(csr_n_T_45_10_), .A2(csr_add_x_379_n359), 
        .A3(csr_add_x_379_n343), .A4(csr_add_x_379_n344), .Y(csr_n_T_44[4]) );
  AND3X1_LVT csr_add_x_379_U310 ( .A1(csr_n_T_45_54_), .A2(csr_n_T_45_55_), 
        .A3(csr_add_x_379_n330), .Y(csr_add_x_379_n358) );
  HADDX1_LVT csr_add_x_379_U309 ( .A0(csr_n_T_45_56_), .B0(csr_add_x_379_n358), 
        .SO(csr_n_T_44[50]) );
  AND4X1_LVT csr_add_x_379_U308 ( .A1(csr_n_T_45_54_), .A2(csr_n_T_45_55_), 
        .A3(csr_n_T_45_56_), .A4(csr_add_x_379_n330), .Y(csr_add_x_379_n357)
         );
  HADDX1_LVT csr_add_x_379_U307 ( .A0(csr_n_T_45_57_), .B0(csr_add_x_379_n357), 
        .SO(csr_n_T_44[51]) );
  AND4X1_LVT csr_add_x_379_U306 ( .A1(csr_n_T_45_54_), .A2(csr_n_T_45_55_), 
        .A3(csr_n_T_45_57_), .A4(csr_n_T_45_56_), .Y(csr_add_x_379_n356) );
  NAND2X0_LVT csr_add_x_379_U305 ( .A1(csr_add_x_379_n356), .A2(
        csr_add_x_379_n330), .Y(csr_add_x_379_n355) );
  AND2X1_LVT csr_add_x_379_U304 ( .A1(csr_add_x_379_n328), .A2(csr_n_T_45_58_), 
        .Y(csr_add_x_379_n354) );
  HADDX1_LVT csr_add_x_379_U303 ( .A0(csr_add_x_379_n354), .B0(csr_n_T_45_59_), 
        .SO(csr_n_T_44[53]) );
  AND3X1_LVT csr_add_x_379_U302 ( .A1(csr_n_T_45_58_), .A2(csr_n_T_45_59_), 
        .A3(csr_add_x_379_n328), .Y(csr_add_x_379_n351) );
  HADDX1_LVT csr_add_x_379_U301 ( .A0(csr_n_T_45_60_), .B0(csr_add_x_379_n351), 
        .SO(csr_n_T_44[54]) );
  AND2X1_LVT csr_add_x_379_U300 ( .A1(csr_add_x_379_n351), .A2(csr_n_T_45_60_), 
        .Y(csr_add_x_379_n353) );
  HADDX1_LVT csr_add_x_379_U299 ( .A0(csr_add_x_379_n353), .B0(csr_n_T_45_61_), 
        .SO(csr_n_T_44[55]) );
  AND3X1_LVT csr_add_x_379_U298 ( .A1(csr_n_T_45_61_), .A2(csr_n_T_45_60_), 
        .A3(csr_add_x_379_n351), .Y(csr_add_x_379_n352) );
  HADDX1_LVT csr_add_x_379_U297 ( .A0(csr_add_x_379_n352), .B0(csr_n_T_45_62_), 
        .SO(csr_n_T_44[56]) );
  AND4X1_LVT csr_add_x_379_U296 ( .A1(csr_n_T_45_61_), .A2(csr_n_T_45_60_), 
        .A3(csr_add_x_379_n351), .A4(csr_n_T_45_62_), .Y(csr_add_x_379_n350)
         );
  HADDX1_LVT csr_add_x_379_U295 ( .A0(csr_n_T_45_63_), .B0(csr_add_x_379_n350), 
        .SO(csr_n_T_44[57]) );
  AND2X1_LVT csr_add_x_379_U294 ( .A1(csr_add_x_379_n344), .A2(csr_n_T_45_10_), 
        .Y(csr_add_x_379_n349) );
  HADDX1_LVT csr_add_x_379_U293 ( .A0(csr_add_x_379_n349), .B0(csr_n_T_45_11_), 
        .SO(csr_n_T_44[5]) );
  HADDX1_LVT csr_add_x_379_U292 ( .A0(csr_n_T_45_12_), .B0(csr_add_x_379_n348), 
        .SO(csr_n_T_44[6]) );
  AND2X1_LVT csr_add_x_379_U291 ( .A1(csr_n_T_45_12_), .A2(csr_add_x_379_n348), 
        .Y(csr_add_x_379_n347) );
  HADDX1_LVT csr_add_x_379_U290 ( .A0(csr_n_T_45_13_), .B0(csr_add_x_379_n347), 
        .SO(csr_n_T_44[7]) );
  AO22X1_LVT csr_add_x_379_U289 ( .A1(csr_add_x_379_n342), .A2(
        csr_add_x_379_n341), .A3(csr_add_x_379_n346), .A4(csr_n_T_45_14_), .Y(
        csr_n_T_44[8]) );
  AND2X1_LVT csr_add_x_379_U288 ( .A1(csr_n_T_45_14_), .A2(csr_add_x_379_n342), 
        .Y(csr_add_x_379_n345) );
  HADDX1_LVT csr_add_x_379_U287 ( .A0(csr_add_x_379_n345), .B0(csr_n_T_45_15_), 
        .SO(csr_n_T_44[9]) );
  INVX1_LVT csr_add_x_379_U286 ( .A(csr_add_x_379_n359), .Y(csr_add_x_379_n344) );
  INVX1_LVT csr_add_x_379_U285 ( .A(csr_n_T_45_10_), .Y(csr_add_x_379_n343) );
  INVX1_LVT csr_add_x_379_U284 ( .A(csr_add_x_379_n346), .Y(csr_add_x_379_n342) );
  INVX1_LVT csr_add_x_379_U283 ( .A(csr_add_x_379_n408), .Y(csr_add_x_379_n340) );
  INVX1_LVT csr_add_x_379_U282 ( .A(csr_n_T_45_18_), .Y(csr_add_x_379_n339) );
  INVX1_LVT csr_add_x_379_U281 ( .A(csr_n_T_45_22_), .Y(csr_add_x_379_n337) );
  INVX1_LVT csr_add_x_379_U280 ( .A(csr_add_x_379_n371), .Y(csr_add_x_379_n333) );
  INVX1_LVT csr_add_x_379_U279 ( .A(csr_add_x_379_n367), .Y(csr_add_x_379_n331) );
  INVX1_LVT csr_add_x_379_U278 ( .A(csr_add_x_379_n361), .Y(csr_add_x_379_n330) );
  INVX1_LVT csr_add_x_379_U277 ( .A(csr_add_x_379_n355), .Y(csr_add_x_379_n328) );
  INVX1_LVT csr_add_x_379_U276 ( .A(csr_add_x_379_n404), .Y(csr_add_x_379_n338) );
  INVX1_LVT csr_add_x_379_U275 ( .A(csr_add_x_379_n393), .Y(csr_add_x_379_n336) );
  INVX1_LVT csr_add_x_379_U274 ( .A(csr_add_x_379_n383), .Y(csr_add_x_379_n334) );
  INVX0_LVT csr_add_x_379_U273 ( .A(csr_n_T_45_46_), .Y(csr_add_x_379_n332) );
  INVX0_LVT csr_add_x_379_U272 ( .A(csr_n_T_45_54_), .Y(csr_add_x_379_n329) );
  INVX0_LVT csr_add_x_379_U271 ( .A(csr_n_T_45_14_), .Y(csr_add_x_379_n341) );
  INVX0_LVT csr_add_x_379_U270 ( .A(csr_n_T_45_30_), .Y(csr_add_x_379_n335) );
  AO22X1_LVT csr_add_x_379_U269 ( .A1(csr_n_T_45_38_), .A2(csr_add_x_379_n383), 
        .A3(csr_add_x_379_n327), .A4(csr_add_x_379_n334), .Y(csr_n_T_44[32])
         );
  INVX0_LVT csr_add_x_379_U268 ( .A(csr_n_T_45_38_), .Y(csr_add_x_379_n327) );
  AO22X1_LVT csr_add_x_379_U267 ( .A1(csr_n_T_45_50_), .A2(csr_add_x_379_n367), 
        .A3(csr_add_x_379_n326), .A4(csr_add_x_379_n331), .Y(csr_n_T_44[44])
         );
  INVX0_LVT csr_add_x_379_U266 ( .A(csr_n_T_45_50_), .Y(csr_add_x_379_n326) );
  AO22X1_LVT csr_add_x_379_U265 ( .A1(csr_n_T_45_58_), .A2(csr_add_x_379_n355), 
        .A3(csr_add_x_379_n325), .A4(csr_add_x_379_n328), .Y(csr_n_T_44[52])
         );
  INVX0_LVT csr_add_x_379_U264 ( .A(csr_n_T_45_58_), .Y(csr_add_x_379_n325) );
  HADDX1_LVT csr_add_x_379_U259 ( .A0(csr_n_T_45_7_), .B0(csr_n_T_45_6_), .C1(
        csr_add_x_379_n203), .SO(csr_n_T_44[1]) );
  AND3X1_LVT bpu_U173 ( .A1(bpu_n166), .A2(csr_io_bp_0_control_w), .A3(bpu_n69), .Y(bpu_io_xcpt_st) );
  AND2X1_LVT bpu_U172 ( .A1(bpu_n165), .A2(bpu_n69), .Y(bpu_io_xcpt_ld) );
  AND3X1_LVT bpu_U171 ( .A1(csr_io_bp_0_control_action), .A2(bpu_n166), .A3(
        csr_io_bp_0_control_w), .Y(bpu_io_debug_st) );
  AND2X1_LVT bpu_U170 ( .A1(csr_io_bp_0_control_action), .A2(bpu_n165), .Y(
        bpu_io_debug_ld) );
  AND2X1_LVT bpu_U169 ( .A1(bpu_n166), .A2(csr_io_bp_0_control_r), .Y(bpu_n165) );
  OA221X1_LVT bpu_U168 ( .A1(csr_io_bp_0_control_tmatch[1]), .A2(bpu_n164), 
        .A3(bpu_n163), .A4(bpu_n162), .A5(bpu_n67), .Y(bpu_n166) );
  AO22X1_LVT bpu_U167 ( .A1(csr_io_bp_0_control_tmatch[0]), .A2(bpu_n161), 
        .A3(bpu_n70), .A4(bpu_n_T_9), .Y(bpu_n162) );
  OA221X1_LVT bpu_U166 ( .A1(bpu_n148), .A2(n_T_918[6]), .A3(bpu_n147), .A4(
        n_T_918[7]), .A5(bpu_n146), .Y(bpu_n149) );
  AOI22X1_LVT bpu_U165 ( .A1(bpu_n148), .A2(n_T_918[6]), .A3(bpu_n147), .A4(
        n_T_918[7]), .Y(bpu_n146) );
  OA221X1_LVT bpu_U164 ( .A1(bpu_n145), .A2(n_T_918[8]), .A3(bpu_n144), .A4(
        n_T_918[14]), .A5(bpu_n143), .Y(bpu_n150) );
  AOI22X1_LVT bpu_U163 ( .A1(bpu_n144), .A2(n_T_918[14]), .A3(bpu_n145), .A4(
        n_T_918[8]), .Y(bpu_n143) );
  OA221X1_LVT bpu_U162 ( .A1(bpu_n142), .A2(n_T_918[11]), .A3(bpu_n141), .A4(
        n_T_918[17]), .A5(bpu_n140), .Y(bpu_n151) );
  AOI22X1_LVT bpu_U161 ( .A1(bpu_n142), .A2(n_T_918[11]), .A3(bpu_n141), .A4(
        n_T_918[17]), .Y(bpu_n140) );
  OA221X1_LVT bpu_U160 ( .A1(bpu_n139), .A2(n_T_918[24]), .A3(bpu_n138), .A4(
        n_T_918[21]), .A5(bpu_n137), .Y(bpu_n152) );
  AOI22X1_LVT bpu_U159 ( .A1(bpu_n138), .A2(n_T_918[21]), .A3(bpu_n139), .A4(
        n_T_918[24]), .Y(bpu_n137) );
  AO221X1_LVT bpu_U158 ( .A1(csr_io_bp_0_address[2]), .A2(bpu_n136), .A3(
        bpu_n135), .A4(n_T_918[2]), .A5(bpu_n134), .Y(bpu_n153) );
  OA222X1_LVT bpu_U157 ( .A1(csr_io_bp_0_address[1]), .A2(n_T_918[1]), .A3(
        bpu_n133), .A4(bpu_n132), .A5(bpu_n70), .A6(bpu_n131), .Y(bpu_n134) );
  OA221X1_LVT bpu_U156 ( .A1(bpu_n126), .A2(n_T_918[29]), .A3(bpu_n125), .A4(
        n_T_918[28]), .A5(bpu_n124), .Y(bpu_n127) );
  AOI22X1_LVT bpu_U155 ( .A1(bpu_n126), .A2(n_T_918[29]), .A3(bpu_n125), .A4(
        n_T_918[28]), .Y(bpu_n124) );
  OA221X1_LVT bpu_U154 ( .A1(bpu_n123), .A2(n_T_918[37]), .A3(bpu_n122), .A4(
        n_T_918[27]), .A5(bpu_n121), .Y(bpu_n128) );
  AOI22X1_LVT bpu_U153 ( .A1(bpu_n122), .A2(n_T_918[27]), .A3(bpu_n123), .A4(
        n_T_918[37]), .Y(bpu_n121) );
  OA221X1_LVT bpu_U152 ( .A1(bpu_n120), .A2(n_T_918[5]), .A3(bpu_n119), .A4(
        n_T_918[4]), .A5(bpu_n118), .Y(bpu_n129) );
  AOI22X1_LVT bpu_U151 ( .A1(bpu_n120), .A2(n_T_918[5]), .A3(bpu_n119), .A4(
        n_T_918[4]), .Y(bpu_n118) );
  OA221X1_LVT bpu_U150 ( .A1(bpu_n117), .A2(n_T_918[12]), .A3(bpu_n116), .A4(
        n_T_918[15]), .A5(bpu_n115), .Y(bpu_n130) );
  AOI22X1_LVT bpu_U149 ( .A1(bpu_n117), .A2(n_T_918[12]), .A3(bpu_n116), .A4(
        n_T_918[15]), .Y(bpu_n115) );
  NAND4X0_LVT bpu_U148 ( .A1(bpu_n114), .A2(bpu_n113), .A3(bpu_n112), .A4(
        bpu_n111), .Y(bpu_n156) );
  OA221X1_LVT bpu_U147 ( .A1(bpu_n110), .A2(n_T_918[16]), .A3(bpu_n109), .A4(
        n_T_918[20]), .A5(bpu_n108), .Y(bpu_n111) );
  AOI22X1_LVT bpu_U146 ( .A1(bpu_n109), .A2(n_T_918[20]), .A3(bpu_n110), .A4(
        n_T_918[16]), .Y(bpu_n108) );
  OA221X1_LVT bpu_U145 ( .A1(bpu_n107), .A2(n_T_918[19]), .A3(bpu_n106), .A4(
        n_T_918[38]), .A5(bpu_n105), .Y(bpu_n112) );
  AOI22X1_LVT bpu_U144 ( .A1(bpu_n107), .A2(n_T_918[19]), .A3(bpu_n106), .A4(
        n_T_918[38]), .Y(bpu_n105) );
  OA221X1_LVT bpu_U143 ( .A1(bpu_n104), .A2(n_T_918[34]), .A3(bpu_n103), .A4(
        n_T_918[32]), .A5(bpu_n102), .Y(bpu_n113) );
  AOI22X1_LVT bpu_U142 ( .A1(bpu_n104), .A2(n_T_918[34]), .A3(bpu_n103), .A4(
        n_T_918[32]), .Y(bpu_n102) );
  OA221X1_LVT bpu_U141 ( .A1(bpu_n101), .A2(n_T_918[31]), .A3(bpu_n100), .A4(
        n_T_918[30]), .A5(bpu_n99), .Y(bpu_n114) );
  AOI22X1_LVT bpu_U140 ( .A1(bpu_n101), .A2(n_T_918[31]), .A3(bpu_n100), .A4(
        n_T_918[30]), .Y(bpu_n99) );
  NAND4X0_LVT bpu_U139 ( .A1(bpu_n98), .A2(bpu_n97), .A3(bpu_n96), .A4(bpu_n95), .Y(bpu_n159) );
  OA221X1_LVT bpu_U138 ( .A1(bpu_n94), .A2(n_T_918[18]), .A3(bpu_n93), .A4(
        n_T_918[13]), .A5(bpu_n92), .Y(bpu_n95) );
  AOI22X1_LVT bpu_U137 ( .A1(bpu_n94), .A2(n_T_918[18]), .A3(bpu_n93), .A4(
        n_T_918[13]), .Y(bpu_n92) );
  OA221X1_LVT bpu_U136 ( .A1(bpu_n91), .A2(n_T_918[25]), .A3(bpu_n90), .A4(
        n_T_918[10]), .A5(bpu_n89), .Y(bpu_n96) );
  AOI22X1_LVT bpu_U135 ( .A1(bpu_n91), .A2(n_T_918[25]), .A3(bpu_n90), .A4(
        n_T_918[10]), .Y(bpu_n89) );
  OA221X1_LVT bpu_U134 ( .A1(bpu_n88), .A2(n_T_918[35]), .A3(bpu_n87), .A4(
        n_T_918[36]), .A5(bpu_n86), .Y(bpu_n97) );
  AOI22X1_LVT bpu_U133 ( .A1(bpu_n87), .A2(n_T_918[36]), .A3(bpu_n88), .A4(
        n_T_918[35]), .Y(bpu_n86) );
  OA221X1_LVT bpu_U132 ( .A1(bpu_n85), .A2(n_T_918[9]), .A3(bpu_n84), .A4(
        n_T_918[23]), .A5(bpu_n83), .Y(bpu_n98) );
  AOI22X1_LVT bpu_U131 ( .A1(bpu_n84), .A2(n_T_918[23]), .A3(bpu_n85), .A4(
        n_T_918[9]), .Y(bpu_n83) );
  NAND3X0_LVT bpu_U130 ( .A1(bpu_n82), .A2(bpu_n81), .A3(bpu_n80), .Y(bpu_n160) );
  AO222X1_LVT bpu_U129 ( .A1(csr_io_bp_0_address[3]), .A2(n_T_918[3]), .A3(
        bpu_n79), .A4(bpu_n78), .A5(bpu_n68), .A6(csr_io_bp_0_address[2]), .Y(
        bpu_n80) );
  OA222X1_LVT bpu_U128 ( .A1(csr_io_bp_0_address[22]), .A2(bpu_n77), .A3(
        bpu_n76), .A4(n_T_918[22]), .A5(csr_io_bp_0_control_tmatch[0]), .A6(
        bpu_n75), .Y(bpu_n81) );
  AO22X1_LVT bpu_U127 ( .A1(csr_io_bp_0_address[0]), .A2(n_T_918[0]), .A3(
        bpu_n131), .A4(bpu_n74), .Y(bpu_n75) );
  OA221X1_LVT bpu_U126 ( .A1(bpu_n73), .A2(n_T_918[33]), .A3(bpu_n72), .A4(
        n_T_918[26]), .A5(bpu_n71), .Y(bpu_n82) );
  AOI22X1_LVT bpu_U125 ( .A1(bpu_n73), .A2(n_T_918[33]), .A3(bpu_n72), .A4(
        n_T_918[26]), .Y(bpu_n71) );
  AND2X1_LVT bpu_U122 ( .A1(bpu_n66), .A2(bpu_n69), .Y(bpu_io_xcpt_if) );
  AND2X1_LVT bpu_U121 ( .A1(bpu_n66), .A2(csr_io_bp_0_control_action), .Y(
        bpu_io_debug_if) );
  AND3X1_LVT bpu_U120 ( .A1(bpu_n65), .A2(bpu_n67), .A3(csr_io_bp_0_control_x), 
        .Y(bpu_n66) );
  MUX21X1_LVT bpu_U119 ( .A1(bpu_n64), .A2(bpu_n63), .S0(
        csr_io_bp_0_control_tmatch[1]), .Y(bpu_n65) );
  NOR4X1_LVT bpu_U118 ( .A1(bpu_n62), .A2(bpu_n61), .A3(bpu_n60), .A4(bpu_n59), 
        .Y(bpu_n64) );
  NAND4X0_LVT bpu_U117 ( .A1(bpu_n58), .A2(bpu_n57), .A3(bpu_n56), .A4(bpu_n55), .Y(bpu_n59) );
  AND4X1_LVT bpu_U116 ( .A1(bpu_n54), .A2(bpu_n53), .A3(bpu_n52), .A4(bpu_n51), 
        .Y(bpu_n55) );
  OA22X1_LVT bpu_U115 ( .A1(bpu_n68), .A2(bpu_n50), .A3(
        csr_io_bp_0_control_tmatch[0]), .A4(bpu_n49), .Y(bpu_n56) );
  AND4X1_LVT bpu_U114 ( .A1(bpu_n48), .A2(bpu_n47), .A3(bpu_n46), .A4(bpu_n45), 
        .Y(bpu_n57) );
  AO21X1_LVT bpu_U113 ( .A1(csr_io_bp_0_address[2]), .A2(bpu_n68), .A3(bpu_n44), .Y(bpu_n48) );
  NOR4X1_LVT bpu_U112 ( .A1(bpu_n43), .A2(bpu_n42), .A3(bpu_n41), .A4(bpu_n40), 
        .Y(bpu_n58) );
  NAND4X0_LVT bpu_U111 ( .A1(bpu_n39), .A2(bpu_n38), .A3(bpu_n37), .A4(bpu_n36), .Y(bpu_n40) );
  NAND4X0_LVT bpu_U110 ( .A1(bpu_n35), .A2(bpu_n34), .A3(bpu_n33), .A4(bpu_n32), .Y(bpu_n41) );
  NAND4X0_LVT bpu_U109 ( .A1(bpu_n31), .A2(bpu_n30), .A3(bpu_n29), .A4(bpu_n28), .Y(bpu_n42) );
  NAND4X0_LVT bpu_U108 ( .A1(bpu_n27), .A2(bpu_n26), .A3(bpu_n25), .A4(bpu_n24), .Y(bpu_n43) );
  AO21X1_LVT bpu_U107 ( .A1(bpu_n23), .A2(bpu_n22), .A3(bpu_n21), .Y(bpu_n60)
         );
  NAND4X0_LVT bpu_U106 ( .A1(bpu_n20), .A2(bpu_n19), .A3(bpu_n18), .A4(bpu_n17), .Y(bpu_n21) );
  INVX1_LVT bpu_U105 ( .A(bpu_n16), .Y(bpu_n22) );
  NAND4X0_LVT bpu_U104 ( .A1(bpu_n15), .A2(bpu_n14), .A3(bpu_n13), .A4(bpu_n12), .Y(bpu_n61) );
  NAND4X0_LVT bpu_U103 ( .A1(bpu_n11), .A2(bpu_n10), .A3(bpu_n9), .A4(bpu_n8), 
        .Y(bpu_n62) );
  INVX1_LVT bpu_U102 ( .A(csr_io_bp_0_control_action), .Y(bpu_n69) );
  INVX1_LVT bpu_U101 ( .A(csr_io_bp_0_address[7]), .Y(bpu_n147) );
  INVX1_LVT bpu_U100 ( .A(csr_io_bp_0_address[15]), .Y(bpu_n116) );
  INVX1_LVT bpu_U99 ( .A(csr_io_bp_0_address[13]), .Y(bpu_n93) );
  INVX1_LVT bpu_U98 ( .A(csr_io_bp_0_address[18]), .Y(bpu_n94) );
  INVX1_LVT bpu_U97 ( .A(csr_io_bp_0_address[9]), .Y(bpu_n85) );
  AND2X1_LVT bpu_U96 ( .A1(bpu_n16), .A2(csr_io_bp_0_address[1]), .Y(bpu_n68)
         );
  AND2X1_LVT bpu_U95 ( .A1(csr_io_bp_0_address[0]), .A2(
        csr_io_bp_0_control_tmatch[0]), .Y(bpu_n16) );
  INVX1_LVT bpu_U94 ( .A(csr_io_bp_0_address[0]), .Y(bpu_n131) );
  NAND3X0_LVT bpu_U93 ( .A1(bpu_n5), .A2(bpu_n6), .A3(bpu_n7), .Y(bpu_n155) );
  NAND2X0_LVT bpu_U92 ( .A1(bpu_n154), .A2(bpu_n153), .Y(bpu_n7) );
  AND4X1_LVT bpu_U91 ( .A1(bpu_n130), .A2(bpu_n129), .A3(bpu_n128), .A4(
        bpu_n127), .Y(bpu_n6) );
  AND4X1_LVT bpu_U90 ( .A1(bpu_n152), .A2(bpu_n151), .A3(bpu_n150), .A4(
        bpu_n149), .Y(bpu_n5) );
  XOR2X1_LVT bpu_U89 ( .A1(ibuf_io_pc[26]), .A2(bpu_n72), .Y(bpu_n19) );
  XOR2X1_LVT bpu_U88 ( .A1(ibuf_io_pc[32]), .A2(bpu_n103), .Y(bpu_n26) );
  XOR2X1_LVT bpu_U87 ( .A1(ibuf_io_pc[30]), .A2(bpu_n100), .Y(bpu_n25) );
  XOR2X1_LVT bpu_U86 ( .A1(ibuf_io_pc[16]), .A2(bpu_n110), .Y(bpu_n24) );
  XOR2X1_LVT bpu_U85 ( .A1(ibuf_io_pc[19]), .A2(bpu_n107), .Y(bpu_n31) );
  XOR2X1_LVT bpu_U84 ( .A1(ibuf_io_pc[8]), .A2(bpu_n145), .Y(bpu_n29) );
  XOR2X1_LVT bpu_U83 ( .A1(ibuf_io_pc[25]), .A2(bpu_n91), .Y(bpu_n28) );
  XOR2X1_LVT bpu_U82 ( .A1(ibuf_io_pc[22]), .A2(bpu_n76), .Y(bpu_n35) );
  XOR2X1_LVT bpu_U81 ( .A1(ibuf_io_pc[24]), .A2(bpu_n139), .Y(bpu_n34) );
  XOR2X1_LVT bpu_U80 ( .A1(ibuf_io_pc[17]), .A2(bpu_n141), .Y(bpu_n33) );
  XOR2X1_LVT bpu_U79 ( .A1(ibuf_io_pc[21]), .A2(bpu_n138), .Y(bpu_n32) );
  XOR2X1_LVT bpu_U78 ( .A1(ibuf_io_pc[11]), .A2(bpu_n142), .Y(bpu_n39) );
  XOR2X1_LVT bpu_U77 ( .A1(ibuf_io_pc[6]), .A2(bpu_n148), .Y(bpu_n38) );
  XOR2X1_LVT bpu_U76 ( .A1(ibuf_io_pc[10]), .A2(bpu_n90), .Y(bpu_n37) );
  XOR2X1_LVT bpu_U75 ( .A1(ibuf_io_pc[36]), .A2(bpu_n87), .Y(bpu_n36) );
  XOR2X1_LVT bpu_U74 ( .A1(ibuf_io_pc[12]), .A2(bpu_n117), .Y(bpu_n47) );
  XOR2X1_LVT bpu_U73 ( .A1(ibuf_io_pc[14]), .A2(bpu_n144), .Y(bpu_n46) );
  XOR2X1_LVT bpu_U72 ( .A1(ibuf_io_pc[4]), .A2(bpu_n119), .Y(bpu_n45) );
  XOR2X1_LVT bpu_U71 ( .A1(ibuf_io_pc[2]), .A2(bpu_n135), .Y(bpu_n50) );
  XOR2X1_LVT bpu_U70 ( .A1(ibuf_io_pc[37]), .A2(bpu_n123), .Y(bpu_n54) );
  XOR2X1_LVT bpu_U69 ( .A1(ibuf_io_pc[5]), .A2(bpu_n120), .Y(bpu_n53) );
  XOR2X1_LVT bpu_U68 ( .A1(ibuf_io_pc[33]), .A2(bpu_n73), .Y(bpu_n52) );
  XOR2X1_LVT bpu_U67 ( .A1(ibuf_io_pc[34]), .A2(bpu_n104), .Y(bpu_n51) );
  NOR4X1_LVT bpu_U66 ( .A1(bpu_n160), .A2(bpu_n159), .A3(bpu_n156), .A4(
        bpu_n155), .Y(bpu_n164) );
  XOR2X1_LVT bpu_U65 ( .A1(ibuf_io_pc[38]), .A2(bpu_n106), .Y(bpu_n11) );
  XOR2X1_LVT bpu_U64 ( .A1(ibuf_io_pc[29]), .A2(bpu_n126), .Y(bpu_n20) );
  XOR2X1_LVT bpu_U63 ( .A1(ibuf_io_pc[27]), .A2(bpu_n122), .Y(bpu_n18) );
  XOR2X1_LVT bpu_U62 ( .A1(ibuf_io_pc[31]), .A2(bpu_n101), .Y(bpu_n27) );
  XOR2X1_LVT bpu_U61 ( .A1(ibuf_io_pc[7]), .A2(bpu_n147), .Y(bpu_n30) );
  XOR2X1_LVT bpu_U60 ( .A1(ibuf_io_pc[3]), .A2(bpu_n79), .Y(bpu_n44) );
  XOR2X1_LVT bpu_U59 ( .A1(ibuf_io_pc[0]), .A2(bpu_n131), .Y(bpu_n49) );
  XOR2X1_LVT bpu_U58 ( .A1(ibuf_io_pc[1]), .A2(csr_io_bp_0_address[1]), .Y(
        bpu_n23) );
  XOR2X1_LVT bpu_U57 ( .A1(ibuf_io_pc[35]), .A2(bpu_n88), .Y(bpu_n10) );
  XOR2X1_LVT bpu_U56 ( .A1(ibuf_io_pc[18]), .A2(bpu_n94), .Y(bpu_n9) );
  XOR2X1_LVT bpu_U55 ( .A1(ibuf_io_pc[23]), .A2(bpu_n84), .Y(bpu_n8) );
  XOR2X1_LVT bpu_U54 ( .A1(ibuf_io_pc[13]), .A2(bpu_n93), .Y(bpu_n15) );
  XOR2X1_LVT bpu_U53 ( .A1(ibuf_io_pc[15]), .A2(bpu_n116), .Y(bpu_n14) );
  XOR2X1_LVT bpu_U52 ( .A1(ibuf_io_pc[9]), .A2(bpu_n85), .Y(bpu_n13) );
  XOR2X1_LVT bpu_U51 ( .A1(ibuf_io_pc[28]), .A2(bpu_n125), .Y(bpu_n12) );
  XOR2X1_LVT bpu_U50 ( .A1(ibuf_io_pc[20]), .A2(bpu_n109), .Y(bpu_n17) );
  INVX0_LVT bpu_U49 ( .A(bpu_n68), .Y(bpu_n154) );
  INVX0_LVT bpu_U48 ( .A(bpu_n_T_9), .Y(bpu_n161) );
  XOR2X1_LVT bpu_U47 ( .A1(bpu_n_T_73), .A2(csr_io_bp_0_control_tmatch[0]), 
        .Y(bpu_n63) );
  INVX1_LVT bpu_U46 ( .A(n_T_918[2]), .Y(bpu_n136) );
  INVX1_LVT bpu_U45 ( .A(n_T_918[3]), .Y(bpu_n78) );
  INVX1_LVT bpu_U44 ( .A(n_T_918[0]), .Y(bpu_n74) );
  INVX1_LVT bpu_U43 ( .A(n_T_918[22]), .Y(bpu_n77) );
  INVX1_LVT bpu_U42 ( .A(n_T_918[1]), .Y(bpu_n132) );
  INVX1_LVT bpu_U41 ( .A(csr_io_bp_0_control_tmatch[1]), .Y(bpu_n163) );
  INVX1_LVT bpu_U40 ( .A(csr_io_bp_0_control_tmatch[0]), .Y(bpu_n70) );
  INVX1_LVT bpu_U39 ( .A(csr_io_bp_0_address[23]), .Y(bpu_n84) );
  INVX1_LVT bpu_U38 ( .A(csr_io_bp_0_address[36]), .Y(bpu_n87) );
  INVX1_LVT bpu_U37 ( .A(csr_io_bp_0_address[35]), .Y(bpu_n88) );
  INVX1_LVT bpu_U36 ( .A(csr_io_bp_0_address[25]), .Y(bpu_n91) );
  INVX1_LVT bpu_U35 ( .A(csr_io_bp_0_address[10]), .Y(bpu_n90) );
  INVX1_LVT bpu_U34 ( .A(csr_io_bp_0_address[31]), .Y(bpu_n101) );
  INVX1_LVT bpu_U33 ( .A(csr_io_bp_0_address[30]), .Y(bpu_n100) );
  INVX1_LVT bpu_U32 ( .A(csr_io_bp_0_address[34]), .Y(bpu_n104) );
  INVX1_LVT bpu_U31 ( .A(csr_io_bp_0_address[32]), .Y(bpu_n103) );
  INVX1_LVT bpu_U30 ( .A(csr_io_bp_0_address[19]), .Y(bpu_n107) );
  INVX1_LVT bpu_U29 ( .A(csr_io_bp_0_address[38]), .Y(bpu_n106) );
  INVX0_LVT bpu_U28 ( .A(csr_io_bp_0_address[20]), .Y(bpu_n109) );
  INVX1_LVT bpu_U27 ( .A(csr_io_bp_0_address[16]), .Y(bpu_n110) );
  INVX1_LVT bpu_U26 ( .A(csr_io_bp_0_address[21]), .Y(bpu_n138) );
  INVX1_LVT bpu_U25 ( .A(csr_io_bp_0_address[24]), .Y(bpu_n139) );
  INVX1_LVT bpu_U24 ( .A(csr_io_bp_0_address[3]), .Y(bpu_n79) );
  INVX1_LVT bpu_U23 ( .A(csr_io_bp_0_address[33]), .Y(bpu_n73) );
  INVX1_LVT bpu_U22 ( .A(csr_io_bp_0_address[26]), .Y(bpu_n72) );
  INVX1_LVT bpu_U21 ( .A(csr_io_bp_0_address[22]), .Y(bpu_n76) );
  INVX1_LVT bpu_U20 ( .A(csr_io_bp_0_address[11]), .Y(bpu_n142) );
  INVX1_LVT bpu_U19 ( .A(csr_io_bp_0_address[17]), .Y(bpu_n141) );
  INVX1_LVT bpu_U18 ( .A(csr_io_bp_0_address[14]), .Y(bpu_n144) );
  INVX1_LVT bpu_U17 ( .A(csr_io_bp_0_address[8]), .Y(bpu_n145) );
  INVX1_LVT bpu_U16 ( .A(csr_io_bp_0_address[6]), .Y(bpu_n148) );
  INVX1_LVT bpu_U15 ( .A(csr_io_bp_0_address[12]), .Y(bpu_n117) );
  INVX1_LVT bpu_U14 ( .A(csr_io_bp_0_address[5]), .Y(bpu_n120) );
  INVX1_LVT bpu_U13 ( .A(csr_io_bp_0_address[4]), .Y(bpu_n119) );
  INVX1_LVT bpu_U12 ( .A(csr_io_bp_0_address[37]), .Y(bpu_n123) );
  INVX1_LVT bpu_U11 ( .A(csr_io_bp_0_address[27]), .Y(bpu_n122) );
  INVX1_LVT bpu_U10 ( .A(csr_io_bp_0_address[2]), .Y(bpu_n135) );
  INVX1_LVT bpu_U9 ( .A(csr_io_bp_0_address[1]), .Y(bpu_n133) );
  INVX1_LVT bpu_U8 ( .A(csr_io_bp_0_address[29]), .Y(bpu_n126) );
  INVX0_LVT bpu_U7 ( .A(csr_io_bp_0_address[28]), .Y(bpu_n125) );
  OA221X1_LVT bpu_U6 ( .A1(io_ptw_status_prv[0]), .A2(bpu_n2), .A3(bpu_n3), 
        .A4(bpu_n4), .A5(n9516), .Y(bpu_n67) );
  AO22X1_LVT bpu_U5 ( .A1(io_ptw_status_prv[1]), .A2(csr_io_bp_0_control_m), 
        .A3(bpu_n1), .A4(csr_io_bp_0_control_s), .Y(bpu_n4) );
  INVX0_LVT bpu_U4 ( .A(io_ptw_status_prv[0]), .Y(bpu_n3) );
  AND2X1_LVT bpu_U3 ( .A1(csr_io_bp_0_control_u), .A2(bpu_n1), .Y(bpu_n2) );
  INVX0_LVT bpu_U2 ( .A(io_ptw_status_prv[1]), .Y(bpu_n1) );
  AO22X1_LVT bpu_gte_x_5_U340 ( .A1(bpu_gte_x_5_n343), .A2(
        csr_io_bp_0_address[36]), .A3(bpu_gte_x_5_n344), .A4(
        csr_io_bp_0_address[35]), .Y(bpu_gte_x_5_n417) );
  AO221X1_LVT bpu_gte_x_5_U339 ( .A1(bpu_gte_x_5_n421), .A2(bpu_gte_x_5_n416), 
        .A3(bpu_gte_x_5_n421), .A4(bpu_gte_x_5_n422), .A5(bpu_gte_x_5_n417), 
        .Y(bpu_gte_x_5_n418) );
  OR2X1_LVT bpu_gte_x_5_U338 ( .A1(bpu_gte_x_5_n344), .A2(
        csr_io_bp_0_address[35]), .Y(bpu_gte_x_5_n420) );
  AO222X1_LVT bpu_gte_x_5_U337 ( .A1(csr_io_bp_0_address[36]), .A2(
        bpu_gte_x_5_n420), .A3(bpu_gte_x_5_n343), .A4(bpu_gte_x_5_n420), .A5(
        csr_io_bp_0_address[36]), .A6(bpu_gte_x_5_n343), .Y(bpu_gte_x_5_n419)
         );
  OA22X1_LVT bpu_gte_x_5_U336 ( .A1(ibuf_io_pc[37]), .A2(bpu_gte_x_5_n335), 
        .A3(ibuf_io_pc[38]), .A4(bpu_gte_x_5_n337), .Y(bpu_gte_x_5_n364) );
  AOI22X1_LVT bpu_gte_x_5_U335 ( .A1(csr_io_bp_0_address[32]), .A2(
        bpu_gte_x_5_n346), .A3(csr_io_bp_0_address[31]), .A4(bpu_gte_x_5_n347), 
        .Y(bpu_gte_x_5_n415) );
  AND4X1_LVT bpu_gte_x_5_U334 ( .A1(bpu_gte_x_5_n338), .A2(bpu_gte_x_5_n339), 
        .A3(bpu_gte_x_5_n364), .A4(bpu_gte_x_5_n415), .Y(bpu_gte_x_5_n365) );
  NAND2X0_LVT bpu_gte_x_5_U333 ( .A1(csr_io_bp_0_address[20]), .A2(
        bpu_gte_x_5_n354), .Y(bpu_gte_x_5_n413) );
  NAND2X0_LVT bpu_gte_x_5_U332 ( .A1(ibuf_io_pc[19]), .A2(bpu_gte_x_5_n413), 
        .Y(bpu_gte_x_5_n414) );
  OA22X1_LVT bpu_gte_x_5_U331 ( .A1(bpu_gte_x_5_n354), .A2(
        csr_io_bp_0_address[20]), .A3(bpu_gte_x_5_n414), .A4(
        csr_io_bp_0_address[19]), .Y(bpu_gte_x_5_n407) );
  NAND2X0_LVT bpu_gte_x_5_U330 ( .A1(csr_io_bp_0_address[16]), .A2(
        bpu_gte_x_5_n356), .Y(bpu_gte_x_5_n390) );
  AO22X1_LVT bpu_gte_x_5_U329 ( .A1(bpu_gte_x_5_n411), .A2(bpu_gte_x_5_n412), 
        .A3(bpu_gte_x_5_n411), .A4(bpu_gte_x_5_n387), .Y(bpu_gte_x_5_n408) );
  OA22X1_LVT bpu_gte_x_5_U328 ( .A1(bpu_gte_x_5_n353), .A2(
        csr_io_bp_0_address[22]), .A3(bpu_gte_x_5_n410), .A4(
        csr_io_bp_0_address[21]), .Y(bpu_gte_x_5_n409) );
  NAND2X0_LVT bpu_gte_x_5_U327 ( .A1(csr_io_bp_0_address[28]), .A2(
        bpu_gte_x_5_n349), .Y(bpu_gte_x_5_n382) );
  NAND2X0_LVT bpu_gte_x_5_U326 ( .A1(csr_io_bp_0_address[23]), .A2(
        bpu_gte_x_5_n352), .Y(bpu_gte_x_5_n405) );
  NAND2X0_LVT bpu_gte_x_5_U325 ( .A1(csr_io_bp_0_address[24]), .A2(
        bpu_gte_x_5_n351), .Y(bpu_gte_x_5_n379) );
  NAND4X0_LVT bpu_gte_x_5_U324 ( .A1(bpu_gte_x_5_n380), .A2(bpu_gte_x_5_n340), 
        .A3(bpu_gte_x_5_n405), .A4(bpu_gte_x_5_n379), .Y(bpu_gte_x_5_n368) );
  NAND2X0_LVT bpu_gte_x_5_U323 ( .A1(csr_io_bp_0_address[12]), .A2(
        bpu_gte_x_5_n358), .Y(bpu_gte_x_5_n404) );
  NAND2X0_LVT bpu_gte_x_5_U322 ( .A1(csr_io_bp_0_address[8]), .A2(
        bpu_gte_x_5_n360), .Y(bpu_gte_x_5_n399) );
  OR3X1_LVT bpu_gte_x_5_U321 ( .A1(bpu_gte_x_5_n396), .A2(bpu_gte_x_5_n397), 
        .A3(bpu_gte_x_5_n398), .Y(bpu_gte_x_5_n384) );
  NAND2X0_LVT bpu_gte_x_5_U320 ( .A1(csr_io_bp_0_address[4]), .A2(
        bpu_gte_x_5_n362), .Y(bpu_gte_x_5_n395) );
  OA221X1_LVT bpu_gte_x_5_U319 ( .A1(bpu_gte_x_5_n391), .A2(bpu_gte_x_5_n392), 
        .A3(bpu_gte_x_5_n393), .A4(bpu_gte_x_5_n392), .A5(bpu_gte_x_5_n394), 
        .Y(bpu_gte_x_5_n385) );
  OR3X1_LVT bpu_gte_x_5_U318 ( .A1(bpu_gte_x_5_n387), .A2(bpu_gte_x_5_n388), 
        .A3(bpu_gte_x_5_n389), .Y(bpu_gte_x_5_n386) );
  AO221X1_LVT bpu_gte_x_5_U317 ( .A1(bpu_gte_x_5_n383), .A2(bpu_gte_x_5_n384), 
        .A3(bpu_gte_x_5_n383), .A4(bpu_gte_x_5_n385), .A5(bpu_gte_x_5_n386), 
        .Y(bpu_gte_x_5_n369) );
  NAND2X0_LVT bpu_gte_x_5_U316 ( .A1(ibuf_io_pc[27]), .A2(bpu_gte_x_5_n382), 
        .Y(bpu_gte_x_5_n381) );
  OA22X1_LVT bpu_gte_x_5_U315 ( .A1(bpu_gte_x_5_n349), .A2(
        csr_io_bp_0_address[28]), .A3(bpu_gte_x_5_n381), .A4(
        csr_io_bp_0_address[27]), .Y(bpu_gte_x_5_n372) );
  AO22X1_LVT bpu_gte_x_5_U314 ( .A1(bpu_gte_x_5_n376), .A2(bpu_gte_x_5_n377), 
        .A3(bpu_gte_x_5_n376), .A4(bpu_gte_x_5_n378), .Y(bpu_gte_x_5_n373) );
  OA22X1_LVT bpu_gte_x_5_U313 ( .A1(bpu_gte_x_5_n348), .A2(
        csr_io_bp_0_address[30]), .A3(bpu_gte_x_5_n375), .A4(
        csr_io_bp_0_address[29]), .Y(bpu_gte_x_5_n374) );
  OAI221X1_LVT bpu_gte_x_5_U312 ( .A1(bpu_gte_x_5_n367), .A2(bpu_gte_x_5_n368), 
        .A3(bpu_gte_x_5_n369), .A4(bpu_gte_x_5_n368), .A5(bpu_gte_x_5_n370), 
        .Y(bpu_gte_x_5_n366) );
  AO222X1_LVT bpu_gte_x_5_U311 ( .A1(bpu_gte_x_5_n363), .A2(bpu_gte_x_5_n364), 
        .A3(bpu_gte_x_5_n337), .A4(ibuf_io_pc[38]), .A5(bpu_gte_x_5_n365), 
        .A6(bpu_gte_x_5_n366), .Y(bpu_n_T_73) );
  INVX1_LVT bpu_gte_x_5_U310 ( .A(bpu_gte_x_5_n378), .Y(bpu_gte_x_5_n340) );
  INVX1_LVT bpu_gte_x_5_U309 ( .A(bpu_gte_x_5_n417), .Y(bpu_gte_x_5_n338) );
  INVX1_LVT bpu_gte_x_5_U308 ( .A(csr_io_bp_0_address[38]), .Y(
        bpu_gte_x_5_n337) );
  NAND2X0_LVT bpu_gte_x_5_U307 ( .A1(bpu_gte_x_5_n335), .A2(ibuf_io_pc[37]), 
        .Y(bpu_gte_x_5_n334) );
  INVX1_LVT bpu_gte_x_5_U306 ( .A(csr_io_bp_0_address[37]), .Y(
        bpu_gte_x_5_n335) );
  AND2X1_LVT bpu_gte_x_5_U305 ( .A1(bpu_gte_x_5_n419), .A2(bpu_gte_x_5_n418), 
        .Y(bpu_gte_x_5_n333) );
  NAND2X0_LVT bpu_gte_x_5_U304 ( .A1(bpu_gte_x_5_n333), .A2(bpu_gte_x_5_n334), 
        .Y(bpu_gte_x_5_n363) );
  OA221X1_LVT bpu_gte_x_5_U303 ( .A1(bpu_gte_x_5_n408), .A2(bpu_gte_x_5_n388), 
        .A3(bpu_gte_x_5_n407), .A4(bpu_gte_x_5_n406), .A5(bpu_gte_x_5_n409), 
        .Y(bpu_gte_x_5_n367) );
  OA221X1_LVT bpu_gte_x_5_U302 ( .A1(bpu_gte_x_5_n402), .A2(bpu_gte_x_5_n397), 
        .A3(bpu_gte_x_5_n401), .A4(bpu_gte_x_5_n400), .A5(bpu_gte_x_5_n403), 
        .Y(bpu_gte_x_5_n383) );
  OA221X1_LVT bpu_gte_x_5_U301 ( .A1(bpu_gte_x_5_n373), .A2(bpu_gte_x_5_n336), 
        .A3(bpu_gte_x_5_n372), .A4(bpu_gte_x_5_n371), .A5(bpu_gte_x_5_n374), 
        .Y(bpu_gte_x_5_n370) );
  OAI21X1_LVT bpu_gte_x_5_U300 ( .A1(ibuf_io_pc[7]), .A2(bpu_gte_x_5_n342), 
        .A3(bpu_gte_x_5_n399), .Y(bpu_gte_x_5_n398) );
  OAI21X1_LVT bpu_gte_x_5_U299 ( .A1(ibuf_io_pc[15]), .A2(bpu_gte_x_5_n341), 
        .A3(bpu_gte_x_5_n390), .Y(bpu_gte_x_5_n389) );
  INVX0_LVT bpu_gte_x_5_U298 ( .A(bpu_gte_x_5_n416), .Y(bpu_gte_x_5_n339) );
  INVX0_LVT bpu_gte_x_5_U297 ( .A(bpu_gte_x_5_n380), .Y(bpu_gte_x_5_n336) );
  INVX1_LVT bpu_gte_x_5_U296 ( .A(ibuf_io_pc[30]), .Y(bpu_gte_x_5_n348) );
  INVX1_LVT bpu_gte_x_5_U295 ( .A(ibuf_io_pc[28]), .Y(bpu_gte_x_5_n349) );
  INVX1_LVT bpu_gte_x_5_U294 ( .A(ibuf_io_pc[26]), .Y(bpu_gte_x_5_n350) );
  INVX1_LVT bpu_gte_x_5_U293 ( .A(ibuf_io_pc[20]), .Y(bpu_gte_x_5_n354) );
  INVX1_LVT bpu_gte_x_5_U292 ( .A(ibuf_io_pc[22]), .Y(bpu_gte_x_5_n353) );
  INVX1_LVT bpu_gte_x_5_U291 ( .A(ibuf_io_pc[18]), .Y(bpu_gte_x_5_n355) );
  INVX1_LVT bpu_gte_x_5_U290 ( .A(ibuf_io_pc[6]), .Y(bpu_gte_x_5_n361) );
  INVX1_LVT bpu_gte_x_5_U289 ( .A(ibuf_io_pc[24]), .Y(bpu_gte_x_5_n351) );
  INVX1_LVT bpu_gte_x_5_U288 ( .A(ibuf_io_pc[23]), .Y(bpu_gte_x_5_n352) );
  INVX1_LVT bpu_gte_x_5_U287 ( .A(ibuf_io_pc[16]), .Y(bpu_gte_x_5_n356) );
  INVX1_LVT bpu_gte_x_5_U286 ( .A(csr_io_bp_0_address[15]), .Y(
        bpu_gte_x_5_n341) );
  INVX1_LVT bpu_gte_x_5_U285 ( .A(csr_io_bp_0_address[7]), .Y(bpu_gte_x_5_n342) );
  INVX1_LVT bpu_gte_x_5_U284 ( .A(ibuf_io_pc[8]), .Y(bpu_gte_x_5_n360) );
  INVX1_LVT bpu_gte_x_5_U283 ( .A(ibuf_io_pc[35]), .Y(bpu_gte_x_5_n344) );
  INVX1_LVT bpu_gte_x_5_U282 ( .A(ibuf_io_pc[10]), .Y(bpu_gte_x_5_n359) );
  INVX1_LVT bpu_gte_x_5_U281 ( .A(ibuf_io_pc[36]), .Y(bpu_gte_x_5_n343) );
  INVX1_LVT bpu_gte_x_5_U280 ( .A(ibuf_io_pc[12]), .Y(bpu_gte_x_5_n358) );
  INVX1_LVT bpu_gte_x_5_U279 ( .A(ibuf_io_pc[31]), .Y(bpu_gte_x_5_n347) );
  INVX1_LVT bpu_gte_x_5_U278 ( .A(ibuf_io_pc[32]), .Y(bpu_gte_x_5_n346) );
  INVX1_LVT bpu_gte_x_5_U277 ( .A(ibuf_io_pc[34]), .Y(bpu_gte_x_5_n345) );
  INVX1_LVT bpu_gte_x_5_U276 ( .A(ibuf_io_pc[4]), .Y(bpu_gte_x_5_n362) );
  INVX1_LVT bpu_gte_x_5_U275 ( .A(ibuf_io_pc[14]), .Y(bpu_gte_x_5_n357) );
  INVX0_LVT bpu_gte_x_5_U273 ( .A(bpu_gte_x_5_n404), .Y(bpu_gte_x_5_n331) );
  INVX0_LVT bpu_gte_x_5_U272 ( .A(ibuf_io_pc[11]), .Y(bpu_gte_x_5_n330) );
  AO22X1_LVT bpu_gte_x_5_U271 ( .A1(bpu_gte_x_5_n361), .A2(
        csr_io_bp_0_address[6]), .A3(csr_io_bp_0_address[5]), .A4(
        bpu_gte_x_5_n329), .Y(bpu_gte_x_5_n392) );
  INVX0_LVT bpu_gte_x_5_U270 ( .A(ibuf_io_pc[5]), .Y(bpu_gte_x_5_n329) );
  NAND2X0_LVT bpu_gte_x_5_U269 ( .A1(ibuf_io_pc[21]), .A2(bpu_gte_x_5_n328), 
        .Y(bpu_gte_x_5_n410) );
  NAND2X0_LVT bpu_gte_x_5_U268 ( .A1(bpu_gte_x_5_n353), .A2(
        csr_io_bp_0_address[22]), .Y(bpu_gte_x_5_n328) );
  NAND2X0_LVT bpu_gte_x_5_U267 ( .A1(ibuf_io_pc[29]), .A2(bpu_gte_x_5_n327), 
        .Y(bpu_gte_x_5_n375) );
  NAND2X0_LVT bpu_gte_x_5_U266 ( .A1(bpu_gte_x_5_n348), .A2(
        csr_io_bp_0_address[30]), .Y(bpu_gte_x_5_n327) );
  OA22X1_LVT bpu_gte_x_5_U265 ( .A1(csr_io_bp_0_address[24]), .A2(
        bpu_gte_x_5_n351), .A3(csr_io_bp_0_address[23]), .A4(bpu_gte_x_5_n326), 
        .Y(bpu_gte_x_5_n377) );
  NAND2X0_LVT bpu_gte_x_5_U264 ( .A1(bpu_gte_x_5_n379), .A2(ibuf_io_pc[23]), 
        .Y(bpu_gte_x_5_n326) );
  AO22X1_LVT bpu_gte_x_5_U263 ( .A1(bpu_gte_x_5_n359), .A2(
        csr_io_bp_0_address[10]), .A3(csr_io_bp_0_address[9]), .A4(
        bpu_gte_x_5_n325), .Y(bpu_gte_x_5_n396) );
  INVX0_LVT bpu_gte_x_5_U262 ( .A(ibuf_io_pc[9]), .Y(bpu_gte_x_5_n325) );
  OA22X1_LVT bpu_gte_x_5_U261 ( .A1(bpu_gte_x_5_n357), .A2(
        csr_io_bp_0_address[14]), .A3(csr_io_bp_0_address[13]), .A4(
        bpu_gte_x_5_n324), .Y(bpu_gte_x_5_n403) );
  NAND2X0_LVT bpu_gte_x_5_U260 ( .A1(ibuf_io_pc[13]), .A2(bpu_gte_x_5_n323), 
        .Y(bpu_gte_x_5_n324) );
  NAND2X0_LVT bpu_gte_x_5_U259 ( .A1(bpu_gte_x_5_n357), .A2(
        csr_io_bp_0_address[14]), .Y(bpu_gte_x_5_n323) );
  OA22X1_LVT bpu_gte_x_5_U258 ( .A1(csr_io_bp_0_address[16]), .A2(
        bpu_gte_x_5_n356), .A3(csr_io_bp_0_address[15]), .A4(bpu_gte_x_5_n322), 
        .Y(bpu_gte_x_5_n412) );
  NAND2X0_LVT bpu_gte_x_5_U257 ( .A1(bpu_gte_x_5_n390), .A2(ibuf_io_pc[15]), 
        .Y(bpu_gte_x_5_n322) );
  INVX0_LVT bpu_gte_x_5_U256 ( .A(bpu_gte_x_5_n413), .Y(bpu_gte_x_5_n321) );
  INVX0_LVT bpu_gte_x_5_U255 ( .A(ibuf_io_pc[19]), .Y(bpu_gte_x_5_n320) );
  OA22X1_LVT bpu_gte_x_5_U253 ( .A1(csr_io_bp_0_address[4]), .A2(
        bpu_gte_x_5_n362), .A3(csr_io_bp_0_address[3]), .A4(bpu_gte_x_5_n318), 
        .Y(bpu_gte_x_5_n393) );
  NAND2X0_LVT bpu_gte_x_5_U252 ( .A1(bpu_gte_x_5_n395), .A2(ibuf_io_pc[3]), 
        .Y(bpu_gte_x_5_n318) );
  AO22X1_LVT bpu_gte_x_5_U251 ( .A1(csr_io_bp_0_address[33]), .A2(
        bpu_gte_x_5_n317), .A3(csr_io_bp_0_address[34]), .A4(bpu_gte_x_5_n345), 
        .Y(bpu_gte_x_5_n416) );
  INVX0_LVT bpu_gte_x_5_U250 ( .A(ibuf_io_pc[33]), .Y(bpu_gte_x_5_n317) );
  OA22X1_LVT bpu_gte_x_5_U249 ( .A1(bpu_gte_x_5_n346), .A2(
        csr_io_bp_0_address[32]), .A3(csr_io_bp_0_address[31]), .A4(
        bpu_gte_x_5_n316), .Y(bpu_gte_x_5_n422) );
  NAND2X0_LVT bpu_gte_x_5_U248 ( .A1(ibuf_io_pc[31]), .A2(bpu_gte_x_5_n315), 
        .Y(bpu_gte_x_5_n316) );
  NAND2X0_LVT bpu_gte_x_5_U247 ( .A1(bpu_gte_x_5_n346), .A2(
        csr_io_bp_0_address[32]), .Y(bpu_gte_x_5_n315) );
  OA22X1_LVT bpu_gte_x_5_U246 ( .A1(csr_io_bp_0_address[12]), .A2(
        bpu_gte_x_5_n358), .A3(csr_io_bp_0_address[11]), .A4(bpu_gte_x_5_n314), 
        .Y(bpu_gte_x_5_n401) );
  NAND2X0_LVT bpu_gte_x_5_U245 ( .A1(bpu_gte_x_5_n404), .A2(ibuf_io_pc[11]), 
        .Y(bpu_gte_x_5_n314) );
  AO22X1_LVT bpu_gte_x_5_U244 ( .A1(bpu_gte_x_5_n357), .A2(
        csr_io_bp_0_address[14]), .A3(csr_io_bp_0_address[13]), .A4(
        bpu_gte_x_5_n313), .Y(bpu_gte_x_5_n400) );
  INVX0_LVT bpu_gte_x_5_U243 ( .A(ibuf_io_pc[13]), .Y(bpu_gte_x_5_n313) );
  OA222X1_LVT bpu_gte_x_5_U242 ( .A1(bpu_gte_x_5_n310), .A2(
        csr_io_bp_0_address[9]), .A3(bpu_gte_x_5_n359), .A4(
        csr_io_bp_0_address[10]), .A5(bpu_gte_x_5_n396), .A6(bpu_gte_x_5_n312), 
        .Y(bpu_gte_x_5_n402) );
  OA22X1_LVT bpu_gte_x_5_U241 ( .A1(csr_io_bp_0_address[8]), .A2(
        bpu_gte_x_5_n360), .A3(csr_io_bp_0_address[7]), .A4(bpu_gte_x_5_n311), 
        .Y(bpu_gte_x_5_n312) );
  NAND2X0_LVT bpu_gte_x_5_U240 ( .A1(bpu_gte_x_5_n399), .A2(ibuf_io_pc[7]), 
        .Y(bpu_gte_x_5_n311) );
  NAND2X0_LVT bpu_gte_x_5_U239 ( .A1(ibuf_io_pc[9]), .A2(bpu_gte_x_5_n309), 
        .Y(bpu_gte_x_5_n310) );
  NAND2X0_LVT bpu_gte_x_5_U238 ( .A1(bpu_gte_x_5_n359), .A2(
        csr_io_bp_0_address[10]), .Y(bpu_gte_x_5_n309) );
  AO22X1_LVT bpu_gte_x_5_U237 ( .A1(bpu_gte_x_5_n353), .A2(
        csr_io_bp_0_address[22]), .A3(csr_io_bp_0_address[21]), .A4(
        bpu_gte_x_5_n308), .Y(bpu_gte_x_5_n406) );
  INVX0_LVT bpu_gte_x_5_U236 ( .A(ibuf_io_pc[21]), .Y(bpu_gte_x_5_n308) );
  OA22X1_LVT bpu_gte_x_5_U235 ( .A1(bpu_gte_x_5_n345), .A2(
        csr_io_bp_0_address[34]), .A3(csr_io_bp_0_address[33]), .A4(
        bpu_gte_x_5_n307), .Y(bpu_gte_x_5_n421) );
  NAND2X0_LVT bpu_gte_x_5_U234 ( .A1(ibuf_io_pc[33]), .A2(bpu_gte_x_5_n306), 
        .Y(bpu_gte_x_5_n307) );
  NAND2X0_LVT bpu_gte_x_5_U233 ( .A1(bpu_gte_x_5_n345), .A2(
        csr_io_bp_0_address[34]), .Y(bpu_gte_x_5_n306) );
  OA22X1_LVT bpu_gte_x_5_U232 ( .A1(bpu_gte_x_5_n361), .A2(
        csr_io_bp_0_address[6]), .A3(csr_io_bp_0_address[5]), .A4(
        bpu_gte_x_5_n305), .Y(bpu_gte_x_5_n394) );
  NAND2X0_LVT bpu_gte_x_5_U231 ( .A1(ibuf_io_pc[5]), .A2(bpu_gte_x_5_n304), 
        .Y(bpu_gte_x_5_n305) );
  NAND2X0_LVT bpu_gte_x_5_U230 ( .A1(bpu_gte_x_5_n361), .A2(
        csr_io_bp_0_address[6]), .Y(bpu_gte_x_5_n304) );
  AO22X1_LVT bpu_gte_x_5_U229 ( .A1(bpu_gte_x_5_n355), .A2(
        csr_io_bp_0_address[18]), .A3(csr_io_bp_0_address[17]), .A4(
        bpu_gte_x_5_n303), .Y(bpu_gte_x_5_n387) );
  INVX0_LVT bpu_gte_x_5_U228 ( .A(ibuf_io_pc[17]), .Y(bpu_gte_x_5_n303) );
  AO22X1_LVT bpu_gte_x_5_U227 ( .A1(csr_io_bp_0_address[25]), .A2(
        bpu_gte_x_5_n302), .A3(csr_io_bp_0_address[26]), .A4(bpu_gte_x_5_n350), 
        .Y(bpu_gte_x_5_n378) );
  INVX0_LVT bpu_gte_x_5_U226 ( .A(ibuf_io_pc[25]), .Y(bpu_gte_x_5_n302) );
  OA22X1_LVT bpu_gte_x_5_U225 ( .A1(bpu_gte_x_5_n355), .A2(
        csr_io_bp_0_address[18]), .A3(csr_io_bp_0_address[17]), .A4(
        bpu_gte_x_5_n301), .Y(bpu_gte_x_5_n411) );
  NAND2X0_LVT bpu_gte_x_5_U224 ( .A1(ibuf_io_pc[17]), .A2(bpu_gte_x_5_n300), 
        .Y(bpu_gte_x_5_n301) );
  NAND2X0_LVT bpu_gte_x_5_U223 ( .A1(bpu_gte_x_5_n355), .A2(
        csr_io_bp_0_address[18]), .Y(bpu_gte_x_5_n300) );
  OA22X1_LVT bpu_gte_x_5_U222 ( .A1(bpu_gte_x_5_n350), .A2(
        csr_io_bp_0_address[26]), .A3(csr_io_bp_0_address[25]), .A4(
        bpu_gte_x_5_n299), .Y(bpu_gte_x_5_n376) );
  NAND2X0_LVT bpu_gte_x_5_U221 ( .A1(ibuf_io_pc[25]), .A2(bpu_gte_x_5_n298), 
        .Y(bpu_gte_x_5_n299) );
  NAND2X0_LVT bpu_gte_x_5_U220 ( .A1(bpu_gte_x_5_n350), .A2(
        csr_io_bp_0_address[26]), .Y(bpu_gte_x_5_n298) );
  INVX0_LVT bpu_gte_x_5_U218 ( .A(bpu_gte_x_5_n371), .Y(bpu_gte_x_5_n296) );
  INVX0_LVT bpu_gte_x_5_U217 ( .A(csr_io_bp_0_address[27]), .Y(
        bpu_gte_x_5_n295) );
  NAND3X0_LVT bpu_gte_x_5_U216 ( .A1(bpu_gte_x_5_n294), .A2(bpu_gte_x_5_n395), 
        .A3(bpu_gte_x_5_n293), .Y(bpu_gte_x_5_n391) );
  NAND2X0_LVT bpu_gte_x_5_U215 ( .A1(bpu_gte_x_5_n291), .A2(bpu_gte_x_5_n288), 
        .Y(bpu_gte_x_5_n294) );
  NAND2X0_LVT bpu_gte_x_5_U214 ( .A1(csr_io_bp_0_address[3]), .A2(
        bpu_gte_x_5_n292), .Y(bpu_gte_x_5_n293) );
  INVX0_LVT bpu_gte_x_5_U213 ( .A(ibuf_io_pc[3]), .Y(bpu_gte_x_5_n292) );
  OA22X1_LVT bpu_gte_x_5_U212 ( .A1(csr_io_bp_0_address[2]), .A2(
        bpu_gte_x_5_n286), .A3(csr_io_bp_0_address[1]), .A4(bpu_gte_x_5_n290), 
        .Y(bpu_gte_x_5_n291) );
  NAND2X0_LVT bpu_gte_x_5_U211 ( .A1(ibuf_io_pc[1]), .A2(bpu_gte_x_5_n289), 
        .Y(bpu_gte_x_5_n290) );
  NAND2X0_LVT bpu_gte_x_5_U210 ( .A1(csr_io_bp_0_address[2]), .A2(
        bpu_gte_x_5_n286), .Y(bpu_gte_x_5_n289) );
  AO222X1_LVT bpu_gte_x_5_U209 ( .A1(bpu_gte_x_5_n285), .A2(
        csr_io_bp_0_address[0]), .A3(bpu_gte_x_5_n286), .A4(
        csr_io_bp_0_address[2]), .A5(bpu_gte_x_5_n287), .A6(
        csr_io_bp_0_address[1]), .Y(bpu_gte_x_5_n288) );
  INVX0_LVT bpu_gte_x_5_U208 ( .A(ibuf_io_pc[1]), .Y(bpu_gte_x_5_n287) );
  INVX0_LVT bpu_gte_x_5_U207 ( .A(ibuf_io_pc[2]), .Y(bpu_gte_x_5_n286) );
  INVX0_LVT bpu_gte_x_5_U206 ( .A(ibuf_io_pc[0]), .Y(bpu_gte_x_5_n285) );
  AO22X1_LVT bpu_gte_x_5_U205 ( .A1(csr_io_bp_0_address[29]), .A2(
        bpu_gte_x_5_n284), .A3(csr_io_bp_0_address[30]), .A4(bpu_gte_x_5_n348), 
        .Y(bpu_gte_x_5_n371) );
  INVX0_LVT bpu_gte_x_5_U204 ( .A(ibuf_io_pc[29]), .Y(bpu_gte_x_5_n284) );
  OA221X1_LVT bpu_gte_x_5_U203 ( .A1(1'b0), .A2(bpu_gte_x_5_n382), .A3(
        ibuf_io_pc[27]), .A4(bpu_gte_x_5_n295), .A5(bpu_gte_x_5_n296), .Y(
        bpu_gte_x_5_n380) );
  AO221X1_LVT bpu_gte_x_5_U202 ( .A1(1'b1), .A2(bpu_gte_x_5_n406), .A3(
        csr_io_bp_0_address[19]), .A4(bpu_gte_x_5_n320), .A5(bpu_gte_x_5_n321), 
        .Y(bpu_gte_x_5_n388) );
  AO221X1_LVT bpu_gte_x_5_U201 ( .A1(1'b1), .A2(bpu_gte_x_5_n400), .A3(
        csr_io_bp_0_address[11]), .A4(bpu_gte_x_5_n330), .A5(bpu_gte_x_5_n331), 
        .Y(bpu_gte_x_5_n397) );
  NAND2X0_LVT bpu_gte_x_2_U341 ( .A1(csr_io_bp_0_address[34]), .A2(
        bpu_gte_x_2_n320), .Y(bpu_gte_x_2_n423) );
  NAND2X0_LVT bpu_gte_x_2_U340 ( .A1(n_T_918[33]), .A2(bpu_gte_x_2_n423), .Y(
        bpu_gte_x_2_n422) );
  OA22X1_LVT bpu_gte_x_2_U339 ( .A1(csr_io_bp_0_address[34]), .A2(
        bpu_gte_x_2_n320), .A3(csr_io_bp_0_address[33]), .A4(bpu_gte_x_2_n422), 
        .Y(bpu_gte_x_2_n418) );
  AO22X1_LVT bpu_gte_x_2_U338 ( .A1(bpu_gte_x_2_n321), .A2(
        csr_io_bp_0_address[33]), .A3(bpu_gte_x_2_n320), .A4(
        csr_io_bp_0_address[34]), .Y(bpu_gte_x_2_n413) );
  NAND2X0_LVT bpu_gte_x_2_U337 ( .A1(csr_io_bp_0_address[32]), .A2(
        bpu_gte_x_2_n322), .Y(bpu_gte_x_2_n421) );
  NAND2X0_LVT bpu_gte_x_2_U336 ( .A1(n_T_918[31]), .A2(bpu_gte_x_2_n421), .Y(
        bpu_gte_x_2_n420) );
  OA22X1_LVT bpu_gte_x_2_U335 ( .A1(bpu_gte_x_2_n420), .A2(
        csr_io_bp_0_address[31]), .A3(bpu_gte_x_2_n322), .A4(
        csr_io_bp_0_address[32]), .Y(bpu_gte_x_2_n419) );
  AO22X1_LVT bpu_gte_x_2_U334 ( .A1(bpu_gte_x_2_n318), .A2(
        csr_io_bp_0_address[36]), .A3(bpu_gte_x_2_n319), .A4(
        csr_io_bp_0_address[35]), .Y(bpu_gte_x_2_n414) );
  AO221X1_LVT bpu_gte_x_2_U333 ( .A1(bpu_gte_x_2_n418), .A2(bpu_gte_x_2_n413), 
        .A3(bpu_gte_x_2_n418), .A4(bpu_gte_x_2_n419), .A5(bpu_gte_x_2_n414), 
        .Y(bpu_gte_x_2_n415) );
  OR2X1_LVT bpu_gte_x_2_U332 ( .A1(bpu_gte_x_2_n319), .A2(
        csr_io_bp_0_address[35]), .Y(bpu_gte_x_2_n417) );
  AO222X1_LVT bpu_gte_x_2_U331 ( .A1(csr_io_bp_0_address[36]), .A2(
        bpu_gte_x_2_n417), .A3(bpu_gte_x_2_n318), .A4(bpu_gte_x_2_n417), .A5(
        csr_io_bp_0_address[36]), .A6(bpu_gte_x_2_n318), .Y(bpu_gte_x_2_n416)
         );
  OA22X1_LVT bpu_gte_x_2_U330 ( .A1(n_T_918[37]), .A2(bpu_gte_x_2_n309), .A3(
        n_T_918[38]), .A4(bpu_gte_x_2_n311), .Y(bpu_gte_x_2_n347) );
  AOI22X1_LVT bpu_gte_x_2_U329 ( .A1(csr_io_bp_0_address[32]), .A2(
        bpu_gte_x_2_n322), .A3(csr_io_bp_0_address[31]), .A4(bpu_gte_x_2_n323), 
        .Y(bpu_gte_x_2_n412) );
  AND4X1_LVT bpu_gte_x_2_U328 ( .A1(bpu_gte_x_2_n312), .A2(bpu_gte_x_2_n313), 
        .A3(bpu_gte_x_2_n347), .A4(bpu_gte_x_2_n412), .Y(bpu_gte_x_2_n348) );
  AO22X1_LVT bpu_gte_x_2_U327 ( .A1(csr_io_bp_0_address[21]), .A2(
        bpu_gte_x_2_n332), .A3(csr_io_bp_0_address[22]), .A4(bpu_gte_x_2_n331), 
        .Y(bpu_gte_x_2_n399) );
  NAND2X0_LVT bpu_gte_x_2_U326 ( .A1(csr_io_bp_0_address[20]), .A2(
        bpu_gte_x_2_n333), .Y(bpu_gte_x_2_n410) );
  NAND2X0_LVT bpu_gte_x_2_U325 ( .A1(n_T_918[19]), .A2(bpu_gte_x_2_n410), .Y(
        bpu_gte_x_2_n411) );
  OA22X1_LVT bpu_gte_x_2_U324 ( .A1(bpu_gte_x_2_n333), .A2(
        csr_io_bp_0_address[20]), .A3(bpu_gte_x_2_n411), .A4(
        csr_io_bp_0_address[19]), .Y(bpu_gte_x_2_n400) );
  NAND2X0_LVT bpu_gte_x_2_U323 ( .A1(csr_io_bp_0_address[18]), .A2(
        bpu_gte_x_2_n334), .Y(bpu_gte_x_2_n409) );
  NAND2X0_LVT bpu_gte_x_2_U322 ( .A1(n_T_918[17]), .A2(bpu_gte_x_2_n409), .Y(
        bpu_gte_x_2_n408) );
  OA22X1_LVT bpu_gte_x_2_U321 ( .A1(csr_io_bp_0_address[18]), .A2(
        bpu_gte_x_2_n334), .A3(csr_io_bp_0_address[17]), .A4(bpu_gte_x_2_n408), 
        .Y(bpu_gte_x_2_n405) );
  NAND2X0_LVT bpu_gte_x_2_U320 ( .A1(csr_io_bp_0_address[16]), .A2(
        bpu_gte_x_2_n336), .Y(bpu_gte_x_2_n377) );
  NAND2X0_LVT bpu_gte_x_2_U319 ( .A1(n_T_918[15]), .A2(bpu_gte_x_2_n377), .Y(
        bpu_gte_x_2_n407) );
  OA22X1_LVT bpu_gte_x_2_U318 ( .A1(bpu_gte_x_2_n336), .A2(
        csr_io_bp_0_address[16]), .A3(bpu_gte_x_2_n407), .A4(
        csr_io_bp_0_address[15]), .Y(bpu_gte_x_2_n406) );
  AO22X1_LVT bpu_gte_x_2_U317 ( .A1(csr_io_bp_0_address[17]), .A2(
        bpu_gte_x_2_n335), .A3(csr_io_bp_0_address[18]), .A4(bpu_gte_x_2_n334), 
        .Y(bpu_gte_x_2_n374) );
  AO22X1_LVT bpu_gte_x_2_U316 ( .A1(bpu_gte_x_2_n405), .A2(bpu_gte_x_2_n406), 
        .A3(bpu_gte_x_2_n405), .A4(bpu_gte_x_2_n374), .Y(bpu_gte_x_2_n401) );
  NAND2X0_LVT bpu_gte_x_2_U315 ( .A1(csr_io_bp_0_address[22]), .A2(
        bpu_gte_x_2_n331), .Y(bpu_gte_x_2_n404) );
  NAND2X0_LVT bpu_gte_x_2_U314 ( .A1(n_T_918[21]), .A2(bpu_gte_x_2_n404), .Y(
        bpu_gte_x_2_n403) );
  OA22X1_LVT bpu_gte_x_2_U313 ( .A1(bpu_gte_x_2_n331), .A2(
        csr_io_bp_0_address[22]), .A3(bpu_gte_x_2_n403), .A4(
        csr_io_bp_0_address[21]), .Y(bpu_gte_x_2_n402) );
  AO22X1_LVT bpu_gte_x_2_U312 ( .A1(bpu_gte_x_2_n325), .A2(
        csr_io_bp_0_address[29]), .A3(bpu_gte_x_2_n324), .A4(
        csr_io_bp_0_address[30]), .Y(bpu_gte_x_2_n354) );
  NAND2X0_LVT bpu_gte_x_2_U311 ( .A1(csr_io_bp_0_address[28]), .A2(
        bpu_gte_x_2_n326), .Y(bpu_gte_x_2_n369) );
  AO22X1_LVT bpu_gte_x_2_U310 ( .A1(bpu_gte_x_2_n328), .A2(
        csr_io_bp_0_address[25]), .A3(bpu_gte_x_2_n327), .A4(
        csr_io_bp_0_address[26]), .Y(bpu_gte_x_2_n362) );
  NAND2X0_LVT bpu_gte_x_2_U309 ( .A1(csr_io_bp_0_address[23]), .A2(
        bpu_gte_x_2_n330), .Y(bpu_gte_x_2_n398) );
  NAND2X0_LVT bpu_gte_x_2_U308 ( .A1(csr_io_bp_0_address[24]), .A2(
        bpu_gte_x_2_n329), .Y(bpu_gte_x_2_n364) );
  NAND4X0_LVT bpu_gte_x_2_U307 ( .A1(bpu_gte_x_2_n367), .A2(bpu_gte_x_2_n315), 
        .A3(bpu_gte_x_2_n398), .A4(bpu_gte_x_2_n364), .Y(bpu_gte_x_2_n351) );
  AO22X1_LVT bpu_gte_x_2_U306 ( .A1(csr_io_bp_0_address[13]), .A2(
        bpu_gte_x_2_n338), .A3(csr_io_bp_0_address[14]), .A4(bpu_gte_x_2_n337), 
        .Y(bpu_gte_x_2_n390) );
  NAND2X0_LVT bpu_gte_x_2_U305 ( .A1(csr_io_bp_0_address[12]), .A2(
        bpu_gte_x_2_n339), .Y(bpu_gte_x_2_n396) );
  NAND2X0_LVT bpu_gte_x_2_U304 ( .A1(n_T_918[11]), .A2(bpu_gte_x_2_n396), .Y(
        bpu_gte_x_2_n397) );
  OA22X1_LVT bpu_gte_x_2_U303 ( .A1(bpu_gte_x_2_n339), .A2(
        csr_io_bp_0_address[12]), .A3(bpu_gte_x_2_n397), .A4(
        csr_io_bp_0_address[11]), .Y(bpu_gte_x_2_n391) );
  NAND2X0_LVT bpu_gte_x_2_U302 ( .A1(csr_io_bp_0_address[8]), .A2(
        bpu_gte_x_2_n342), .Y(bpu_gte_x_2_n389) );
  AO22X1_LVT bpu_gte_x_2_U301 ( .A1(csr_io_bp_0_address[9]), .A2(
        bpu_gte_x_2_n341), .A3(csr_io_bp_0_address[10]), .A4(bpu_gte_x_2_n340), 
        .Y(bpu_gte_x_2_n386) );
  NAND2X0_LVT bpu_gte_x_2_U300 ( .A1(csr_io_bp_0_address[14]), .A2(
        bpu_gte_x_2_n337), .Y(bpu_gte_x_2_n395) );
  NAND2X0_LVT bpu_gte_x_2_U299 ( .A1(n_T_918[13]), .A2(bpu_gte_x_2_n395), .Y(
        bpu_gte_x_2_n394) );
  OA22X1_LVT bpu_gte_x_2_U298 ( .A1(bpu_gte_x_2_n337), .A2(
        csr_io_bp_0_address[14]), .A3(bpu_gte_x_2_n394), .A4(
        csr_io_bp_0_address[13]), .Y(bpu_gte_x_2_n393) );
  OAI21X1_LVT bpu_gte_x_2_U297 ( .A1(n_T_918[7]), .A2(bpu_gte_x_2_n317), .A3(
        bpu_gte_x_2_n389), .Y(bpu_gte_x_2_n388) );
  OR3X1_LVT bpu_gte_x_2_U296 ( .A1(bpu_gte_x_2_n386), .A2(bpu_gte_x_2_n387), 
        .A3(bpu_gte_x_2_n388), .Y(bpu_gte_x_2_n371) );
  NAND2X0_LVT bpu_gte_x_2_U295 ( .A1(csr_io_bp_0_address[4]), .A2(
        bpu_gte_x_2_n345), .Y(bpu_gte_x_2_n385) );
  AO22X1_LVT bpu_gte_x_2_U294 ( .A1(csr_io_bp_0_address[5]), .A2(
        bpu_gte_x_2_n344), .A3(csr_io_bp_0_address[6]), .A4(bpu_gte_x_2_n343), 
        .Y(bpu_gte_x_2_n379) );
  NAND2X0_LVT bpu_gte_x_2_U293 ( .A1(n_T_918[3]), .A2(bpu_gte_x_2_n385), .Y(
        bpu_gte_x_2_n384) );
  OA22X1_LVT bpu_gte_x_2_U292 ( .A1(bpu_gte_x_2_n384), .A2(
        csr_io_bp_0_address[3]), .A3(bpu_gte_x_2_n345), .A4(
        csr_io_bp_0_address[4]), .Y(bpu_gte_x_2_n380) );
  NAND2X0_LVT bpu_gte_x_2_U291 ( .A1(csr_io_bp_0_address[6]), .A2(
        bpu_gte_x_2_n343), .Y(bpu_gte_x_2_n383) );
  NAND2X0_LVT bpu_gte_x_2_U290 ( .A1(n_T_918[5]), .A2(bpu_gte_x_2_n383), .Y(
        bpu_gte_x_2_n382) );
  OA22X1_LVT bpu_gte_x_2_U289 ( .A1(bpu_gte_x_2_n343), .A2(
        csr_io_bp_0_address[6]), .A3(bpu_gte_x_2_n382), .A4(
        csr_io_bp_0_address[5]), .Y(bpu_gte_x_2_n381) );
  OA221X1_LVT bpu_gte_x_2_U288 ( .A1(bpu_gte_x_2_n378), .A2(bpu_gte_x_2_n379), 
        .A3(bpu_gte_x_2_n380), .A4(bpu_gte_x_2_n379), .A5(bpu_gte_x_2_n381), 
        .Y(bpu_gte_x_2_n372) );
  OAI21X1_LVT bpu_gte_x_2_U287 ( .A1(n_T_918[15]), .A2(bpu_gte_x_2_n316), .A3(
        bpu_gte_x_2_n377), .Y(bpu_gte_x_2_n376) );
  OR3X1_LVT bpu_gte_x_2_U286 ( .A1(bpu_gte_x_2_n374), .A2(bpu_gte_x_2_n375), 
        .A3(bpu_gte_x_2_n376), .Y(bpu_gte_x_2_n373) );
  AO221X1_LVT bpu_gte_x_2_U285 ( .A1(bpu_gte_x_2_n370), .A2(bpu_gte_x_2_n371), 
        .A3(bpu_gte_x_2_n370), .A4(bpu_gte_x_2_n372), .A5(bpu_gte_x_2_n373), 
        .Y(bpu_gte_x_2_n352) );
  NAND2X0_LVT bpu_gte_x_2_U284 ( .A1(n_T_918[27]), .A2(bpu_gte_x_2_n369), .Y(
        bpu_gte_x_2_n368) );
  OA22X1_LVT bpu_gte_x_2_U283 ( .A1(bpu_gte_x_2_n326), .A2(
        csr_io_bp_0_address[28]), .A3(bpu_gte_x_2_n368), .A4(
        csr_io_bp_0_address[27]), .Y(bpu_gte_x_2_n355) );
  NAND2X0_LVT bpu_gte_x_2_U282 ( .A1(csr_io_bp_0_address[26]), .A2(
        bpu_gte_x_2_n327), .Y(bpu_gte_x_2_n366) );
  NAND2X0_LVT bpu_gte_x_2_U281 ( .A1(n_T_918[25]), .A2(bpu_gte_x_2_n366), .Y(
        bpu_gte_x_2_n365) );
  OA22X1_LVT bpu_gte_x_2_U280 ( .A1(csr_io_bp_0_address[26]), .A2(
        bpu_gte_x_2_n327), .A3(csr_io_bp_0_address[25]), .A4(bpu_gte_x_2_n365), 
        .Y(bpu_gte_x_2_n360) );
  NAND2X0_LVT bpu_gte_x_2_U279 ( .A1(n_T_918[23]), .A2(bpu_gte_x_2_n364), .Y(
        bpu_gte_x_2_n363) );
  OA22X1_LVT bpu_gte_x_2_U278 ( .A1(bpu_gte_x_2_n329), .A2(
        csr_io_bp_0_address[24]), .A3(bpu_gte_x_2_n363), .A4(
        csr_io_bp_0_address[23]), .Y(bpu_gte_x_2_n361) );
  AO22X1_LVT bpu_gte_x_2_U277 ( .A1(bpu_gte_x_2_n360), .A2(bpu_gte_x_2_n361), 
        .A3(bpu_gte_x_2_n360), .A4(bpu_gte_x_2_n362), .Y(bpu_gte_x_2_n356) );
  NAND2X0_LVT bpu_gte_x_2_U276 ( .A1(csr_io_bp_0_address[30]), .A2(
        bpu_gte_x_2_n324), .Y(bpu_gte_x_2_n359) );
  NAND2X0_LVT bpu_gte_x_2_U275 ( .A1(n_T_918[29]), .A2(bpu_gte_x_2_n359), .Y(
        bpu_gte_x_2_n358) );
  OA22X1_LVT bpu_gte_x_2_U274 ( .A1(bpu_gte_x_2_n324), .A2(
        csr_io_bp_0_address[30]), .A3(bpu_gte_x_2_n358), .A4(
        csr_io_bp_0_address[29]), .Y(bpu_gte_x_2_n357) );
  OAI221X1_LVT bpu_gte_x_2_U273 ( .A1(bpu_gte_x_2_n350), .A2(bpu_gte_x_2_n351), 
        .A3(bpu_gte_x_2_n352), .A4(bpu_gte_x_2_n351), .A5(bpu_gte_x_2_n353), 
        .Y(bpu_gte_x_2_n349) );
  AO222X1_LVT bpu_gte_x_2_U272 ( .A1(bpu_gte_x_2_n346), .A2(bpu_gte_x_2_n347), 
        .A3(bpu_gte_x_2_n311), .A4(n_T_918[38]), .A5(bpu_gte_x_2_n348), .A6(
        bpu_gte_x_2_n349), .Y(bpu_n_T_9) );
  INVX1_LVT bpu_gte_x_2_U271 ( .A(bpu_gte_x_2_n362), .Y(bpu_gte_x_2_n315) );
  INVX1_LVT bpu_gte_x_2_U270 ( .A(bpu_gte_x_2_n413), .Y(bpu_gte_x_2_n313) );
  INVX1_LVT bpu_gte_x_2_U269 ( .A(bpu_gte_x_2_n414), .Y(bpu_gte_x_2_n312) );
  NAND2X0_LVT bpu_gte_x_2_U268 ( .A1(bpu_gte_x_2_n309), .A2(n_T_918[37]), .Y(
        bpu_gte_x_2_n308) );
  AND2X1_LVT bpu_gte_x_2_U267 ( .A1(bpu_gte_x_2_n416), .A2(bpu_gte_x_2_n415), 
        .Y(bpu_gte_x_2_n307) );
  NAND2X0_LVT bpu_gte_x_2_U266 ( .A1(bpu_gte_x_2_n307), .A2(bpu_gte_x_2_n308), 
        .Y(bpu_gte_x_2_n346) );
  OA221X1_LVT bpu_gte_x_2_U265 ( .A1(bpu_gte_x_2_n401), .A2(bpu_gte_x_2_n375), 
        .A3(bpu_gte_x_2_n400), .A4(bpu_gte_x_2_n399), .A5(bpu_gte_x_2_n402), 
        .Y(bpu_gte_x_2_n350) );
  NAND2X0_LVT bpu_gte_x_2_U264 ( .A1(bpu_gte_x_2_n306), .A2(
        csr_io_bp_0_address[27]), .Y(bpu_gte_x_2_n305) );
  AND2X1_LVT bpu_gte_x_2_U263 ( .A1(bpu_gte_x_2_n369), .A2(bpu_gte_x_2_n314), 
        .Y(bpu_gte_x_2_n304) );
  AND2X1_LVT bpu_gte_x_2_U262 ( .A1(bpu_gte_x_2_n304), .A2(bpu_gte_x_2_n305), 
        .Y(bpu_gte_x_2_n367) );
  OA221X1_LVT bpu_gte_x_2_U261 ( .A1(bpu_gte_x_2_n392), .A2(bpu_gte_x_2_n387), 
        .A3(bpu_gte_x_2_n391), .A4(bpu_gte_x_2_n390), .A5(bpu_gte_x_2_n393), 
        .Y(bpu_gte_x_2_n370) );
  OA221X1_LVT bpu_gte_x_2_U260 ( .A1(bpu_gte_x_2_n356), .A2(bpu_gte_x_2_n310), 
        .A3(bpu_gte_x_2_n355), .A4(bpu_gte_x_2_n354), .A5(bpu_gte_x_2_n357), 
        .Y(bpu_gte_x_2_n353) );
  INVX0_LVT bpu_gte_x_2_U259 ( .A(bpu_gte_x_2_n354), .Y(bpu_gte_x_2_n314) );
  INVX0_LVT bpu_gte_x_2_U258 ( .A(bpu_gte_x_2_n367), .Y(bpu_gte_x_2_n310) );
  INVX1_LVT bpu_gte_x_2_U257 ( .A(n_T_918[26]), .Y(bpu_gte_x_2_n327) );
  INVX1_LVT bpu_gte_x_2_U256 ( .A(n_T_918[27]), .Y(bpu_gte_x_2_n306) );
  INVX1_LVT bpu_gte_x_2_U255 ( .A(n_T_918[28]), .Y(bpu_gte_x_2_n326) );
  INVX1_LVT bpu_gte_x_2_U254 ( .A(n_T_918[29]), .Y(bpu_gte_x_2_n325) );
  INVX1_LVT bpu_gte_x_2_U253 ( .A(n_T_918[30]), .Y(bpu_gte_x_2_n324) );
  INVX1_LVT bpu_gte_x_2_U252 ( .A(n_T_918[18]), .Y(bpu_gte_x_2_n334) );
  INVX1_LVT bpu_gte_x_2_U251 ( .A(n_T_918[21]), .Y(bpu_gte_x_2_n332) );
  INVX1_LVT bpu_gte_x_2_U250 ( .A(n_T_918[22]), .Y(bpu_gte_x_2_n331) );
  INVX1_LVT bpu_gte_x_2_U249 ( .A(n_T_918[20]), .Y(bpu_gte_x_2_n333) );
  INVX1_LVT bpu_gte_x_2_U248 ( .A(n_T_918[16]), .Y(bpu_gte_x_2_n336) );
  INVX1_LVT bpu_gte_x_2_U247 ( .A(n_T_918[23]), .Y(bpu_gte_x_2_n330) );
  INVX1_LVT bpu_gte_x_2_U246 ( .A(n_T_918[24]), .Y(bpu_gte_x_2_n329) );
  INVX1_LVT bpu_gte_x_2_U245 ( .A(n_T_918[25]), .Y(bpu_gte_x_2_n328) );
  INVX1_LVT bpu_gte_x_2_U244 ( .A(n_T_918[17]), .Y(bpu_gte_x_2_n335) );
  INVX1_LVT bpu_gte_x_2_U243 ( .A(n_T_918[36]), .Y(bpu_gte_x_2_n318) );
  INVX1_LVT bpu_gte_x_2_U242 ( .A(n_T_918[35]), .Y(bpu_gte_x_2_n319) );
  INVX1_LVT bpu_gte_x_2_U241 ( .A(n_T_918[33]), .Y(bpu_gte_x_2_n321) );
  INVX1_LVT bpu_gte_x_2_U240 ( .A(n_T_918[34]), .Y(bpu_gte_x_2_n320) );
  INVX1_LVT bpu_gte_x_2_U239 ( .A(n_T_918[32]), .Y(bpu_gte_x_2_n322) );
  INVX1_LVT bpu_gte_x_2_U238 ( .A(n_T_918[31]), .Y(bpu_gte_x_2_n323) );
  INVX1_LVT bpu_gte_x_2_U237 ( .A(n_T_918[4]), .Y(bpu_gte_x_2_n345) );
  INVX1_LVT bpu_gte_x_2_U236 ( .A(n_T_918[5]), .Y(bpu_gte_x_2_n344) );
  INVX1_LVT bpu_gte_x_2_U235 ( .A(n_T_918[6]), .Y(bpu_gte_x_2_n343) );
  INVX1_LVT bpu_gte_x_2_U234 ( .A(n_T_918[8]), .Y(bpu_gte_x_2_n342) );
  INVX1_LVT bpu_gte_x_2_U233 ( .A(n_T_918[9]), .Y(bpu_gte_x_2_n341) );
  INVX1_LVT bpu_gte_x_2_U232 ( .A(n_T_918[10]), .Y(bpu_gte_x_2_n340) );
  INVX1_LVT bpu_gte_x_2_U231 ( .A(n_T_918[14]), .Y(bpu_gte_x_2_n337) );
  INVX1_LVT bpu_gte_x_2_U230 ( .A(n_T_918[12]), .Y(bpu_gte_x_2_n339) );
  INVX1_LVT bpu_gte_x_2_U229 ( .A(n_T_918[13]), .Y(bpu_gte_x_2_n338) );
  INVX1_LVT bpu_gte_x_2_U228 ( .A(csr_io_bp_0_address[7]), .Y(bpu_gte_x_2_n317) );
  INVX1_LVT bpu_gte_x_2_U227 ( .A(csr_io_bp_0_address[15]), .Y(
        bpu_gte_x_2_n316) );
  INVX1_LVT bpu_gte_x_2_U226 ( .A(csr_io_bp_0_address[37]), .Y(
        bpu_gte_x_2_n309) );
  INVX1_LVT bpu_gte_x_2_U225 ( .A(csr_io_bp_0_address[38]), .Y(
        bpu_gte_x_2_n311) );
  INVX0_LVT bpu_gte_x_2_U224 ( .A(bpu_gte_x_2_n396), .Y(bpu_gte_x_2_n303) );
  INVX0_LVT bpu_gte_x_2_U223 ( .A(n_T_918[11]), .Y(bpu_gte_x_2_n302) );
  INVX0_LVT bpu_gte_x_2_U221 ( .A(bpu_gte_x_2_n410), .Y(bpu_gte_x_2_n300) );
  INVX0_LVT bpu_gte_x_2_U220 ( .A(n_T_918[19]), .Y(bpu_gte_x_2_n299) );
  NAND3X0_LVT bpu_gte_x_2_U218 ( .A1(bpu_gte_x_2_n297), .A2(bpu_gte_x_2_n385), 
        .A3(bpu_gte_x_2_n296), .Y(bpu_gte_x_2_n378) );
  NAND2X0_LVT bpu_gte_x_2_U217 ( .A1(bpu_gte_x_2_n294), .A2(bpu_gte_x_2_n291), 
        .Y(bpu_gte_x_2_n297) );
  NAND2X0_LVT bpu_gte_x_2_U216 ( .A1(csr_io_bp_0_address[3]), .A2(
        bpu_gte_x_2_n295), .Y(bpu_gte_x_2_n296) );
  INVX0_LVT bpu_gte_x_2_U215 ( .A(n_T_918[3]), .Y(bpu_gte_x_2_n295) );
  OA22X1_LVT bpu_gte_x_2_U214 ( .A1(csr_io_bp_0_address[1]), .A2(
        bpu_gte_x_2_n293), .A3(csr_io_bp_0_address[2]), .A4(bpu_gte_x_2_n290), 
        .Y(bpu_gte_x_2_n294) );
  NAND2X0_LVT bpu_gte_x_2_U213 ( .A1(n_T_918[1]), .A2(bpu_gte_x_2_n292), .Y(
        bpu_gte_x_2_n293) );
  NAND2X0_LVT bpu_gte_x_2_U212 ( .A1(csr_io_bp_0_address[2]), .A2(
        bpu_gte_x_2_n290), .Y(bpu_gte_x_2_n292) );
  AO222X1_LVT bpu_gte_x_2_U211 ( .A1(bpu_gte_x_2_n288), .A2(
        csr_io_bp_0_address[0]), .A3(bpu_gte_x_2_n289), .A4(
        csr_io_bp_0_address[1]), .A5(bpu_gte_x_2_n290), .A6(
        csr_io_bp_0_address[2]), .Y(bpu_gte_x_2_n291) );
  INVX0_LVT bpu_gte_x_2_U210 ( .A(n_T_918[2]), .Y(bpu_gte_x_2_n290) );
  INVX0_LVT bpu_gte_x_2_U209 ( .A(n_T_918[1]), .Y(bpu_gte_x_2_n289) );
  INVX0_LVT bpu_gte_x_2_U208 ( .A(n_T_918[0]), .Y(bpu_gte_x_2_n288) );
  OA222X1_LVT bpu_gte_x_2_U207 ( .A1(bpu_gte_x_2_n285), .A2(
        csr_io_bp_0_address[9]), .A3(bpu_gte_x_2_n340), .A4(
        csr_io_bp_0_address[10]), .A5(bpu_gte_x_2_n386), .A6(bpu_gte_x_2_n287), 
        .Y(bpu_gte_x_2_n392) );
  OA22X1_LVT bpu_gte_x_2_U206 ( .A1(csr_io_bp_0_address[8]), .A2(
        bpu_gte_x_2_n342), .A3(csr_io_bp_0_address[7]), .A4(bpu_gte_x_2_n286), 
        .Y(bpu_gte_x_2_n287) );
  NAND2X0_LVT bpu_gte_x_2_U205 ( .A1(bpu_gte_x_2_n389), .A2(n_T_918[7]), .Y(
        bpu_gte_x_2_n286) );
  NAND2X0_LVT bpu_gte_x_2_U204 ( .A1(n_T_918[9]), .A2(bpu_gte_x_2_n284), .Y(
        bpu_gte_x_2_n285) );
  NAND2X0_LVT bpu_gte_x_2_U203 ( .A1(bpu_gte_x_2_n340), .A2(
        csr_io_bp_0_address[10]), .Y(bpu_gte_x_2_n284) );
  AO221X1_LVT bpu_gte_x_2_U202 ( .A1(1'b1), .A2(bpu_gte_x_2_n399), .A3(
        csr_io_bp_0_address[19]), .A4(bpu_gte_x_2_n299), .A5(bpu_gte_x_2_n300), 
        .Y(bpu_gte_x_2_n375) );
  AO221X1_LVT bpu_gte_x_2_U201 ( .A1(1'b1), .A2(bpu_gte_x_2_n390), .A3(
        csr_io_bp_0_address[11]), .A4(bpu_gte_x_2_n302), .A5(bpu_gte_x_2_n303), 
        .Y(bpu_gte_x_2_n387) );
  AO21X1_LVT alu_U803 ( .A1(alu_n602), .A2(alu_n608), .A3(alu_n601), .Y(
        alu_io_out[62]) );
  NAND3X0_LVT alu_U802 ( .A1(alu_n115), .A2(alu_n600), .A3(alu_n599), .Y(
        alu_n601) );
  NAND2X0_LVT alu_U801 ( .A1(alu_n_T_101_1_), .A2(alu_n598), .Y(alu_n599) );
  AND3X1_LVT alu_U800 ( .A1(alu_n597), .A2(alu_n596), .A3(alu_n595), .Y(
        alu_n600) );
  NAND3X0_LVT alu_U799 ( .A1(alu_io_in2[62]), .A2(alu_n603), .A3(
        alu_io_in1[62]), .Y(alu_n595) );
  NAND2X0_LVT alu_U798 ( .A1(alu_n594), .A2(alu_n593), .Y(alu_n596) );
  NAND2X0_LVT alu_U797 ( .A1(alu_n_T_101_62_), .A2(alu_n124), .Y(alu_n597) );
  AO21X1_LVT alu_U796 ( .A1(alu_n602), .A2(alu_n609), .A3(alu_n592), .Y(
        alu_io_out[61]) );
  NAND4X0_LVT alu_U795 ( .A1(alu_n115), .A2(alu_n591), .A3(alu_n590), .A4(
        alu_n589), .Y(alu_n592) );
  NAND2X0_LVT alu_U794 ( .A1(alu_n_T_101_2_), .A2(alu_n598), .Y(alu_n589) );
  NAND2X0_LVT alu_U793 ( .A1(alu_n_T_101_61_), .A2(alu_n124), .Y(alu_n590) );
  OA21X1_LVT alu_U792 ( .A1(alu_n605), .A2(alu_n588), .A3(alu_n587), .Y(
        alu_n591) );
  NAND3X0_LVT alu_U791 ( .A1(alu_io_in2[61]), .A2(alu_n603), .A3(
        alu_io_in1[61]), .Y(alu_n587) );
  NAND3X0_LVT alu_U790 ( .A1(alu_n586), .A2(alu_n585), .A3(alu_n115), .Y(
        alu_io_out[60]) );
  AND4X1_LVT alu_U789 ( .A1(alu_n584), .A2(alu_n583), .A3(alu_n582), .A4(
        alu_n581), .Y(alu_n585) );
  NAND3X0_LVT alu_U788 ( .A1(alu_io_in2[60]), .A2(alu_n603), .A3(
        alu_io_in1[60]), .Y(alu_n581) );
  NAND2X0_LVT alu_U787 ( .A1(alu_n580), .A2(alu_n593), .Y(alu_n582) );
  NAND2X0_LVT alu_U786 ( .A1(alu_n_T_101_60_), .A2(alu_n124), .Y(alu_n583) );
  NAND2X0_LVT alu_U785 ( .A1(alu_n_T_101_3_), .A2(alu_n598), .Y(alu_n584) );
  NAND2X0_LVT alu_U784 ( .A1(alu_n610), .A2(alu_n602), .Y(alu_n586) );
  NAND3X0_LVT alu_U783 ( .A1(alu_n579), .A2(alu_n578), .A3(alu_n115), .Y(
        alu_io_out[59]) );
  AND4X1_LVT alu_U782 ( .A1(alu_n577), .A2(alu_n576), .A3(alu_n575), .A4(
        alu_n574), .Y(alu_n578) );
  NAND3X0_LVT alu_U781 ( .A1(alu_io_in2[59]), .A2(alu_n603), .A3(
        alu_io_in1[59]), .Y(alu_n574) );
  NAND2X0_LVT alu_U780 ( .A1(alu_n573), .A2(alu_n593), .Y(alu_n575) );
  NAND2X0_LVT alu_U779 ( .A1(alu_n_T_101_4_), .A2(alu_n598), .Y(alu_n576) );
  NAND2X0_LVT alu_U778 ( .A1(alu_n_T_101_59_), .A2(alu_n124), .Y(alu_n577) );
  NAND2X0_LVT alu_U777 ( .A1(alu_n611), .A2(alu_n602), .Y(alu_n579) );
  AO21X1_LVT alu_U776 ( .A1(alu_n602), .A2(alu_n612), .A3(alu_n572), .Y(
        alu_io_out[58]) );
  NAND4X0_LVT alu_U775 ( .A1(alu_n115), .A2(alu_n571), .A3(alu_n570), .A4(
        alu_n569), .Y(alu_n572) );
  NAND2X0_LVT alu_U774 ( .A1(alu_n_T_101_58_), .A2(alu_n124), .Y(alu_n569) );
  NAND2X0_LVT alu_U773 ( .A1(alu_n_T_101_5_), .A2(alu_n598), .Y(alu_n570) );
  OA21X1_LVT alu_U772 ( .A1(alu_n605), .A2(alu_n568), .A3(alu_n567), .Y(
        alu_n571) );
  NAND3X0_LVT alu_U771 ( .A1(alu_io_in2[58]), .A2(alu_n603), .A3(
        alu_io_in1[58]), .Y(alu_n567) );
  AO21X1_LVT alu_U770 ( .A1(alu_n602), .A2(alu_n613), .A3(alu_n566), .Y(
        alu_io_out[57]) );
  NAND4X0_LVT alu_U769 ( .A1(alu_n115), .A2(alu_n565), .A3(alu_n564), .A4(
        alu_n563), .Y(alu_n566) );
  NAND2X0_LVT alu_U768 ( .A1(alu_n_T_101_6_), .A2(alu_n598), .Y(alu_n563) );
  NAND2X0_LVT alu_U767 ( .A1(alu_n_T_101_57_), .A2(alu_n124), .Y(alu_n564) );
  OA21X1_LVT alu_U766 ( .A1(alu_n605), .A2(alu_n562), .A3(alu_n561), .Y(
        alu_n565) );
  NAND3X0_LVT alu_U765 ( .A1(alu_io_in2[57]), .A2(alu_n603), .A3(
        alu_io_in1[57]), .Y(alu_n561) );
  AO21X1_LVT alu_U764 ( .A1(alu_n602), .A2(alu_n614), .A3(alu_n560), .Y(
        alu_io_out[56]) );
  NAND4X0_LVT alu_U763 ( .A1(alu_n115), .A2(alu_n559), .A3(alu_n558), .A4(
        alu_n557), .Y(alu_n560) );
  NAND2X0_LVT alu_U762 ( .A1(alu_n_T_101_56_), .A2(alu_n124), .Y(alu_n557) );
  NAND2X0_LVT alu_U761 ( .A1(alu_n_T_101_7_), .A2(alu_n598), .Y(alu_n558) );
  OA21X1_LVT alu_U760 ( .A1(alu_n605), .A2(alu_n556), .A3(alu_n555), .Y(
        alu_n559) );
  NAND3X0_LVT alu_U759 ( .A1(alu_io_in2[56]), .A2(alu_n603), .A3(
        alu_io_in1[56]), .Y(alu_n555) );
  AO21X1_LVT alu_U758 ( .A1(alu_n602), .A2(alu_n615), .A3(alu_n554), .Y(
        alu_io_out[55]) );
  NAND4X0_LVT alu_U757 ( .A1(alu_n606), .A2(alu_n553), .A3(alu_n552), .A4(
        alu_n551), .Y(alu_n554) );
  NAND2X0_LVT alu_U756 ( .A1(alu_n_T_101_8_), .A2(alu_n598), .Y(alu_n551) );
  NAND2X0_LVT alu_U755 ( .A1(alu_n_T_101_55_), .A2(alu_n124), .Y(alu_n552) );
  OA21X1_LVT alu_U754 ( .A1(alu_n605), .A2(alu_n550), .A3(alu_n549), .Y(
        alu_n553) );
  NAND3X0_LVT alu_U753 ( .A1(alu_io_in2[55]), .A2(alu_n603), .A3(
        alu_io_in1[55]), .Y(alu_n549) );
  AO21X1_LVT alu_U752 ( .A1(alu_n602), .A2(alu_n616), .A3(alu_n548), .Y(
        alu_io_out[54]) );
  NAND4X0_LVT alu_U751 ( .A1(alu_n606), .A2(alu_n547), .A3(alu_n546), .A4(
        alu_n545), .Y(alu_n548) );
  NAND2X0_LVT alu_U750 ( .A1(alu_n_T_101_54_), .A2(alu_n124), .Y(alu_n545) );
  NAND2X0_LVT alu_U749 ( .A1(alu_n_T_101_9_), .A2(alu_n598), .Y(alu_n546) );
  OA21X1_LVT alu_U748 ( .A1(alu_n605), .A2(alu_n544), .A3(alu_n543), .Y(
        alu_n547) );
  NAND3X0_LVT alu_U747 ( .A1(alu_io_in2[54]), .A2(alu_n603), .A3(
        alu_io_in1[54]), .Y(alu_n543) );
  AO21X1_LVT alu_U746 ( .A1(alu_n602), .A2(alu_n617), .A3(alu_n542), .Y(
        alu_io_out[53]) );
  NAND4X0_LVT alu_U745 ( .A1(alu_n606), .A2(alu_n541), .A3(alu_n540), .A4(
        alu_n539), .Y(alu_n542) );
  NAND2X0_LVT alu_U744 ( .A1(alu_n_T_101_10_), .A2(alu_n598), .Y(alu_n539) );
  NAND2X0_LVT alu_U743 ( .A1(alu_n_T_101_53_), .A2(alu_n124), .Y(alu_n540) );
  OA21X1_LVT alu_U742 ( .A1(alu_n605), .A2(alu_n538), .A3(alu_n537), .Y(
        alu_n541) );
  NAND3X0_LVT alu_U741 ( .A1(alu_io_in2[53]), .A2(alu_n603), .A3(
        alu_io_in1[53]), .Y(alu_n537) );
  AO21X1_LVT alu_U740 ( .A1(alu_n602), .A2(alu_n618), .A3(alu_n536), .Y(
        alu_io_out[52]) );
  NAND4X0_LVT alu_U739 ( .A1(alu_n606), .A2(alu_n535), .A3(alu_n534), .A4(
        alu_n533), .Y(alu_n536) );
  NAND2X0_LVT alu_U738 ( .A1(alu_n_T_101_52_), .A2(alu_n124), .Y(alu_n533) );
  NAND2X0_LVT alu_U737 ( .A1(alu_n_T_101_11_), .A2(alu_n598), .Y(alu_n534) );
  OA21X1_LVT alu_U736 ( .A1(alu_n605), .A2(alu_n532), .A3(alu_n531), .Y(
        alu_n535) );
  NAND3X0_LVT alu_U735 ( .A1(alu_io_in2[52]), .A2(alu_n603), .A3(
        alu_io_in1[52]), .Y(alu_n531) );
  AO21X1_LVT alu_U734 ( .A1(alu_n602), .A2(alu_n619), .A3(alu_n530), .Y(
        alu_io_out[51]) );
  NAND4X0_LVT alu_U733 ( .A1(alu_n606), .A2(alu_n529), .A3(alu_n528), .A4(
        alu_n527), .Y(alu_n530) );
  NAND2X0_LVT alu_U732 ( .A1(alu_n_T_101_12_), .A2(alu_n598), .Y(alu_n527) );
  NAND2X0_LVT alu_U731 ( .A1(alu_n_T_101_51_), .A2(alu_n124), .Y(alu_n528) );
  OA21X1_LVT alu_U730 ( .A1(alu_n605), .A2(alu_n526), .A3(alu_n525), .Y(
        alu_n529) );
  NAND3X0_LVT alu_U729 ( .A1(alu_io_in2[51]), .A2(alu_n603), .A3(
        alu_io_in1[51]), .Y(alu_n525) );
  AO21X1_LVT alu_U728 ( .A1(alu_n602), .A2(alu_n620), .A3(alu_n524), .Y(
        alu_io_out[50]) );
  NAND4X0_LVT alu_U727 ( .A1(alu_n606), .A2(alu_n523), .A3(alu_n522), .A4(
        alu_n521), .Y(alu_n524) );
  NAND2X0_LVT alu_U726 ( .A1(alu_n_T_101_50_), .A2(alu_n124), .Y(alu_n521) );
  NAND2X0_LVT alu_U725 ( .A1(alu_n_T_101_13_), .A2(alu_n598), .Y(alu_n522) );
  OA21X1_LVT alu_U724 ( .A1(alu_n605), .A2(alu_n520), .A3(alu_n519), .Y(
        alu_n523) );
  NAND3X0_LVT alu_U723 ( .A1(alu_io_in2[50]), .A2(alu_n603), .A3(
        alu_io_in1[50]), .Y(alu_n519) );
  AO21X1_LVT alu_U722 ( .A1(alu_n602), .A2(alu_n621), .A3(alu_n518), .Y(
        alu_io_out[49]) );
  NAND4X0_LVT alu_U721 ( .A1(alu_n606), .A2(alu_n517), .A3(alu_n516), .A4(
        alu_n515), .Y(alu_n518) );
  NAND2X0_LVT alu_U720 ( .A1(alu_n_T_101_14_), .A2(alu_n598), .Y(alu_n515) );
  NAND2X0_LVT alu_U719 ( .A1(alu_n_T_101_49_), .A2(alu_n124), .Y(alu_n516) );
  OA21X1_LVT alu_U718 ( .A1(alu_n605), .A2(alu_n514), .A3(alu_n513), .Y(
        alu_n517) );
  NAND3X0_LVT alu_U717 ( .A1(alu_io_in2[49]), .A2(alu_n603), .A3(
        alu_io_in1[49]), .Y(alu_n513) );
  AO21X1_LVT alu_U716 ( .A1(alu_n602), .A2(alu_n622), .A3(alu_n512), .Y(
        alu_io_out[48]) );
  NAND4X0_LVT alu_U715 ( .A1(alu_n606), .A2(alu_n511), .A3(alu_n510), .A4(
        alu_n509), .Y(alu_n512) );
  NAND2X0_LVT alu_U714 ( .A1(alu_n_T_101_48_), .A2(alu_n124), .Y(alu_n509) );
  NAND2X0_LVT alu_U713 ( .A1(alu_n_T_101_15_), .A2(alu_n598), .Y(alu_n510) );
  OA21X1_LVT alu_U712 ( .A1(alu_n605), .A2(alu_n508), .A3(alu_n507), .Y(
        alu_n511) );
  NAND3X0_LVT alu_U711 ( .A1(alu_io_in2[48]), .A2(alu_n603), .A3(
        alu_io_in1[48]), .Y(alu_n507) );
  NAND4X0_LVT alu_U710 ( .A1(alu_n606), .A2(alu_n506), .A3(alu_n505), .A4(
        alu_n504), .Y(alu_io_out[47]) );
  NAND2X0_LVT alu_U709 ( .A1(alu_n_T_101_47_), .A2(alu_n124), .Y(alu_n504) );
  OA21X1_LVT alu_U708 ( .A1(alu_n123), .A2(alu_n503), .A3(alu_n502), .Y(
        alu_n505) );
  OA21X1_LVT alu_U707 ( .A1(alu_n605), .A2(alu_n501), .A3(alu_n500), .Y(
        alu_n502) );
  NAND3X0_LVT alu_U706 ( .A1(alu_io_in2[47]), .A2(alu_n603), .A3(
        alu_io_in1[47]), .Y(alu_n500) );
  NAND2X0_LVT alu_U705 ( .A1(alu_n623), .A2(alu_n602), .Y(alu_n506) );
  AO21X1_LVT alu_U704 ( .A1(alu_n602), .A2(alu_n624), .A3(alu_n499), .Y(
        alu_io_out[46]) );
  NAND4X0_LVT alu_U703 ( .A1(alu_n606), .A2(alu_n498), .A3(alu_n497), .A4(
        alu_n496), .Y(alu_n499) );
  NAND2X0_LVT alu_U702 ( .A1(alu_n_T_101_46_), .A2(alu_n124), .Y(alu_n496) );
  NAND2X0_LVT alu_U701 ( .A1(alu_n_T_101_17_), .A2(alu_n598), .Y(alu_n497) );
  OA21X1_LVT alu_U700 ( .A1(alu_n605), .A2(alu_n495), .A3(alu_n494), .Y(
        alu_n498) );
  NAND3X0_LVT alu_U699 ( .A1(alu_io_in2[46]), .A2(alu_n603), .A3(
        alu_io_in1[46]), .Y(alu_n494) );
  AO21X1_LVT alu_U698 ( .A1(alu_n602), .A2(alu_n625), .A3(alu_n493), .Y(
        alu_io_out[45]) );
  NAND4X0_LVT alu_U697 ( .A1(alu_n606), .A2(alu_n492), .A3(alu_n491), .A4(
        alu_n490), .Y(alu_n493) );
  NAND2X0_LVT alu_U696 ( .A1(alu_n_T_101_18_), .A2(alu_n598), .Y(alu_n490) );
  NAND2X0_LVT alu_U695 ( .A1(alu_n_T_101_45_), .A2(alu_n124), .Y(alu_n491) );
  OA21X1_LVT alu_U694 ( .A1(alu_n605), .A2(alu_n489), .A3(alu_n488), .Y(
        alu_n492) );
  NAND3X0_LVT alu_U693 ( .A1(alu_io_in2[45]), .A2(alu_n603), .A3(
        alu_io_in1[45]), .Y(alu_n488) );
  AO21X1_LVT alu_U692 ( .A1(alu_n602), .A2(alu_n626), .A3(alu_n487), .Y(
        alu_io_out[44]) );
  NAND4X0_LVT alu_U691 ( .A1(alu_n115), .A2(alu_n486), .A3(alu_n485), .A4(
        alu_n484), .Y(alu_n487) );
  NAND2X0_LVT alu_U690 ( .A1(alu_n_T_101_44_), .A2(alu_n124), .Y(alu_n484) );
  NAND2X0_LVT alu_U689 ( .A1(alu_n_T_101_19_), .A2(alu_n598), .Y(alu_n485) );
  OA21X1_LVT alu_U688 ( .A1(alu_n605), .A2(alu_n483), .A3(alu_n482), .Y(
        alu_n486) );
  NAND3X0_LVT alu_U687 ( .A1(alu_io_in2[44]), .A2(alu_n603), .A3(
        alu_io_in1[44]), .Y(alu_n482) );
  AO21X1_LVT alu_U686 ( .A1(alu_n602), .A2(alu_n627), .A3(alu_n481), .Y(
        alu_io_out[43]) );
  NAND4X0_LVT alu_U685 ( .A1(alu_n115), .A2(alu_n480), .A3(alu_n479), .A4(
        alu_n478), .Y(alu_n481) );
  NAND2X0_LVT alu_U684 ( .A1(alu_n_T_101_20_), .A2(alu_n598), .Y(alu_n478) );
  NAND2X0_LVT alu_U683 ( .A1(alu_n_T_101_43_), .A2(alu_n124), .Y(alu_n479) );
  OA21X1_LVT alu_U682 ( .A1(alu_n605), .A2(alu_n477), .A3(alu_n476), .Y(
        alu_n480) );
  NAND3X0_LVT alu_U681 ( .A1(alu_io_in2[43]), .A2(alu_n603), .A3(
        alu_io_in1[43]), .Y(alu_n476) );
  AO21X1_LVT alu_U680 ( .A1(alu_n602), .A2(alu_n628), .A3(alu_n475), .Y(
        alu_io_out[42]) );
  NAND4X0_LVT alu_U679 ( .A1(alu_n115), .A2(alu_n474), .A3(alu_n473), .A4(
        alu_n472), .Y(alu_n475) );
  NAND2X0_LVT alu_U678 ( .A1(alu_n_T_101_42_), .A2(alu_n124), .Y(alu_n472) );
  NAND2X0_LVT alu_U677 ( .A1(alu_n_T_101_21_), .A2(alu_n598), .Y(alu_n473) );
  OA21X1_LVT alu_U676 ( .A1(alu_n605), .A2(alu_n471), .A3(alu_n470), .Y(
        alu_n474) );
  NAND3X0_LVT alu_U675 ( .A1(alu_io_in2[42]), .A2(alu_n603), .A3(
        alu_io_in1[42]), .Y(alu_n470) );
  AO21X1_LVT alu_U674 ( .A1(alu_n602), .A2(alu_n629), .A3(alu_n469), .Y(
        alu_io_out[41]) );
  NAND4X0_LVT alu_U673 ( .A1(alu_n115), .A2(alu_n468), .A3(alu_n467), .A4(
        alu_n466), .Y(alu_n469) );
  NAND2X0_LVT alu_U672 ( .A1(alu_n_T_101_22_), .A2(alu_n598), .Y(alu_n466) );
  NAND2X0_LVT alu_U671 ( .A1(alu_n_T_101_41_), .A2(alu_n124), .Y(alu_n467) );
  OA21X1_LVT alu_U670 ( .A1(alu_n605), .A2(alu_n465), .A3(alu_n464), .Y(
        alu_n468) );
  NAND3X0_LVT alu_U669 ( .A1(alu_io_in2[41]), .A2(alu_n603), .A3(
        alu_io_in1[41]), .Y(alu_n464) );
  AO21X1_LVT alu_U668 ( .A1(alu_n602), .A2(alu_n630), .A3(alu_n463), .Y(
        alu_io_out[40]) );
  NAND4X0_LVT alu_U667 ( .A1(alu_n606), .A2(alu_n462), .A3(alu_n461), .A4(
        alu_n460), .Y(alu_n463) );
  NAND2X0_LVT alu_U666 ( .A1(alu_n_T_101_40_), .A2(alu_n124), .Y(alu_n460) );
  NAND2X0_LVT alu_U665 ( .A1(alu_n_T_101_23_), .A2(alu_n598), .Y(alu_n461) );
  OA21X1_LVT alu_U664 ( .A1(alu_n605), .A2(alu_n459), .A3(alu_n458), .Y(
        alu_n462) );
  NAND3X0_LVT alu_U663 ( .A1(alu_io_in2[40]), .A2(alu_n603), .A3(
        alu_io_in1[40]), .Y(alu_n458) );
  NAND4X0_LVT alu_U662 ( .A1(alu_n115), .A2(alu_n451), .A3(alu_n450), .A4(
        alu_n449), .Y(alu_io_out[33]) );
  NAND2X0_LVT alu_U661 ( .A1(alu_n_T_101_33_), .A2(alu_n124), .Y(alu_n449) );
  OA21X1_LVT alu_U660 ( .A1(alu_n123), .A2(alu_n448), .A3(alu_n447), .Y(
        alu_n450) );
  OA21X1_LVT alu_U659 ( .A1(alu_n605), .A2(alu_n446), .A3(alu_n445), .Y(
        alu_n447) );
  NAND3X0_LVT alu_U658 ( .A1(alu_io_in2[33]), .A2(alu_n603), .A3(
        alu_io_in1[33]), .Y(alu_n445) );
  NAND2X0_LVT alu_U657 ( .A1(io_dmem_req_bits_addr[33]), .A2(alu_n602), .Y(
        alu_n451) );
  NAND4X0_LVT alu_U656 ( .A1(alu_n444), .A2(alu_n443), .A3(alu_n115), .A4(
        alu_n442), .Y(alu_io_out[32]) );
  NAND2X0_LVT alu_U655 ( .A1(alu_n_T_101_31_), .A2(alu_n598), .Y(alu_n442) );
  NAND2X0_LVT alu_U654 ( .A1(alu_io_out[31]), .A2(alu_n440), .Y(alu_n606) );
  OA21X1_LVT alu_U653 ( .A1(alu_n117), .A2(alu_n439), .A3(alu_n438), .Y(
        alu_n443) );
  OA21X1_LVT alu_U652 ( .A1(alu_n605), .A2(alu_n437), .A3(alu_n436), .Y(
        alu_n438) );
  NAND3X0_LVT alu_U651 ( .A1(alu_io_in2[32]), .A2(alu_n603), .A3(
        alu_io_in1[32]), .Y(alu_n436) );
  AND2X1_LVT alu_U650 ( .A1(alu_n435), .A2(alu_io_dw), .Y(alu_n593) );
  NAND2X0_LVT alu_U649 ( .A1(io_dmem_req_bits_addr[32]), .A2(alu_n602), .Y(
        alu_n444) );
  AO21X1_LVT alu_U648 ( .A1(alu_n434), .A2(io_dmem_req_bits_addr[31]), .A3(
        alu_n433), .Y(alu_io_out[31]) );
  NAND4X0_LVT alu_U647 ( .A1(alu_n432), .A2(alu_n431), .A3(alu_n430), .A4(
        alu_n429), .Y(alu_n433) );
  NAND3X0_LVT alu_U646 ( .A1(alu_io_in2[31]), .A2(alu_n122), .A3(
        alu_io_in1[31]), .Y(alu_n429) );
  NAND2X0_LVT alu_U645 ( .A1(alu_n428), .A2(alu_n435), .Y(alu_n430) );
  NAND2X0_LVT alu_U644 ( .A1(alu_n_T_101_32_), .A2(alu_n441), .Y(alu_n431) );
  NAND2X0_LVT alu_U643 ( .A1(alu_n_T_101_31_), .A2(alu_n121), .Y(alu_n432) );
  NAND4X0_LVT alu_U642 ( .A1(alu_n427), .A2(alu_n426), .A3(alu_n425), .A4(
        alu_n424), .Y(alu_io_out[30]) );
  NAND2X0_LVT alu_U641 ( .A1(alu_n_T_101_30_), .A2(alu_n121), .Y(alu_n424) );
  NAND2X0_LVT alu_U640 ( .A1(alu_n_T_101_33_), .A2(alu_n441), .Y(alu_n425) );
  OA21X1_LVT alu_U639 ( .A1(alu_n423), .A2(alu_n422), .A3(alu_n421), .Y(
        alu_n426) );
  NAND3X0_LVT alu_U638 ( .A1(alu_io_in2[30]), .A2(alu_n122), .A3(
        alu_io_in1[30]), .Y(alu_n421) );
  NAND2X0_LVT alu_U637 ( .A1(io_dmem_req_bits_addr[30]), .A2(alu_n434), .Y(
        alu_n427) );
  NAND4X0_LVT alu_U636 ( .A1(alu_n420), .A2(alu_n419), .A3(alu_n418), .A4(
        alu_n417), .Y(alu_io_out[29]) );
  NAND2X0_LVT alu_U635 ( .A1(alu_n_T_101_34_), .A2(alu_n441), .Y(alu_n417) );
  NAND2X0_LVT alu_U634 ( .A1(alu_n_T_101_29_), .A2(alu_n121), .Y(alu_n418) );
  OA21X1_LVT alu_U633 ( .A1(alu_n423), .A2(alu_n416), .A3(alu_n415), .Y(
        alu_n419) );
  NAND3X0_LVT alu_U632 ( .A1(alu_io_in2[29]), .A2(alu_n122), .A3(
        alu_io_in1[29]), .Y(alu_n415) );
  NAND2X0_LVT alu_U631 ( .A1(io_dmem_req_bits_addr[29]), .A2(alu_n434), .Y(
        alu_n420) );
  NAND4X0_LVT alu_U630 ( .A1(alu_n414), .A2(alu_n413), .A3(alu_n412), .A4(
        alu_n411), .Y(alu_io_out[28]) );
  NAND2X0_LVT alu_U629 ( .A1(alu_n_T_101_28_), .A2(alu_n121), .Y(alu_n411) );
  NAND2X0_LVT alu_U628 ( .A1(alu_n_T_101_35_), .A2(alu_n441), .Y(alu_n412) );
  OA21X1_LVT alu_U627 ( .A1(alu_n423), .A2(alu_n410), .A3(alu_n409), .Y(
        alu_n413) );
  NAND3X0_LVT alu_U626 ( .A1(alu_io_in2[28]), .A2(alu_n122), .A3(
        alu_io_in1[28]), .Y(alu_n409) );
  NAND2X0_LVT alu_U625 ( .A1(io_dmem_req_bits_addr[28]), .A2(alu_n434), .Y(
        alu_n414) );
  NAND4X0_LVT alu_U624 ( .A1(alu_n408), .A2(alu_n407), .A3(alu_n406), .A4(
        alu_n405), .Y(alu_io_out[27]) );
  NAND2X0_LVT alu_U623 ( .A1(alu_n_T_101_36_), .A2(alu_n441), .Y(alu_n405) );
  NAND2X0_LVT alu_U622 ( .A1(alu_n_T_101_27_), .A2(alu_n121), .Y(alu_n406) );
  OA21X1_LVT alu_U621 ( .A1(alu_n423), .A2(alu_n404), .A3(alu_n403), .Y(
        alu_n407) );
  NAND3X0_LVT alu_U620 ( .A1(alu_io_in2[27]), .A2(alu_n122), .A3(
        alu_io_in1[27]), .Y(alu_n403) );
  NAND2X0_LVT alu_U619 ( .A1(io_dmem_req_bits_addr[27]), .A2(alu_n434), .Y(
        alu_n408) );
  NAND4X0_LVT alu_U618 ( .A1(alu_n402), .A2(alu_n401), .A3(alu_n400), .A4(
        alu_n399), .Y(alu_io_out[26]) );
  NAND2X0_LVT alu_U617 ( .A1(alu_n_T_101_26_), .A2(alu_n121), .Y(alu_n399) );
  NAND2X0_LVT alu_U616 ( .A1(alu_n_T_101_37_), .A2(alu_n441), .Y(alu_n400) );
  OA21X1_LVT alu_U615 ( .A1(alu_n423), .A2(alu_n398), .A3(alu_n397), .Y(
        alu_n401) );
  NAND3X0_LVT alu_U614 ( .A1(alu_io_in2[26]), .A2(alu_n122), .A3(
        alu_io_in1[26]), .Y(alu_n397) );
  NAND2X0_LVT alu_U613 ( .A1(io_dmem_req_bits_addr[26]), .A2(alu_n434), .Y(
        alu_n402) );
  NAND4X0_LVT alu_U612 ( .A1(alu_n396), .A2(alu_n395), .A3(alu_n394), .A4(
        alu_n393), .Y(alu_io_out[25]) );
  NAND2X0_LVT alu_U611 ( .A1(alu_n_T_101_38_), .A2(alu_n441), .Y(alu_n393) );
  NAND2X0_LVT alu_U610 ( .A1(alu_n_T_101_25_), .A2(alu_n121), .Y(alu_n394) );
  OA21X1_LVT alu_U609 ( .A1(alu_n423), .A2(alu_n392), .A3(alu_n391), .Y(
        alu_n395) );
  NAND3X0_LVT alu_U608 ( .A1(alu_io_in2[25]), .A2(alu_n122), .A3(
        alu_io_in1[25]), .Y(alu_n391) );
  NAND2X0_LVT alu_U607 ( .A1(io_dmem_req_bits_addr[25]), .A2(alu_n434), .Y(
        alu_n396) );
  NAND4X0_LVT alu_U606 ( .A1(alu_n390), .A2(alu_n389), .A3(alu_n388), .A4(
        alu_n387), .Y(alu_io_out[24]) );
  NAND2X0_LVT alu_U605 ( .A1(alu_n_T_101_24_), .A2(alu_n121), .Y(alu_n387) );
  NAND2X0_LVT alu_U604 ( .A1(alu_n_T_101_39_), .A2(alu_n441), .Y(alu_n388) );
  OA21X1_LVT alu_U603 ( .A1(alu_n423), .A2(alu_n386), .A3(alu_n385), .Y(
        alu_n389) );
  NAND3X0_LVT alu_U602 ( .A1(alu_io_in2[24]), .A2(alu_n122), .A3(
        alu_io_in1[24]), .Y(alu_n385) );
  NAND2X0_LVT alu_U601 ( .A1(io_dmem_req_bits_addr[24]), .A2(alu_n434), .Y(
        alu_n390) );
  NAND4X0_LVT alu_U600 ( .A1(alu_n384), .A2(alu_n383), .A3(alu_n382), .A4(
        alu_n381), .Y(alu_io_out[23]) );
  NAND2X0_LVT alu_U599 ( .A1(alu_n_T_101_40_), .A2(alu_n441), .Y(alu_n381) );
  NAND2X0_LVT alu_U598 ( .A1(alu_n_T_101_23_), .A2(alu_n121), .Y(alu_n382) );
  OA21X1_LVT alu_U597 ( .A1(alu_n423), .A2(alu_n380), .A3(alu_n379), .Y(
        alu_n383) );
  NAND3X0_LVT alu_U596 ( .A1(alu_io_in2[23]), .A2(alu_n122), .A3(
        alu_io_in1[23]), .Y(alu_n379) );
  NAND2X0_LVT alu_U595 ( .A1(io_dmem_req_bits_addr[23]), .A2(alu_n434), .Y(
        alu_n384) );
  NAND4X0_LVT alu_U594 ( .A1(alu_n378), .A2(alu_n377), .A3(alu_n376), .A4(
        alu_n375), .Y(alu_io_out[22]) );
  NAND2X0_LVT alu_U593 ( .A1(alu_n_T_101_22_), .A2(alu_n121), .Y(alu_n375) );
  NAND2X0_LVT alu_U592 ( .A1(alu_n_T_101_41_), .A2(alu_n441), .Y(alu_n376) );
  OA21X1_LVT alu_U591 ( .A1(alu_n423), .A2(alu_n374), .A3(alu_n373), .Y(
        alu_n377) );
  NAND3X0_LVT alu_U590 ( .A1(alu_io_in2[22]), .A2(alu_n122), .A3(
        alu_io_in1[22]), .Y(alu_n373) );
  NAND2X0_LVT alu_U589 ( .A1(io_dmem_req_bits_addr[22]), .A2(alu_n434), .Y(
        alu_n378) );
  NAND4X0_LVT alu_U588 ( .A1(alu_n372), .A2(alu_n371), .A3(alu_n370), .A4(
        alu_n369), .Y(alu_io_out[21]) );
  NAND2X0_LVT alu_U587 ( .A1(alu_n_T_101_42_), .A2(alu_n441), .Y(alu_n369) );
  NAND2X0_LVT alu_U586 ( .A1(alu_n_T_101_21_), .A2(alu_n121), .Y(alu_n370) );
  OA21X1_LVT alu_U585 ( .A1(alu_n423), .A2(alu_n368), .A3(alu_n367), .Y(
        alu_n371) );
  NAND3X0_LVT alu_U584 ( .A1(alu_io_in2[21]), .A2(alu_n122), .A3(
        alu_io_in1[21]), .Y(alu_n367) );
  NAND2X0_LVT alu_U583 ( .A1(io_dmem_req_bits_addr[21]), .A2(alu_n434), .Y(
        alu_n372) );
  NAND4X0_LVT alu_U582 ( .A1(alu_n366), .A2(alu_n365), .A3(alu_n364), .A4(
        alu_n363), .Y(alu_io_out[20]) );
  NAND2X0_LVT alu_U581 ( .A1(alu_n_T_101_20_), .A2(alu_n121), .Y(alu_n363) );
  NAND2X0_LVT alu_U580 ( .A1(alu_n_T_101_43_), .A2(alu_n441), .Y(alu_n364) );
  OA21X1_LVT alu_U579 ( .A1(alu_n423), .A2(alu_n362), .A3(alu_n361), .Y(
        alu_n365) );
  NAND3X0_LVT alu_U578 ( .A1(alu_io_in2[20]), .A2(alu_n122), .A3(
        alu_io_in1[20]), .Y(alu_n361) );
  NAND2X0_LVT alu_U577 ( .A1(io_dmem_req_bits_addr[20]), .A2(alu_n434), .Y(
        alu_n366) );
  NAND4X0_LVT alu_U576 ( .A1(alu_n360), .A2(alu_n359), .A3(alu_n358), .A4(
        alu_n357), .Y(alu_io_out[19]) );
  NAND2X0_LVT alu_U575 ( .A1(alu_n_T_101_44_), .A2(alu_n441), .Y(alu_n357) );
  NAND2X0_LVT alu_U574 ( .A1(alu_n_T_101_19_), .A2(alu_n121), .Y(alu_n358) );
  OA21X1_LVT alu_U573 ( .A1(alu_n423), .A2(alu_n356), .A3(alu_n355), .Y(
        alu_n359) );
  NAND3X0_LVT alu_U572 ( .A1(alu_io_in2[19]), .A2(alu_n122), .A3(
        alu_io_in1[19]), .Y(alu_n355) );
  NAND2X0_LVT alu_U571 ( .A1(io_dmem_req_bits_addr[19]), .A2(alu_n434), .Y(
        alu_n360) );
  NAND4X0_LVT alu_U570 ( .A1(alu_n354), .A2(alu_n353), .A3(alu_n352), .A4(
        alu_n351), .Y(alu_io_out[18]) );
  NAND2X0_LVT alu_U569 ( .A1(alu_n_T_101_18_), .A2(alu_n121), .Y(alu_n351) );
  NAND2X0_LVT alu_U568 ( .A1(alu_n_T_101_45_), .A2(alu_n441), .Y(alu_n352) );
  OA21X1_LVT alu_U567 ( .A1(alu_n423), .A2(alu_n350), .A3(alu_n349), .Y(
        alu_n353) );
  NAND3X0_LVT alu_U566 ( .A1(alu_io_in2[18]), .A2(alu_n122), .A3(
        alu_io_in1[18]), .Y(alu_n349) );
  NAND2X0_LVT alu_U565 ( .A1(io_dmem_req_bits_addr[18]), .A2(alu_n434), .Y(
        alu_n354) );
  NAND4X0_LVT alu_U564 ( .A1(alu_n348), .A2(alu_n347), .A3(alu_n346), .A4(
        alu_n345), .Y(alu_io_out[17]) );
  NAND2X0_LVT alu_U563 ( .A1(alu_n_T_101_46_), .A2(alu_n441), .Y(alu_n345) );
  NAND2X0_LVT alu_U562 ( .A1(alu_n_T_101_17_), .A2(alu_n121), .Y(alu_n346) );
  OA21X1_LVT alu_U561 ( .A1(alu_n423), .A2(alu_n344), .A3(alu_n343), .Y(
        alu_n347) );
  NAND3X0_LVT alu_U560 ( .A1(alu_io_in2[17]), .A2(alu_n122), .A3(
        alu_io_in1[17]), .Y(alu_n343) );
  NAND2X0_LVT alu_U559 ( .A1(io_dmem_req_bits_addr[17]), .A2(alu_n434), .Y(
        alu_n348) );
  NAND4X0_LVT alu_U558 ( .A1(alu_n342), .A2(alu_n341), .A3(alu_n340), .A4(
        alu_n339), .Y(alu_io_out[16]) );
  NAND2X0_LVT alu_U557 ( .A1(alu_n_T_101_16_), .A2(alu_n121), .Y(alu_n339) );
  NAND2X0_LVT alu_U556 ( .A1(alu_n_T_101_47_), .A2(alu_n441), .Y(alu_n340) );
  OA21X1_LVT alu_U555 ( .A1(alu_n423), .A2(alu_n338), .A3(alu_n337), .Y(
        alu_n341) );
  NAND3X0_LVT alu_U554 ( .A1(alu_io_in2[16]), .A2(alu_n122), .A3(
        alu_io_in1[16]), .Y(alu_n337) );
  NAND2X0_LVT alu_U553 ( .A1(io_dmem_req_bits_addr[16]), .A2(alu_n434), .Y(
        alu_n342) );
  AO21X1_LVT alu_U552 ( .A1(io_dmem_req_bits_addr[15]), .A2(alu_n434), .A3(
        alu_n336), .Y(alu_io_out[15]) );
  NAND4X0_LVT alu_U551 ( .A1(alu_n335), .A2(alu_n334), .A3(alu_n333), .A4(
        alu_n332), .Y(alu_n336) );
  NAND3X0_LVT alu_U550 ( .A1(alu_io_in2[15]), .A2(alu_n122), .A3(
        alu_io_in1[15]), .Y(alu_n332) );
  OR2X1_LVT alu_U549 ( .A1(alu_n423), .A2(alu_n331), .Y(alu_n333) );
  NAND2X0_LVT alu_U548 ( .A1(alu_n_T_101_48_), .A2(alu_n441), .Y(alu_n334) );
  NAND2X0_LVT alu_U547 ( .A1(alu_n_T_101_15_), .A2(alu_n121), .Y(alu_n335) );
  NAND4X0_LVT alu_U546 ( .A1(alu_n330), .A2(alu_n329), .A3(alu_n328), .A4(
        alu_n327), .Y(alu_io_out[14]) );
  NAND2X0_LVT alu_U545 ( .A1(alu_n_T_101_14_), .A2(alu_n121), .Y(alu_n327) );
  NAND2X0_LVT alu_U544 ( .A1(alu_n_T_101_49_), .A2(alu_n441), .Y(alu_n328) );
  OA21X1_LVT alu_U543 ( .A1(alu_n423), .A2(alu_n326), .A3(alu_n325), .Y(
        alu_n329) );
  NAND3X0_LVT alu_U542 ( .A1(alu_io_in2[14]), .A2(alu_n122), .A3(
        alu_io_in1[14]), .Y(alu_n325) );
  NAND2X0_LVT alu_U541 ( .A1(io_dmem_req_bits_addr[14]), .A2(alu_n434), .Y(
        alu_n330) );
  NAND4X0_LVT alu_U540 ( .A1(alu_n323), .A2(alu_n322), .A3(alu_n321), .A4(
        alu_n320), .Y(alu_io_out[12]) );
  NAND2X0_LVT alu_U539 ( .A1(alu_n_T_101_12_), .A2(alu_n121), .Y(alu_n320) );
  NAND2X0_LVT alu_U538 ( .A1(alu_n_T_101_51_), .A2(alu_n441), .Y(alu_n321) );
  OA21X1_LVT alu_U537 ( .A1(alu_n423), .A2(alu_n319), .A3(alu_n318), .Y(
        alu_n322) );
  NAND3X0_LVT alu_U536 ( .A1(alu_io_in2[12]), .A2(alu_n122), .A3(
        alu_io_in1[12]), .Y(alu_n318) );
  NAND2X0_LVT alu_U535 ( .A1(io_dmem_req_bits_addr[12]), .A2(alu_n434), .Y(
        alu_n323) );
  NAND4X0_LVT alu_U534 ( .A1(alu_n317), .A2(alu_n316), .A3(alu_n315), .A4(
        alu_n314), .Y(alu_io_out[11]) );
  NAND2X0_LVT alu_U533 ( .A1(alu_n_T_101_52_), .A2(alu_n441), .Y(alu_n314) );
  NAND2X0_LVT alu_U532 ( .A1(alu_n_T_101_11_), .A2(alu_n121), .Y(alu_n315) );
  OA21X1_LVT alu_U531 ( .A1(alu_n423), .A2(alu_n313), .A3(alu_n312), .Y(
        alu_n316) );
  NAND3X0_LVT alu_U530 ( .A1(alu_io_in2[11]), .A2(alu_n122), .A3(
        alu_io_in1[11]), .Y(alu_n312) );
  NAND2X0_LVT alu_U529 ( .A1(io_dmem_req_bits_addr[11]), .A2(alu_n434), .Y(
        alu_n317) );
  NAND4X0_LVT alu_U528 ( .A1(alu_n311), .A2(alu_n310), .A3(alu_n309), .A4(
        alu_n308), .Y(alu_io_out[10]) );
  NAND2X0_LVT alu_U527 ( .A1(alu_n_T_101_10_), .A2(alu_n121), .Y(alu_n308) );
  NAND2X0_LVT alu_U526 ( .A1(alu_n_T_101_53_), .A2(alu_n441), .Y(alu_n309) );
  OA21X1_LVT alu_U525 ( .A1(alu_n423), .A2(alu_n307), .A3(alu_n306), .Y(
        alu_n310) );
  NAND3X0_LVT alu_U524 ( .A1(alu_io_in2[10]), .A2(alu_n122), .A3(
        alu_io_in1[10]), .Y(alu_n306) );
  NAND2X0_LVT alu_U523 ( .A1(io_dmem_req_bits_addr[10]), .A2(alu_n434), .Y(
        alu_n311) );
  NAND4X0_LVT alu_U522 ( .A1(alu_n305), .A2(alu_n304), .A3(alu_n303), .A4(
        alu_n302), .Y(alu_io_out[9]) );
  NAND2X0_LVT alu_U521 ( .A1(alu_n_T_101_54_), .A2(alu_n441), .Y(alu_n302) );
  MUX21X1_LVT alu_U520 ( .A1(alu_n301), .A2(alu_n300), .S0(alu_io_in1[9]), .Y(
        alu_n303) );
  OA22X1_LVT alu_U519 ( .A1(alu_io_in2[9]), .A2(alu_n423), .A3(alu_n118), .A4(
        alu_n299), .Y(alu_n300) );
  NAND2X0_LVT alu_U518 ( .A1(alu_io_in2[9]), .A2(alu_n435), .Y(alu_n301) );
  NAND2X0_LVT alu_U517 ( .A1(alu_n_T_101_9_), .A2(alu_n121), .Y(alu_n304) );
  NAND2X0_LVT alu_U516 ( .A1(io_dmem_req_bits_addr[9]), .A2(alu_n434), .Y(
        alu_n305) );
  NAND4X0_LVT alu_U515 ( .A1(alu_n298), .A2(alu_n297), .A3(alu_n296), .A4(
        alu_n295), .Y(alu_io_out[8]) );
  NAND2X0_LVT alu_U514 ( .A1(alu_n_T_101_8_), .A2(alu_n121), .Y(alu_n295) );
  NAND2X0_LVT alu_U513 ( .A1(alu_n_T_101_55_), .A2(alu_n441), .Y(alu_n296) );
  OA21X1_LVT alu_U512 ( .A1(alu_n423), .A2(alu_n294), .A3(alu_n293), .Y(
        alu_n297) );
  NAND3X0_LVT alu_U511 ( .A1(alu_io_in2[8]), .A2(alu_n122), .A3(alu_io_in1[8]), 
        .Y(alu_n293) );
  NAND2X0_LVT alu_U510 ( .A1(io_dmem_req_bits_addr[8]), .A2(alu_n434), .Y(
        alu_n298) );
  NAND4X0_LVT alu_U509 ( .A1(alu_n292), .A2(alu_n291), .A3(alu_n290), .A4(
        alu_n289), .Y(alu_io_out[7]) );
  NAND2X0_LVT alu_U508 ( .A1(alu_n_T_101_56_), .A2(alu_n441), .Y(alu_n289) );
  OA21X1_LVT alu_U507 ( .A1(alu_n423), .A2(alu_n288), .A3(alu_n287), .Y(
        alu_n290) );
  NAND3X0_LVT alu_U506 ( .A1(alu_io_in2[7]), .A2(alu_n122), .A3(alu_io_in1[7]), 
        .Y(alu_n287) );
  NAND2X0_LVT alu_U505 ( .A1(io_dmem_req_bits_addr[7]), .A2(alu_n434), .Y(
        alu_n291) );
  NAND2X0_LVT alu_U504 ( .A1(alu_n_T_101_7_), .A2(alu_n121), .Y(alu_n292) );
  NAND4X0_LVT alu_U503 ( .A1(alu_n286), .A2(alu_n285), .A3(alu_n284), .A4(
        alu_n283), .Y(alu_io_out[6]) );
  NAND2X0_LVT alu_U502 ( .A1(alu_n_T_101_6_), .A2(alu_n121), .Y(alu_n283) );
  NAND2X0_LVT alu_U501 ( .A1(alu_n_T_101_57_), .A2(alu_n441), .Y(alu_n284) );
  OA21X1_LVT alu_U500 ( .A1(alu_n423), .A2(alu_n282), .A3(alu_n281), .Y(
        alu_n285) );
  NAND3X0_LVT alu_U499 ( .A1(alu_io_in2[6]), .A2(alu_n122), .A3(alu_io_in1[6]), 
        .Y(alu_n281) );
  NAND2X0_LVT alu_U498 ( .A1(io_dmem_req_bits_addr[6]), .A2(alu_n434), .Y(
        alu_n286) );
  NAND4X0_LVT alu_U497 ( .A1(alu_n280), .A2(alu_n279), .A3(alu_n278), .A4(
        alu_n277), .Y(alu_io_out[5]) );
  NAND2X0_LVT alu_U496 ( .A1(alu_n_T_101_58_), .A2(alu_n441), .Y(alu_n277) );
  NAND2X0_LVT alu_U495 ( .A1(io_dmem_req_bits_addr[5]), .A2(alu_n434), .Y(
        alu_n278) );
  OA21X1_LVT alu_U494 ( .A1(alu_n423), .A2(alu_n276), .A3(alu_n275), .Y(
        alu_n279) );
  NAND3X0_LVT alu_U493 ( .A1(alu_io_in2[5]), .A2(alu_n122), .A3(alu_io_in1[5]), 
        .Y(alu_n275) );
  NAND2X0_LVT alu_U492 ( .A1(alu_n_T_101_5_), .A2(alu_n121), .Y(alu_n280) );
  NAND4X0_LVT alu_U491 ( .A1(alu_n274), .A2(alu_n273), .A3(alu_n272), .A4(
        alu_n271), .Y(alu_io_out[4]) );
  NAND2X0_LVT alu_U490 ( .A1(io_dmem_req_bits_addr[4]), .A2(alu_n434), .Y(
        alu_n271) );
  NAND2X0_LVT alu_U489 ( .A1(alu_n_T_101_4_), .A2(alu_n121), .Y(alu_n272) );
  OA21X1_LVT alu_U488 ( .A1(alu_n423), .A2(alu_n270), .A3(alu_n269), .Y(
        alu_n273) );
  NAND3X0_LVT alu_U487 ( .A1(alu_io_in2[4]), .A2(alu_n122), .A3(alu_io_in1[4]), 
        .Y(alu_n269) );
  NAND2X0_LVT alu_U486 ( .A1(alu_n_T_101_59_), .A2(alu_n441), .Y(alu_n274) );
  NAND4X0_LVT alu_U485 ( .A1(alu_n268), .A2(alu_n267), .A3(alu_n266), .A4(
        alu_n265), .Y(alu_io_out[3]) );
  NAND2X0_LVT alu_U484 ( .A1(alu_n434), .A2(io_dmem_req_bits_addr[3]), .Y(
        alu_n265) );
  NAND2X0_LVT alu_U483 ( .A1(alu_n_T_101_60_), .A2(alu_n441), .Y(alu_n266) );
  OA21X1_LVT alu_U482 ( .A1(alu_n423), .A2(alu_n264), .A3(alu_n263), .Y(
        alu_n267) );
  NAND3X0_LVT alu_U481 ( .A1(alu_io_in2[3]), .A2(alu_n122), .A3(alu_io_in1[3]), 
        .Y(alu_n263) );
  NAND2X0_LVT alu_U480 ( .A1(alu_n_T_101_3_), .A2(alu_n121), .Y(alu_n268) );
  NAND4X0_LVT alu_U479 ( .A1(alu_n262), .A2(alu_n261), .A3(alu_n260), .A4(
        alu_n259), .Y(alu_io_out[2]) );
  NAND2X0_LVT alu_U478 ( .A1(io_dmem_req_bits_addr[2]), .A2(alu_n434), .Y(
        alu_n259) );
  NAND2X0_LVT alu_U477 ( .A1(alu_n_T_101_2_), .A2(alu_n121), .Y(alu_n260) );
  AOI22X1_LVT alu_U476 ( .A1(alu_io_in2[2]), .A2(alu_n258), .A3(alu_n257), 
        .A4(alu_n435), .Y(alu_n261) );
  AND2X1_LVT alu_U475 ( .A1(alu_io_in1[2]), .A2(alu_n122), .Y(alu_n258) );
  NAND2X0_LVT alu_U474 ( .A1(alu_n_T_101_61_), .A2(alu_n441), .Y(alu_n262) );
  AO21X1_LVT alu_U473 ( .A1(alu_n121), .A2(alu_n_T_101_1_), .A3(alu_n256), .Y(
        alu_io_out[1]) );
  NAND4X0_LVT alu_U472 ( .A1(alu_n255), .A2(alu_n254), .A3(alu_n253), .A4(
        alu_n252), .Y(alu_n256) );
  NAND3X0_LVT alu_U471 ( .A1(alu_io_in2[1]), .A2(alu_n122), .A3(alu_io_in1[1]), 
        .Y(alu_n252) );
  NAND2X0_LVT alu_U470 ( .A1(alu_n251), .A2(alu_n435), .Y(alu_n253) );
  NAND2X0_LVT alu_U469 ( .A1(io_dmem_req_bits_addr[1]), .A2(alu_n434), .Y(
        alu_n254) );
  NAND2X0_LVT alu_U468 ( .A1(alu_n_T_101_62_), .A2(alu_n441), .Y(alu_n255) );
  AO21X1_LVT alu_U467 ( .A1(alu_io_fn[2]), .A2(alu_n250), .A3(alu_n249), .Y(
        alu_io_out[0]) );
  NAND4X0_LVT alu_U466 ( .A1(alu_n248), .A2(alu_n247), .A3(alu_n246), .A4(
        alu_n245), .Y(alu_n249) );
  NAND2X0_LVT alu_U465 ( .A1(io_dmem_req_bits_addr[0]), .A2(alu_n434), .Y(
        alu_n245) );
  NAND2X0_LVT alu_U464 ( .A1(alu_n_T_101_0_), .A2(alu_n121), .Y(alu_n246) );
  OA21X1_LVT alu_U463 ( .A1(alu_n423), .A2(alu_n240), .A3(alu_n239), .Y(
        alu_n247) );
  NAND3X0_LVT alu_U462 ( .A1(alu_io_in2[0]), .A2(alu_n122), .A3(alu_io_in1[0]), 
        .Y(alu_n239) );
  AND3X1_LVT alu_U461 ( .A1(alu_n126), .A2(alu_io_fn[2]), .A3(alu_n237), .Y(
        alu_n435) );
  NAND2X0_LVT alu_U460 ( .A1(alu_n_T_101_63_), .A2(alu_n441), .Y(alu_n248) );
  AND4X1_LVT alu_U459 ( .A1(alu_n241), .A2(alu_n236), .A3(alu_n126), .A4(
        alu_io_fn[0]), .Y(alu_n441) );
  NAND2X0_LVT alu_U458 ( .A1(alu_n234), .A2(alu_n233), .Y(alu_shin_0_) );
  AOI22X1_LVT alu_U457 ( .A1(alu_n121), .A2(alu_io_in1[0]), .A3(alu_io_in1[63]), .A4(alu_n120), .Y(alu_n233) );
  NAND2X0_LVT alu_U456 ( .A1(alu_n234), .A2(alu_n231), .Y(alu_shin_1_) );
  AOI22X1_LVT alu_U455 ( .A1(alu_io_in1[1]), .A2(alu_n121), .A3(alu_io_in1[62]), .A4(alu_n120), .Y(alu_n231) );
  NAND2X0_LVT alu_U454 ( .A1(alu_n234), .A2(alu_n230), .Y(alu_shin_2_) );
  AOI22X1_LVT alu_U453 ( .A1(alu_io_in1[2]), .A2(alu_n121), .A3(alu_io_in1[61]), .A4(alu_n232), .Y(alu_n230) );
  NAND2X0_LVT alu_U452 ( .A1(alu_n234), .A2(alu_n229), .Y(alu_shin_3_) );
  AOI22X1_LVT alu_U451 ( .A1(alu_io_in1[3]), .A2(alu_n121), .A3(alu_io_in1[60]), .A4(alu_n120), .Y(alu_n229) );
  NAND2X0_LVT alu_U450 ( .A1(alu_n234), .A2(alu_n228), .Y(alu_shin_4_) );
  AOI22X1_LVT alu_U449 ( .A1(alu_io_in1[4]), .A2(alu_n121), .A3(alu_io_in1[59]), .A4(alu_n232), .Y(alu_n228) );
  NAND2X0_LVT alu_U448 ( .A1(alu_n234), .A2(alu_n227), .Y(alu_shin_5_) );
  AOI22X1_LVT alu_U447 ( .A1(alu_io_in1[5]), .A2(alu_n121), .A3(alu_io_in1[58]), .A4(alu_n120), .Y(alu_n227) );
  NAND2X0_LVT alu_U446 ( .A1(alu_n234), .A2(alu_n226), .Y(alu_shin_6_) );
  AOI22X1_LVT alu_U445 ( .A1(alu_io_in1[6]), .A2(alu_n121), .A3(alu_io_in1[57]), .A4(alu_n232), .Y(alu_n226) );
  NAND2X0_LVT alu_U444 ( .A1(alu_n234), .A2(alu_n225), .Y(alu_shin_7_) );
  AOI22X1_LVT alu_U443 ( .A1(alu_io_in1[7]), .A2(alu_n121), .A3(alu_io_in1[56]), .A4(alu_n120), .Y(alu_n225) );
  NAND2X0_LVT alu_U442 ( .A1(alu_n234), .A2(alu_n224), .Y(alu_shin_8_) );
  AOI22X1_LVT alu_U441 ( .A1(alu_io_in1[8]), .A2(alu_n121), .A3(alu_io_in1[55]), .A4(alu_n232), .Y(alu_n224) );
  NAND2X0_LVT alu_U440 ( .A1(alu_n234), .A2(alu_n223), .Y(alu_shin_9_) );
  AOI22X1_LVT alu_U439 ( .A1(alu_io_in1[9]), .A2(alu_n121), .A3(alu_io_in1[54]), .A4(alu_n232), .Y(alu_n223) );
  NAND2X0_LVT alu_U438 ( .A1(alu_n234), .A2(alu_n222), .Y(alu_shin_10_) );
  AOI22X1_LVT alu_U437 ( .A1(alu_io_in1[10]), .A2(alu_n121), .A3(
        alu_io_in1[53]), .A4(alu_n232), .Y(alu_n222) );
  NAND2X0_LVT alu_U436 ( .A1(alu_n234), .A2(alu_n221), .Y(alu_shin_11_) );
  AOI22X1_LVT alu_U435 ( .A1(alu_io_in1[11]), .A2(alu_n121), .A3(
        alu_io_in1[52]), .A4(alu_n232), .Y(alu_n221) );
  NAND2X0_LVT alu_U434 ( .A1(alu_n234), .A2(alu_n220), .Y(alu_shin_12_) );
  AOI22X1_LVT alu_U433 ( .A1(alu_io_in1[12]), .A2(alu_n121), .A3(
        alu_io_in1[51]), .A4(alu_n232), .Y(alu_n220) );
  NAND2X0_LVT alu_U432 ( .A1(alu_n234), .A2(alu_n219), .Y(alu_shin_13_) );
  AOI22X1_LVT alu_U431 ( .A1(alu_io_in1[13]), .A2(alu_n121), .A3(
        alu_io_in1[50]), .A4(alu_n120), .Y(alu_n219) );
  NAND2X0_LVT alu_U430 ( .A1(alu_n234), .A2(alu_n218), .Y(alu_shin_14_) );
  AOI22X1_LVT alu_U429 ( .A1(alu_io_in1[14]), .A2(alu_n121), .A3(
        alu_io_in1[49]), .A4(alu_n232), .Y(alu_n218) );
  NAND2X0_LVT alu_U428 ( .A1(alu_n234), .A2(alu_n217), .Y(alu_shin_15_) );
  AOI22X1_LVT alu_U427 ( .A1(alu_io_in1[15]), .A2(alu_n121), .A3(
        alu_io_in1[48]), .A4(alu_n120), .Y(alu_n217) );
  NAND2X0_LVT alu_U426 ( .A1(alu_n234), .A2(alu_n216), .Y(alu_shin_16_) );
  AOI22X1_LVT alu_U425 ( .A1(alu_io_in1[16]), .A2(alu_n121), .A3(
        alu_io_in1[47]), .A4(alu_n232), .Y(alu_n216) );
  NAND2X0_LVT alu_U424 ( .A1(alu_n234), .A2(alu_n215), .Y(alu_shin_17_) );
  AOI22X1_LVT alu_U423 ( .A1(alu_io_in1[17]), .A2(alu_n121), .A3(
        alu_io_in1[46]), .A4(alu_n232), .Y(alu_n215) );
  NAND2X0_LVT alu_U422 ( .A1(alu_n234), .A2(alu_n214), .Y(alu_shin_18_) );
  AOI22X1_LVT alu_U421 ( .A1(alu_io_in1[18]), .A2(alu_n121), .A3(
        alu_io_in1[45]), .A4(alu_n120), .Y(alu_n214) );
  NAND2X0_LVT alu_U420 ( .A1(alu_n234), .A2(alu_n213), .Y(alu_shin_19_) );
  AOI22X1_LVT alu_U419 ( .A1(alu_io_in1[19]), .A2(alu_n121), .A3(
        alu_io_in1[44]), .A4(alu_n232), .Y(alu_n213) );
  NAND2X0_LVT alu_U418 ( .A1(alu_n234), .A2(alu_n212), .Y(alu_shin_20_) );
  AOI22X1_LVT alu_U417 ( .A1(alu_io_in1[20]), .A2(alu_n121), .A3(
        alu_io_in1[43]), .A4(alu_n120), .Y(alu_n212) );
  NAND2X0_LVT alu_U416 ( .A1(alu_n234), .A2(alu_n211), .Y(alu_shin_21_) );
  AOI22X1_LVT alu_U415 ( .A1(alu_io_in1[21]), .A2(alu_n121), .A3(
        alu_io_in1[42]), .A4(alu_n232), .Y(alu_n211) );
  NAND2X0_LVT alu_U414 ( .A1(alu_n234), .A2(alu_n210), .Y(alu_shin_22_) );
  AOI22X1_LVT alu_U413 ( .A1(alu_io_in1[22]), .A2(alu_n121), .A3(
        alu_io_in1[41]), .A4(alu_n232), .Y(alu_n210) );
  NAND2X0_LVT alu_U412 ( .A1(alu_n234), .A2(alu_n209), .Y(alu_shin_23_) );
  AOI22X1_LVT alu_U411 ( .A1(alu_io_in1[23]), .A2(alu_n121), .A3(
        alu_io_in1[40]), .A4(alu_n232), .Y(alu_n209) );
  NAND2X0_LVT alu_U410 ( .A1(alu_n234), .A2(alu_n208), .Y(alu_shin_24_) );
  AOI22X1_LVT alu_U409 ( .A1(alu_io_in1[24]), .A2(alu_n121), .A3(
        alu_io_in1[39]), .A4(alu_n120), .Y(alu_n208) );
  NAND2X0_LVT alu_U408 ( .A1(alu_n234), .A2(alu_n207), .Y(alu_shin_25_) );
  AOI22X1_LVT alu_U407 ( .A1(alu_io_in1[38]), .A2(alu_n120), .A3(alu_n121), 
        .A4(alu_io_in1[25]), .Y(alu_n207) );
  NAND2X0_LVT alu_U406 ( .A1(alu_n234), .A2(alu_n206), .Y(alu_shin_26_) );
  AOI22X1_LVT alu_U405 ( .A1(alu_io_in1[37]), .A2(alu_n120), .A3(alu_n121), 
        .A4(alu_io_in1[26]), .Y(alu_n206) );
  NAND2X0_LVT alu_U404 ( .A1(alu_n234), .A2(alu_n205), .Y(alu_shin_27_) );
  AOI22X1_LVT alu_U403 ( .A1(alu_io_in1[36]), .A2(alu_n120), .A3(alu_n121), 
        .A4(alu_io_in1[27]), .Y(alu_n205) );
  NAND2X0_LVT alu_U402 ( .A1(alu_n234), .A2(alu_n204), .Y(alu_shin_28_) );
  AOI22X1_LVT alu_U401 ( .A1(alu_io_in1[35]), .A2(alu_n120), .A3(alu_n121), 
        .A4(alu_io_in1[28]), .Y(alu_n204) );
  NAND2X0_LVT alu_U400 ( .A1(alu_n234), .A2(alu_n203), .Y(alu_shin_29_) );
  AOI22X1_LVT alu_U399 ( .A1(alu_io_in1[34]), .A2(alu_n120), .A3(alu_n121), 
        .A4(alu_io_in1[29]), .Y(alu_n203) );
  NAND2X0_LVT alu_U398 ( .A1(alu_n234), .A2(alu_n202), .Y(alu_shin_30_) );
  AOI22X1_LVT alu_U397 ( .A1(alu_io_in1[30]), .A2(alu_n121), .A3(
        alu_io_in1[33]), .A4(alu_n120), .Y(alu_n202) );
  NAND2X0_LVT alu_U396 ( .A1(alu_n234), .A2(alu_n201), .Y(alu_shin_31_) );
  AOI22X1_LVT alu_U395 ( .A1(alu_io_in1[32]), .A2(alu_n120), .A3(alu_n121), 
        .A4(alu_io_in1[31]), .Y(alu_n201) );
  NOR2X0_LVT alu_U394 ( .A1(alu_n440), .A2(alu_n121), .Y(alu_n232) );
  NAND2X0_LVT alu_U393 ( .A1(alu_n119), .A2(alu_n198), .Y(alu_shin_32_) );
  AOI22X1_LVT alu_U392 ( .A1(alu_io_in1[32]), .A2(alu_n124), .A3(
        alu_io_in1[31]), .A4(alu_n116), .Y(alu_n198) );
  NAND2X0_LVT alu_U391 ( .A1(alu_n119), .A2(alu_n197), .Y(alu_shin_33_) );
  AOI22X1_LVT alu_U390 ( .A1(alu_io_in1[33]), .A2(alu_n124), .A3(
        alu_io_in1[30]), .A4(alu_n116), .Y(alu_n197) );
  NAND2X0_LVT alu_U389 ( .A1(alu_n119), .A2(alu_n196), .Y(alu_shin_34_) );
  AOI22X1_LVT alu_U388 ( .A1(alu_io_in1[34]), .A2(alu_n124), .A3(
        alu_io_in1[29]), .A4(alu_n116), .Y(alu_n196) );
  NAND2X0_LVT alu_U387 ( .A1(alu_n119), .A2(alu_n195), .Y(alu_shin_35_) );
  AOI22X1_LVT alu_U386 ( .A1(alu_io_in1[35]), .A2(alu_n124), .A3(
        alu_io_in1[28]), .A4(alu_n116), .Y(alu_n195) );
  NAND2X0_LVT alu_U385 ( .A1(alu_n119), .A2(alu_n194), .Y(alu_shin_36_) );
  AOI22X1_LVT alu_U384 ( .A1(alu_io_in1[36]), .A2(alu_n124), .A3(
        alu_io_in1[27]), .A4(alu_n116), .Y(alu_n194) );
  NAND2X0_LVT alu_U383 ( .A1(alu_n119), .A2(alu_n193), .Y(alu_shin_37_) );
  AOI22X1_LVT alu_U382 ( .A1(alu_io_in1[37]), .A2(alu_n124), .A3(
        alu_io_in1[26]), .A4(alu_n116), .Y(alu_n193) );
  NAND2X0_LVT alu_U381 ( .A1(alu_n119), .A2(alu_n192), .Y(alu_shin_38_) );
  AOI22X1_LVT alu_U380 ( .A1(alu_io_in1[38]), .A2(alu_n124), .A3(
        alu_io_in1[25]), .A4(alu_n116), .Y(alu_n192) );
  NAND2X0_LVT alu_U379 ( .A1(alu_n119), .A2(alu_n191), .Y(alu_shin_39_) );
  AOI22X1_LVT alu_U378 ( .A1(alu_io_in1[24]), .A2(alu_n116), .A3(
        alu_io_in1[39]), .A4(alu_n124), .Y(alu_n191) );
  NAND2X0_LVT alu_U377 ( .A1(alu_n119), .A2(alu_n190), .Y(alu_shin_40_) );
  AOI22X1_LVT alu_U376 ( .A1(alu_io_in1[23]), .A2(alu_n116), .A3(
        alu_io_in1[40]), .A4(alu_n124), .Y(alu_n190) );
  NAND2X0_LVT alu_U375 ( .A1(alu_n119), .A2(alu_n189), .Y(alu_shin_41_) );
  AOI22X1_LVT alu_U374 ( .A1(alu_io_in1[22]), .A2(alu_n116), .A3(
        alu_io_in1[41]), .A4(alu_n124), .Y(alu_n189) );
  NAND2X0_LVT alu_U373 ( .A1(alu_n119), .A2(alu_n188), .Y(alu_shin_42_) );
  AOI22X1_LVT alu_U372 ( .A1(alu_io_in1[21]), .A2(alu_n116), .A3(
        alu_io_in1[42]), .A4(alu_n124), .Y(alu_n188) );
  NAND2X0_LVT alu_U371 ( .A1(alu_n119), .A2(alu_n187), .Y(alu_shin_43_) );
  AOI22X1_LVT alu_U370 ( .A1(alu_io_in1[20]), .A2(alu_n116), .A3(
        alu_io_in1[43]), .A4(alu_n124), .Y(alu_n187) );
  NAND2X0_LVT alu_U369 ( .A1(alu_n199), .A2(alu_n186), .Y(alu_shin_44_) );
  AOI22X1_LVT alu_U368 ( .A1(alu_io_in1[19]), .A2(alu_n116), .A3(
        alu_io_in1[44]), .A4(alu_n124), .Y(alu_n186) );
  NAND2X0_LVT alu_U367 ( .A1(alu_n199), .A2(alu_n185), .Y(alu_shin_45_) );
  AOI22X1_LVT alu_U366 ( .A1(alu_io_in1[18]), .A2(alu_n116), .A3(
        alu_io_in1[45]), .A4(alu_n124), .Y(alu_n185) );
  NAND2X0_LVT alu_U365 ( .A1(alu_n199), .A2(alu_n184), .Y(alu_shin_46_) );
  AOI22X1_LVT alu_U364 ( .A1(alu_io_in1[17]), .A2(alu_n116), .A3(
        alu_io_in1[46]), .A4(alu_n124), .Y(alu_n184) );
  NAND2X0_LVT alu_U363 ( .A1(alu_n199), .A2(alu_n183), .Y(alu_shin_47_) );
  AOI22X1_LVT alu_U362 ( .A1(alu_io_in1[16]), .A2(alu_n116), .A3(
        alu_io_in1[47]), .A4(alu_n124), .Y(alu_n183) );
  NAND2X0_LVT alu_U361 ( .A1(alu_n199), .A2(alu_n182), .Y(alu_shin_48_) );
  AOI22X1_LVT alu_U360 ( .A1(alu_io_in1[15]), .A2(alu_n116), .A3(
        alu_io_in1[48]), .A4(alu_n124), .Y(alu_n182) );
  NAND2X0_LVT alu_U359 ( .A1(alu_n199), .A2(alu_n181), .Y(alu_shin_49_) );
  AOI22X1_LVT alu_U358 ( .A1(alu_io_in1[14]), .A2(alu_n116), .A3(
        alu_io_in1[49]), .A4(alu_n124), .Y(alu_n181) );
  NAND2X0_LVT alu_U357 ( .A1(alu_n199), .A2(alu_n180), .Y(alu_shin_50_) );
  AOI22X1_LVT alu_U356 ( .A1(alu_io_in1[13]), .A2(alu_n116), .A3(
        alu_io_in1[50]), .A4(alu_n124), .Y(alu_n180) );
  NAND2X0_LVT alu_U355 ( .A1(alu_n199), .A2(alu_n179), .Y(alu_shin_51_) );
  AOI22X1_LVT alu_U354 ( .A1(alu_io_in1[12]), .A2(alu_n116), .A3(
        alu_io_in1[51]), .A4(alu_n124), .Y(alu_n179) );
  NAND2X0_LVT alu_U353 ( .A1(alu_n199), .A2(alu_n178), .Y(alu_shin_52_) );
  AOI22X1_LVT alu_U352 ( .A1(alu_io_in1[11]), .A2(alu_n116), .A3(
        alu_io_in1[52]), .A4(alu_n124), .Y(alu_n178) );
  NAND2X0_LVT alu_U351 ( .A1(alu_n199), .A2(alu_n177), .Y(alu_shin_53_) );
  AOI22X1_LVT alu_U350 ( .A1(alu_io_in1[10]), .A2(alu_n116), .A3(
        alu_io_in1[53]), .A4(alu_n124), .Y(alu_n177) );
  NAND2X0_LVT alu_U349 ( .A1(alu_n199), .A2(alu_n176), .Y(alu_shin_54_) );
  AOI22X1_LVT alu_U348 ( .A1(alu_io_in1[9]), .A2(alu_n116), .A3(alu_io_in1[54]), .A4(alu_n124), .Y(alu_n176) );
  NAND2X0_LVT alu_U347 ( .A1(alu_n199), .A2(alu_n175), .Y(alu_shin_55_) );
  AOI22X1_LVT alu_U346 ( .A1(alu_io_in1[8]), .A2(alu_n116), .A3(alu_io_in1[55]), .A4(alu_n124), .Y(alu_n175) );
  NAND2X0_LVT alu_U345 ( .A1(alu_n119), .A2(alu_n174), .Y(alu_shin_56_) );
  AOI22X1_LVT alu_U344 ( .A1(alu_io_in1[7]), .A2(alu_n116), .A3(alu_io_in1[56]), .A4(alu_n124), .Y(alu_n174) );
  NAND2X0_LVT alu_U343 ( .A1(alu_n199), .A2(alu_n173), .Y(alu_shin_57_) );
  AOI22X1_LVT alu_U342 ( .A1(alu_io_in1[6]), .A2(alu_n116), .A3(alu_io_in1[57]), .A4(alu_n124), .Y(alu_n173) );
  NAND2X0_LVT alu_U341 ( .A1(alu_n119), .A2(alu_n172), .Y(alu_shin_58_) );
  AOI22X1_LVT alu_U340 ( .A1(alu_io_in1[5]), .A2(alu_n116), .A3(alu_io_in1[58]), .A4(alu_n124), .Y(alu_n172) );
  NAND2X0_LVT alu_U339 ( .A1(alu_n119), .A2(alu_n171), .Y(alu_shin_59_) );
  AOI22X1_LVT alu_U338 ( .A1(alu_io_in1[4]), .A2(alu_n116), .A3(alu_io_in1[59]), .A4(alu_n124), .Y(alu_n171) );
  NAND2X0_LVT alu_U337 ( .A1(alu_n119), .A2(alu_n170), .Y(alu_shin_60_) );
  AOI22X1_LVT alu_U336 ( .A1(alu_io_in1[3]), .A2(alu_n116), .A3(alu_io_in1[60]), .A4(alu_n124), .Y(alu_n170) );
  NAND2X0_LVT alu_U335 ( .A1(alu_n119), .A2(alu_n169), .Y(alu_shin_61_) );
  AOI22X1_LVT alu_U334 ( .A1(alu_io_in1[2]), .A2(alu_n116), .A3(alu_io_in1[61]), .A4(alu_n124), .Y(alu_n169) );
  NAND2X0_LVT alu_U333 ( .A1(alu_n199), .A2(alu_n168), .Y(alu_shin_62_) );
  AOI22X1_LVT alu_U332 ( .A1(alu_io_in1[1]), .A2(alu_n116), .A3(alu_io_in1[62]), .A4(alu_n124), .Y(alu_n168) );
  NAND2X0_LVT alu_U331 ( .A1(alu_n167), .A2(alu_n199), .Y(alu_shin_63_) );
  NAND2X0_LVT alu_U330 ( .A1(alu_io_in1[31]), .A2(alu_n166), .Y(alu_n200) );
  AND2X1_LVT alu_U329 ( .A1(alu_n440), .A2(alu_n125), .Y(alu_n166) );
  INVX1_LVT alu_U328 ( .A(alu_io_dw), .Y(alu_n440) );
  AOI22X1_LVT alu_U327 ( .A1(alu_io_in1[0]), .A2(alu_n116), .A3(alu_io_in1[63]), .A4(alu_n124), .Y(alu_n167) );
  NAND2X0_LVT alu_U326 ( .A1(alu_io_fn[1]), .A2(alu_n126), .Y(alu_n243) );
  MUX21X1_LVT alu_U325 ( .A1(alu_io_fn[1]), .A2(alu_n126), .S0(alu_io_fn[2]), 
        .Y(alu_n165) );
  NAND2X0_LVT alu_U324 ( .A1(alu_n235), .A2(alu_n163), .Y(alu_n164) );
  NAND4X0_LVT alu_U323 ( .A1(alu_n162), .A2(alu_n161), .A3(alu_n160), .A4(
        alu_n159), .Y(alu_n163) );
  NOR4X1_LVT alu_U322 ( .A1(alu_n158), .A2(alu_n157), .A3(alu_n156), .A4(
        alu_n155), .Y(alu_n159) );
  NAND4X0_LVT alu_U321 ( .A1(alu_n368), .A2(alu_n350), .A3(alu_n338), .A4(
        alu_n344), .Y(alu_n155) );
  NAND4X0_LVT alu_U320 ( .A1(alu_n392), .A2(alu_n374), .A3(alu_n380), .A4(
        alu_n362), .Y(alu_n156) );
  NAND4X0_LVT alu_U319 ( .A1(alu_n416), .A2(alu_n398), .A3(alu_n404), .A4(
        alu_n386), .Y(alu_n157) );
  NAND4X0_LVT alu_U318 ( .A1(alu_n307), .A2(alu_n313), .A3(alu_n410), .A4(
        alu_n294), .Y(alu_n158) );
  NOR4X1_LVT alu_U317 ( .A1(alu_n149), .A2(alu_n148), .A3(alu_n147), .A4(
        alu_n146), .Y(alu_n160) );
  NAND4X0_LVT alu_U316 ( .A1(alu_n326), .A2(alu_n331), .A3(alu_n319), .A4(
        alu_n324), .Y(alu_n146) );
  NAND4X0_LVT alu_U315 ( .A1(alu_n453), .A2(alu_n452), .A3(alu_n446), .A4(
        alu_n437), .Y(alu_n147) );
  NAND4X0_LVT alu_U314 ( .A1(alu_n457), .A2(alu_n456), .A3(alu_n455), .A4(
        alu_n454), .Y(alu_n148) );
  NAND4X0_LVT alu_U313 ( .A1(alu_n588), .A2(alu_n568), .A3(alu_n544), .A4(
        alu_n495), .Y(alu_n149) );
  NOR4X1_LVT alu_U312 ( .A1(alu_n145), .A2(alu_n144), .A3(alu_n143), .A4(
        alu_n142), .Y(alu_n161) );
  NAND4X0_LVT alu_U311 ( .A1(alu_n477), .A2(alu_n471), .A3(alu_n465), .A4(
        alu_n459), .Y(alu_n142) );
  NAND4X0_LVT alu_U310 ( .A1(alu_n508), .A2(alu_n501), .A3(alu_n489), .A4(
        alu_n483), .Y(alu_n143) );
  NAND4X0_LVT alu_U309 ( .A1(alu_n532), .A2(alu_n526), .A3(alu_n520), .A4(
        alu_n514), .Y(alu_n144) );
  NAND4X0_LVT alu_U308 ( .A1(alu_n562), .A2(alu_n556), .A3(alu_n538), .A4(
        alu_n550), .Y(alu_n145) );
  NOR4X1_LVT alu_U307 ( .A1(alu_n257), .A2(alu_n251), .A3(alu_n141), .A4(
        alu_n140), .Y(alu_n162) );
  NAND4X0_LVT alu_U306 ( .A1(alu_n139), .A2(alu_n138), .A3(alu_n356), .A4(
        alu_n422), .Y(alu_n140) );
  NOR4X1_LVT alu_U305 ( .A1(alu_n137), .A2(alu_n594), .A3(alu_n580), .A4(
        alu_n573), .Y(alu_n138) );
  NAND2X0_LVT alu_U304 ( .A1(alu_n136), .A2(alu_n126), .Y(alu_n137) );
  AND4X1_LVT alu_U303 ( .A1(alu_n240), .A2(alu_n264), .A3(alu_n270), .A4(
        alu_n282), .Y(alu_n139) );
  NAND4X0_LVT alu_U302 ( .A1(alu_n131), .A2(alu_n604), .A3(alu_n288), .A4(
        alu_n276), .Y(alu_n141) );
  NAND2X0_LVT alu_U301 ( .A1(alu_n129), .A2(alu_n125), .Y(alu_n235) );
  MUX21X1_LVT alu_U300 ( .A1(alu_n128), .A2(alu_n127), .S0(alu_io_in1[63]), 
        .Y(alu_n129) );
  MUX21X1_LVT alu_U299 ( .A1(alu_n241), .A2(alu_n607), .S0(alu_io_in2[63]), 
        .Y(alu_n127) );
  INVX1_LVT alu_U298 ( .A(alu_io_fn[1]), .Y(alu_n241) );
  MUX21X1_LVT alu_U297 ( .A1(alu_n607), .A2(alu_io_fn[1]), .S0(alu_io_in2[63]), 
        .Y(alu_n128) );
  NAND2X0_LVT alu_U296 ( .A1(alu_n238), .A2(alu_io_fn[2]), .Y(alu_n118) );
  NAND2X0_LVT alu_U295 ( .A1(alu_io_dw), .A2(alu_n121), .Y(alu_n117) );
  NBUFFX2_LVT alu_U294 ( .A(alu_n232), .Y(alu_n120) );
  NBUFFX2_LVT alu_U293 ( .A(alu_n199), .Y(alu_n119) );
  XOR2X1_LVT alu_U292 ( .A1(alu_io_in2[9]), .A2(alu_io_fn[3]), .Y(
        alu_in2_inv_9_) );
  XOR2X1_LVT alu_U291 ( .A1(alu_io_in2[7]), .A2(alu_io_fn[3]), .Y(
        alu_in2_inv_7_) );
  XOR2X1_LVT alu_U290 ( .A1(alu_io_in2[3]), .A2(alu_io_fn[3]), .Y(
        alu_in2_inv_3_) );
  INVX1_LVT alu_U289 ( .A(alu_n117), .Y(alu_n124) );
  XNOR2X1_LVT alu_U288 ( .A1(alu_in2_inv_46_), .A2(alu_io_in1[46]), .Y(
        alu_n495) );
  XNOR2X1_LVT alu_U287 ( .A1(alu_in2_inv_54_), .A2(alu_io_in1[54]), .Y(
        alu_n544) );
  XNOR2X1_LVT alu_U286 ( .A1(alu_in2_inv_55_), .A2(alu_io_in1[55]), .Y(
        alu_n550) );
  XNOR2X1_LVT alu_U285 ( .A1(alu_in2_inv_58_), .A2(alu_io_in1[58]), .Y(
        alu_n568) );
  XOR2X1_LVT alu_U284 ( .A1(alu_in2_inv_62_), .A2(alu_io_in1[62]), .Y(alu_n594) );
  XOR2X1_LVT alu_U283 ( .A1(alu_in2_inv_60_), .A2(alu_io_in1[60]), .Y(alu_n580) );
  XOR2X1_LVT alu_U282 ( .A1(alu_in2_inv_59_), .A2(alu_io_in1[59]), .Y(alu_n573) );
  XOR2X1_LVT alu_U281 ( .A1(alu_in2_inv_2_), .A2(alu_io_in1[2]), .Y(alu_n257)
         );
  XOR2X1_LVT alu_U280 ( .A1(alu_in2_inv_1_), .A2(alu_io_in1[1]), .Y(alu_n251)
         );
  XOR2X1_LVT alu_U279 ( .A1(alu_in2_inv_5_), .A2(alu_n130), .Y(alu_n276) );
  XOR2X1_LVT alu_U278 ( .A1(alu_in2_inv_0_), .A2(alu_n132), .Y(alu_n240) );
  XOR2X1_LVT alu_U277 ( .A1(alu_in2_inv_3_), .A2(alu_n133), .Y(alu_n264) );
  XOR2X1_LVT alu_U276 ( .A1(alu_in2_inv_4_), .A2(alu_n134), .Y(alu_n270) );
  XOR2X1_LVT alu_U275 ( .A1(alu_io_in2[9]), .A2(alu_n135), .Y(alu_n136) );
  XNOR2X1_LVT alu_U274 ( .A1(alu_in2_inv_11_), .A2(alu_io_in1[11]), .Y(
        alu_n313) );
  XNOR2X1_LVT alu_U273 ( .A1(alu_in2_inv_28_), .A2(alu_io_in1[28]), .Y(
        alu_n410) );
  XNOR2X1_LVT alu_U272 ( .A1(alu_in2_inv_8_), .A2(alu_io_in1[8]), .Y(alu_n294)
         );
  XOR2X1_LVT alu_U271 ( .A1(alu_in2_inv_24_), .A2(alu_n150), .Y(alu_n386) );
  XOR2X1_LVT alu_U270 ( .A1(alu_in2_inv_22_), .A2(alu_n151), .Y(alu_n374) );
  XOR2X1_LVT alu_U269 ( .A1(alu_in2_inv_23_), .A2(alu_n152), .Y(alu_n380) );
  XOR2X1_LVT alu_U268 ( .A1(alu_in2_inv_20_), .A2(alu_n153), .Y(alu_n362) );
  XOR2X1_LVT alu_U267 ( .A1(alu_in2_inv_21_), .A2(alu_n154), .Y(alu_n368) );
  XOR2X1_LVT alu_U266 ( .A1(alu_n164), .A2(alu_io_fn[0]), .Y(alu_io_cmp_out)
         );
  NAND2X0_LVT alu_U265 ( .A1(alu_n125), .A2(alu_n241), .Y(alu_n242) );
  AND2X1_LVT alu_U264 ( .A1(alu_io_dw), .A2(alu_io_in2[5]), .Y(alu_shamt_5_)
         );
  INVX1_LVT alu_U263 ( .A(alu_n126), .Y(alu_n125) );
  AND3X1_LVT alu_U262 ( .A1(alu_n244), .A2(alu_n243), .A3(alu_n242), .Y(
        alu_n434) );
  AND2X1_LVT alu_U261 ( .A1(alu_io_dw), .A2(alu_n434), .Y(alu_n602) );
  NAND3X0_LVT alu_U260 ( .A1(alu_n165), .A2(alu_io_fn[0]), .A3(alu_n243), .Y(
        alu_n116) );
  INVX1_LVT alu_U259 ( .A(alu_n116), .Y(alu_n121) );
  INVX1_LVT alu_U258 ( .A(alu_n118), .Y(alu_n122) );
  INVX1_LVT alu_U257 ( .A(alu_n593), .Y(alu_n605) );
  AND2X1_LVT alu_U256 ( .A1(alu_n122), .A2(alu_io_dw), .Y(alu_n603) );
  AND2X1_LVT alu_U255 ( .A1(alu_n441), .A2(alu_io_dw), .Y(alu_n598) );
  INVX1_LVT alu_U254 ( .A(alu_n435), .Y(alu_n423) );
  XOR2X1_LVT alu_U253 ( .A1(alu_io_in2[5]), .A2(alu_io_fn[3]), .Y(
        alu_in2_inv_5_) );
  NOR2X1_LVT alu_U252 ( .A1(alu_io_fn[0]), .A2(alu_io_fn[2]), .Y(alu_n244) );
  XOR2X1_LVT alu_U251 ( .A1(alu_io_in2[36]), .A2(alu_n125), .Y(alu_in2_inv_36_) );
  XOR2X1_LVT alu_U250 ( .A1(alu_io_in2[37]), .A2(alu_n125), .Y(alu_in2_inv_37_) );
  XOR2X1_LVT alu_U249 ( .A1(alu_io_in2[40]), .A2(alu_n125), .Y(alu_in2_inv_40_) );
  XOR2X1_LVT alu_U248 ( .A1(alu_io_in2[34]), .A2(alu_n125), .Y(alu_in2_inv_34_) );
  XOR2X1_LVT alu_U247 ( .A1(alu_io_in2[42]), .A2(alu_n125), .Y(alu_in2_inv_42_) );
  XOR2X1_LVT alu_U246 ( .A1(alu_io_in2[33]), .A2(alu_n125), .Y(alu_in2_inv_33_) );
  XOR2X1_LVT alu_U245 ( .A1(alu_io_in2[31]), .A2(alu_n125), .Y(alu_in2_inv_31_) );
  XOR2X1_LVT alu_U244 ( .A1(alu_io_in2[41]), .A2(alu_n125), .Y(alu_in2_inv_41_) );
  XOR2X1_LVT alu_U243 ( .A1(alu_io_in2[32]), .A2(alu_n125), .Y(alu_in2_inv_32_) );
  XOR2X1_LVT alu_U242 ( .A1(alu_io_in2[35]), .A2(alu_n125), .Y(alu_in2_inv_35_) );
  XOR2X1_LVT alu_U241 ( .A1(alu_io_in2[4]), .A2(alu_n125), .Y(alu_in2_inv_4_)
         );
  XOR2X1_LVT alu_U240 ( .A1(alu_io_in2[60]), .A2(alu_n125), .Y(alu_in2_inv_60_) );
  XOR2X1_LVT alu_U239 ( .A1(alu_io_in2[50]), .A2(alu_n125), .Y(alu_in2_inv_50_) );
  XOR2X1_LVT alu_U238 ( .A1(alu_io_in2[59]), .A2(alu_n125), .Y(alu_in2_inv_59_) );
  XOR2X1_LVT alu_U237 ( .A1(alu_io_in2[49]), .A2(alu_n125), .Y(alu_in2_inv_49_) );
  XOR2X1_LVT alu_U236 ( .A1(alu_io_in2[62]), .A2(alu_n125), .Y(alu_in2_inv_62_) );
  XOR2X1_LVT alu_U235 ( .A1(alu_io_in2[47]), .A2(alu_n125), .Y(alu_in2_inv_47_) );
  XOR2X1_LVT alu_U234 ( .A1(alu_io_in2[61]), .A2(alu_n125), .Y(alu_in2_inv_61_) );
  XOR2X1_LVT alu_U233 ( .A1(alu_io_in2[56]), .A2(alu_n125), .Y(alu_in2_inv_56_) );
  XOR2X1_LVT alu_U232 ( .A1(alu_io_in2[48]), .A2(alu_n125), .Y(alu_in2_inv_48_) );
  XOR2X1_LVT alu_U231 ( .A1(alu_io_in2[55]), .A2(alu_n125), .Y(alu_in2_inv_55_) );
  XOR2X1_LVT alu_U230 ( .A1(alu_io_in2[0]), .A2(alu_n125), .Y(alu_in2_inv_0_)
         );
  XOR2X1_LVT alu_U229 ( .A1(alu_io_in2[57]), .A2(alu_n125), .Y(alu_in2_inv_57_) );
  XOR2X1_LVT alu_U228 ( .A1(alu_io_in2[58]), .A2(alu_n125), .Y(alu_in2_inv_58_) );
  XOR2X1_LVT alu_U227 ( .A1(alu_io_in2[39]), .A2(alu_n125), .Y(alu_in2_inv_39_) );
  XOR2X1_LVT alu_U226 ( .A1(alu_io_in2[38]), .A2(alu_n125), .Y(alu_in2_inv_38_) );
  XOR2X1_LVT alu_U225 ( .A1(alu_io_in2[8]), .A2(alu_n125), .Y(alu_in2_inv_8_)
         );
  XOR2X1_LVT alu_U224 ( .A1(alu_io_in2[54]), .A2(alu_n125), .Y(alu_in2_inv_54_) );
  XOR2X1_LVT alu_U223 ( .A1(alu_io_in2[52]), .A2(alu_n125), .Y(alu_in2_inv_52_) );
  XOR2X1_LVT alu_U222 ( .A1(alu_io_in2[53]), .A2(alu_n125), .Y(alu_in2_inv_53_) );
  XOR2X1_LVT alu_U221 ( .A1(alu_io_in2[46]), .A2(alu_n125), .Y(alu_in2_inv_46_) );
  XOR2X1_LVT alu_U220 ( .A1(alu_io_in2[45]), .A2(alu_n125), .Y(alu_in2_inv_45_) );
  XOR2X1_LVT alu_U219 ( .A1(alu_io_in2[43]), .A2(alu_n125), .Y(alu_in2_inv_43_) );
  XOR2X1_LVT alu_U218 ( .A1(alu_io_in2[44]), .A2(alu_n125), .Y(alu_in2_inv_44_) );
  XOR2X1_LVT alu_U217 ( .A1(alu_io_in2[6]), .A2(alu_n125), .Y(alu_in2_inv_6_)
         );
  XOR2X1_LVT alu_U216 ( .A1(alu_io_in2[10]), .A2(alu_n125), .Y(alu_in2_inv_10_) );
  XOR2X1_LVT alu_U215 ( .A1(alu_io_in2[63]), .A2(alu_n125), .Y(alu_in2_inv_63_) );
  XOR2X1_LVT alu_U214 ( .A1(alu_io_in2[51]), .A2(alu_n125), .Y(alu_in2_inv_51_) );
  XOR2X1_LVT alu_U213 ( .A1(alu_io_in2[13]), .A2(alu_n125), .Y(alu_in2_inv_13_) );
  XOR2X1_LVT alu_U212 ( .A1(alu_io_in2[22]), .A2(alu_n125), .Y(alu_in2_inv_22_) );
  XOR2X1_LVT alu_U211 ( .A1(alu_io_in2[21]), .A2(alu_n125), .Y(alu_in2_inv_21_) );
  XOR2X1_LVT alu_U210 ( .A1(alu_io_in2[12]), .A2(alu_n125), .Y(alu_in2_inv_12_) );
  XOR2X1_LVT alu_U209 ( .A1(alu_io_in2[27]), .A2(alu_n125), .Y(alu_in2_inv_27_) );
  XOR2X1_LVT alu_U208 ( .A1(alu_io_in2[28]), .A2(alu_n125), .Y(alu_in2_inv_28_) );
  XOR2X1_LVT alu_U207 ( .A1(alu_io_in2[11]), .A2(alu_n125), .Y(alu_in2_inv_11_) );
  XOR2X1_LVT alu_U206 ( .A1(alu_io_in2[2]), .A2(alu_n125), .Y(alu_in2_inv_2_)
         );
  XOR2X1_LVT alu_U205 ( .A1(alu_io_in2[1]), .A2(alu_n125), .Y(alu_in2_inv_1_)
         );
  XOR2X1_LVT alu_U204 ( .A1(alu_io_in2[26]), .A2(alu_n125), .Y(alu_in2_inv_26_) );
  XOR2X1_LVT alu_U203 ( .A1(alu_io_in2[24]), .A2(alu_n125), .Y(alu_in2_inv_24_) );
  XOR2X1_LVT alu_U202 ( .A1(alu_io_in2[23]), .A2(alu_n125), .Y(alu_in2_inv_23_) );
  XOR2X1_LVT alu_U201 ( .A1(alu_io_in2[20]), .A2(alu_n125), .Y(alu_in2_inv_20_) );
  XOR2X1_LVT alu_U200 ( .A1(alu_io_in2[19]), .A2(alu_n125), .Y(alu_in2_inv_19_) );
  XOR2X1_LVT alu_U199 ( .A1(alu_io_in2[25]), .A2(alu_n125), .Y(alu_in2_inv_25_) );
  XOR2X1_LVT alu_U198 ( .A1(alu_io_in2[18]), .A2(alu_n125), .Y(alu_in2_inv_18_) );
  XOR2X1_LVT alu_U197 ( .A1(alu_io_in2[30]), .A2(alu_io_fn[3]), .Y(
        alu_in2_inv_30_) );
  XOR2X1_LVT alu_U196 ( .A1(alu_io_in2[29]), .A2(alu_n125), .Y(alu_in2_inv_29_) );
  XOR2X1_LVT alu_U195 ( .A1(alu_io_in2[15]), .A2(alu_n125), .Y(alu_in2_inv_15_) );
  XOR2X1_LVT alu_U194 ( .A1(alu_io_in2[17]), .A2(alu_n125), .Y(alu_in2_inv_17_) );
  XOR2X1_LVT alu_U193 ( .A1(alu_io_in2[14]), .A2(alu_n125), .Y(alu_in2_inv_14_) );
  XOR2X1_LVT alu_U192 ( .A1(alu_io_in2[16]), .A2(alu_io_fn[3]), .Y(
        alu_in2_inv_16_) );
  XOR2X1_LVT alu_U191 ( .A1(alu_in2_inv_31_), .A2(alu_io_in1[31]), .Y(alu_n428) );
  INVX0_LVT alu_U190 ( .A(alu_n428), .Y(alu_n131) );
  INVX0_LVT alu_U189 ( .A(alu_n_T_101_16_), .Y(alu_n503) );
  INVX0_LVT alu_U188 ( .A(alu_n_T_101_32_), .Y(alu_n439) );
  INVX0_LVT alu_U187 ( .A(alu_n_T_101_30_), .Y(alu_n448) );
  NBUFFX2_LVT alu_U186 ( .A(alu_n606), .Y(alu_n115) );
  INVX0_LVT alu_U185 ( .A(alu_n235), .Y(alu_n250) );
  INVX1_LVT alu_U184 ( .A(alu_io_fn[3]), .Y(alu_n126) );
  INVX1_LVT alu_U183 ( .A(alu_io_fn[2]), .Y(alu_n236) );
  INVX1_LVT alu_U182 ( .A(alu_io_fn[0]), .Y(alu_n237) );
  INVX0_LVT alu_U181 ( .A(alu_n243), .Y(alu_n238) );
  INVX1_LVT alu_U180 ( .A(alu_n598), .Y(alu_n123) );
  INVX1_LVT alu_U179 ( .A(alu_io_in1[0]), .Y(alu_n132) );
  INVX1_LVT alu_U178 ( .A(alu_io_in1[24]), .Y(alu_n150) );
  INVX1_LVT alu_U177 ( .A(alu_io_in1[22]), .Y(alu_n151) );
  INVX1_LVT alu_U176 ( .A(alu_io_in1[23]), .Y(alu_n152) );
  INVX1_LVT alu_U175 ( .A(alu_io_in1[9]), .Y(alu_n135) );
  INVX1_LVT alu_U174 ( .A(alu_io_in1[5]), .Y(alu_n130) );
  INVX1_LVT alu_U173 ( .A(alu_io_in1[21]), .Y(alu_n154) );
  INVX1_LVT alu_U172 ( .A(alu_io_in1[4]), .Y(alu_n134) );
  INVX1_LVT alu_U171 ( .A(alu_io_in1[20]), .Y(alu_n153) );
  INVX1_LVT alu_U170 ( .A(alu_io_in1[3]), .Y(alu_n133) );
  OR2X1_LVT alu_U169 ( .A1(alu_n116), .A2(alu_n200), .Y(alu_n199) );
  INVX1_LVT alu_U168 ( .A(alu_io_in2[9]), .Y(alu_n299) );
  AND2X2_LVT alu_U167 ( .A1(alu_n125), .A2(alu_shin_63_), .Y(alu_n_T_100_64_)
         );
  OR2X4_LVT alu_U166 ( .A1(alu_n121), .A2(alu_n200), .Y(alu_n234) );
  AO22X1_LVT alu_U165 ( .A1(alu_io_in1[57]), .A2(alu_in2_inv_57_), .A3(
        alu_n113), .A4(alu_n114), .Y(alu_n562) );
  INVX0_LVT alu_U164 ( .A(alu_in2_inv_57_), .Y(alu_n114) );
  INVX0_LVT alu_U163 ( .A(alu_io_in1[57]), .Y(alu_n113) );
  AO22X1_LVT alu_U162 ( .A1(alu_io_in1[56]), .A2(alu_in2_inv_56_), .A3(
        alu_n111), .A4(alu_n112), .Y(alu_n556) );
  INVX0_LVT alu_U161 ( .A(alu_in2_inv_56_), .Y(alu_n112) );
  INVX0_LVT alu_U160 ( .A(alu_io_in1[56]), .Y(alu_n111) );
  AO22X1_LVT alu_U159 ( .A1(alu_io_in1[51]), .A2(alu_in2_inv_51_), .A3(
        alu_n109), .A4(alu_n110), .Y(alu_n526) );
  INVX0_LVT alu_U158 ( .A(alu_in2_inv_51_), .Y(alu_n110) );
  INVX0_LVT alu_U157 ( .A(alu_io_in1[51]), .Y(alu_n109) );
  AO22X1_LVT alu_U156 ( .A1(alu_io_in1[50]), .A2(alu_in2_inv_50_), .A3(
        alu_n107), .A4(alu_n108), .Y(alu_n520) );
  INVX0_LVT alu_U155 ( .A(alu_in2_inv_50_), .Y(alu_n108) );
  INVX0_LVT alu_U154 ( .A(alu_io_in1[50]), .Y(alu_n107) );
  AO22X1_LVT alu_U153 ( .A1(alu_io_in1[49]), .A2(alu_in2_inv_49_), .A3(
        alu_n105), .A4(alu_n106), .Y(alu_n514) );
  INVX0_LVT alu_U152 ( .A(alu_in2_inv_49_), .Y(alu_n106) );
  INVX0_LVT alu_U151 ( .A(alu_io_in1[49]), .Y(alu_n105) );
  AO22X1_LVT alu_U150 ( .A1(alu_io_in1[45]), .A2(alu_in2_inv_45_), .A3(
        alu_n103), .A4(alu_n104), .Y(alu_n489) );
  INVX0_LVT alu_U149 ( .A(alu_in2_inv_45_), .Y(alu_n104) );
  INVX0_LVT alu_U148 ( .A(alu_io_in1[45]), .Y(alu_n103) );
  AO22X1_LVT alu_U147 ( .A1(alu_io_in1[44]), .A2(alu_in2_inv_44_), .A3(
        alu_n101), .A4(alu_n102), .Y(alu_n483) );
  INVX0_LVT alu_U146 ( .A(alu_in2_inv_44_), .Y(alu_n102) );
  INVX0_LVT alu_U145 ( .A(alu_io_in1[44]), .Y(alu_n101) );
  AO22X1_LVT alu_U144 ( .A1(alu_io_in1[43]), .A2(alu_in2_inv_43_), .A3(alu_n99), .A4(alu_n100), .Y(alu_n477) );
  INVX0_LVT alu_U143 ( .A(alu_in2_inv_43_), .Y(alu_n100) );
  INVX0_LVT alu_U142 ( .A(alu_io_in1[43]), .Y(alu_n99) );
  AO22X1_LVT alu_U141 ( .A1(alu_io_in1[42]), .A2(alu_in2_inv_42_), .A3(alu_n97), .A4(alu_n98), .Y(alu_n471) );
  INVX0_LVT alu_U140 ( .A(alu_in2_inv_42_), .Y(alu_n98) );
  INVX0_LVT alu_U139 ( .A(alu_io_in1[42]), .Y(alu_n97) );
  AO22X1_LVT alu_U138 ( .A1(alu_io_in1[41]), .A2(alu_in2_inv_41_), .A3(alu_n95), .A4(alu_n96), .Y(alu_n465) );
  INVX0_LVT alu_U137 ( .A(alu_in2_inv_41_), .Y(alu_n96) );
  INVX0_LVT alu_U136 ( .A(alu_io_in1[41]), .Y(alu_n95) );
  AO22X1_LVT alu_U135 ( .A1(alu_io_in1[40]), .A2(alu_in2_inv_40_), .A3(alu_n93), .A4(alu_n94), .Y(alu_n459) );
  INVX0_LVT alu_U134 ( .A(alu_in2_inv_40_), .Y(alu_n94) );
  INVX0_LVT alu_U133 ( .A(alu_io_in1[40]), .Y(alu_n93) );
  AO22X1_LVT alu_U132 ( .A1(alu_io_in1[33]), .A2(alu_in2_inv_33_), .A3(alu_n91), .A4(alu_n92), .Y(alu_n446) );
  INVX0_LVT alu_U131 ( .A(alu_in2_inv_33_), .Y(alu_n92) );
  INVX0_LVT alu_U130 ( .A(alu_io_in1[33]), .Y(alu_n91) );
  AO22X1_LVT alu_U129 ( .A1(alu_io_in1[53]), .A2(alu_in2_inv_53_), .A3(alu_n89), .A4(alu_n90), .Y(alu_n538) );
  INVX0_LVT alu_U128 ( .A(alu_in2_inv_53_), .Y(alu_n90) );
  INVX0_LVT alu_U127 ( .A(alu_io_in1[53]), .Y(alu_n89) );
  AO22X1_LVT alu_U126 ( .A1(alu_io_in1[48]), .A2(alu_in2_inv_48_), .A3(alu_n87), .A4(alu_n88), .Y(alu_n508) );
  INVX0_LVT alu_U125 ( .A(alu_in2_inv_48_), .Y(alu_n88) );
  INVX0_LVT alu_U124 ( .A(alu_io_in1[48]), .Y(alu_n87) );
  AO22X1_LVT alu_U123 ( .A1(alu_io_in1[47]), .A2(alu_in2_inv_47_), .A3(alu_n85), .A4(alu_n86), .Y(alu_n501) );
  INVX0_LVT alu_U122 ( .A(alu_in2_inv_47_), .Y(alu_n86) );
  INVX0_LVT alu_U121 ( .A(alu_io_in1[47]), .Y(alu_n85) );
  AO22X1_LVT alu_U120 ( .A1(alu_io_in1[38]), .A2(alu_in2_inv_38_), .A3(alu_n83), .A4(alu_n84), .Y(alu_n456) );
  INVX0_LVT alu_U119 ( .A(alu_in2_inv_38_), .Y(alu_n84) );
  INVX0_LVT alu_U118 ( .A(alu_io_in1[38]), .Y(alu_n83) );
  AO22X1_LVT alu_U117 ( .A1(alu_io_in1[27]), .A2(alu_in2_inv_27_), .A3(alu_n81), .A4(alu_n82), .Y(alu_n404) );
  INVX0_LVT alu_U116 ( .A(alu_in2_inv_27_), .Y(alu_n82) );
  INVX0_LVT alu_U115 ( .A(alu_io_in1[27]), .Y(alu_n81) );
  AO22X1_LVT alu_U114 ( .A1(alu_io_in1[19]), .A2(alu_in2_inv_19_), .A3(alu_n79), .A4(alu_n80), .Y(alu_n356) );
  INVX0_LVT alu_U113 ( .A(alu_in2_inv_19_), .Y(alu_n80) );
  INVX0_LVT alu_U112 ( .A(alu_io_in1[19]), .Y(alu_n79) );
  AO22X1_LVT alu_U111 ( .A1(alu_io_in1[61]), .A2(alu_in2_inv_61_), .A3(alu_n77), .A4(alu_n78), .Y(alu_n588) );
  INVX0_LVT alu_U110 ( .A(alu_in2_inv_61_), .Y(alu_n78) );
  INVX0_LVT alu_U109 ( .A(alu_io_in1[61]), .Y(alu_n77) );
  AO22X1_LVT alu_U108 ( .A1(alu_io_in1[52]), .A2(alu_in2_inv_52_), .A3(alu_n75), .A4(alu_n76), .Y(alu_n532) );
  INVX0_LVT alu_U107 ( .A(alu_in2_inv_52_), .Y(alu_n76) );
  INVX0_LVT alu_U106 ( .A(alu_io_in1[52]), .Y(alu_n75) );
  AO22X1_LVT alu_U105 ( .A1(alu_io_in1[37]), .A2(alu_in2_inv_37_), .A3(alu_n73), .A4(alu_n74), .Y(alu_n455) );
  INVX0_LVT alu_U104 ( .A(alu_in2_inv_37_), .Y(alu_n74) );
  INVX0_LVT alu_U103 ( .A(alu_io_in1[37]), .Y(alu_n73) );
  AO22X1_LVT alu_U102 ( .A1(alu_io_in1[36]), .A2(alu_in2_inv_36_), .A3(alu_n71), .A4(alu_n72), .Y(alu_n454) );
  INVX0_LVT alu_U101 ( .A(alu_in2_inv_36_), .Y(alu_n72) );
  INVX0_LVT alu_U100 ( .A(alu_io_in1[36]), .Y(alu_n71) );
  AO22X1_LVT alu_U99 ( .A1(alu_io_in1[34]), .A2(alu_in2_inv_34_), .A3(alu_n69), 
        .A4(alu_n70), .Y(alu_n452) );
  INVX0_LVT alu_U98 ( .A(alu_in2_inv_34_), .Y(alu_n70) );
  INVX0_LVT alu_U97 ( .A(alu_io_in1[34]), .Y(alu_n69) );
  AO22X1_LVT alu_U96 ( .A1(alu_io_in1[32]), .A2(alu_in2_inv_32_), .A3(alu_n67), 
        .A4(alu_n68), .Y(alu_n437) );
  INVX0_LVT alu_U95 ( .A(alu_in2_inv_32_), .Y(alu_n68) );
  INVX0_LVT alu_U94 ( .A(alu_io_in1[32]), .Y(alu_n67) );
  AO22X1_LVT alu_U93 ( .A1(alu_io_in1[29]), .A2(alu_in2_inv_29_), .A3(alu_n65), 
        .A4(alu_n66), .Y(alu_n416) );
  INVX0_LVT alu_U92 ( .A(alu_in2_inv_29_), .Y(alu_n66) );
  INVX0_LVT alu_U91 ( .A(alu_io_in1[29]), .Y(alu_n65) );
  AO22X1_LVT alu_U90 ( .A1(alu_io_in1[17]), .A2(alu_in2_inv_17_), .A3(alu_n63), 
        .A4(alu_n64), .Y(alu_n344) );
  INVX0_LVT alu_U89 ( .A(alu_in2_inv_17_), .Y(alu_n64) );
  INVX0_LVT alu_U88 ( .A(alu_io_in1[17]), .Y(alu_n63) );
  NAND4X0_LVT alu_U87 ( .A1(alu_n60), .A2(alu_n115), .A3(alu_n61), .A4(alu_n62), .Y(alu_io_out[63]) );
  NAND3X0_LVT alu_U86 ( .A1(alu_io_in1[63]), .A2(alu_io_in2[63]), .A3(alu_n603), .Y(alu_n62) );
  AOI22X1_LVT alu_U85 ( .A1(alu_n607), .A2(alu_n602), .A3(alu_n124), .A4(
        alu_n_T_101_63_), .Y(alu_n61) );
  OA22X1_LVT alu_U84 ( .A1(alu_n605), .A2(alu_n604), .A3(alu_n123), .A4(
        alu_n59), .Y(alu_n60) );
  INVX0_LVT alu_U83 ( .A(alu_n_T_101_0_), .Y(alu_n59) );
  AO22X1_LVT alu_U82 ( .A1(alu_io_in1[35]), .A2(alu_in2_inv_35_), .A3(alu_n57), 
        .A4(alu_n58), .Y(alu_n453) );
  INVX0_LVT alu_U81 ( .A(alu_in2_inv_35_), .Y(alu_n58) );
  INVX0_LVT alu_U80 ( .A(alu_io_in1[35]), .Y(alu_n57) );
  AO22X1_LVT alu_U79 ( .A1(alu_io_in1[26]), .A2(alu_in2_inv_26_), .A3(alu_n55), 
        .A4(alu_n56), .Y(alu_n398) );
  INVX0_LVT alu_U78 ( .A(alu_in2_inv_26_), .Y(alu_n56) );
  INVX0_LVT alu_U77 ( .A(alu_io_in1[26]), .Y(alu_n55) );
  AO22X1_LVT alu_U76 ( .A1(alu_io_in1[18]), .A2(alu_in2_inv_18_), .A3(alu_n53), 
        .A4(alu_n54), .Y(alu_n350) );
  INVX0_LVT alu_U75 ( .A(alu_in2_inv_18_), .Y(alu_n54) );
  INVX0_LVT alu_U74 ( .A(alu_io_in1[18]), .Y(alu_n53) );
  NAND4X0_LVT alu_U73 ( .A1(alu_n50), .A2(alu_n115), .A3(alu_n51), .A4(alu_n52), .Y(alu_io_out[39]) );
  NAND3X0_LVT alu_U72 ( .A1(alu_io_in1[39]), .A2(alu_io_in2[39]), .A3(alu_n603), .Y(alu_n52) );
  AOI22X1_LVT alu_U71 ( .A1(alu_n602), .A2(alu_io_adder_out_39_), .A3(alu_n124), .A4(alu_n_T_101_39_), .Y(alu_n51) );
  OA22X1_LVT alu_U70 ( .A1(alu_n605), .A2(alu_n457), .A3(alu_n123), .A4(
        alu_n49), .Y(alu_n50) );
  INVX0_LVT alu_U69 ( .A(alu_n_T_101_24_), .Y(alu_n49) );
  AO22X1_LVT alu_U68 ( .A1(alu_io_in1[30]), .A2(alu_in2_inv_30_), .A3(alu_n47), 
        .A4(alu_n48), .Y(alu_n422) );
  INVX0_LVT alu_U67 ( .A(alu_in2_inv_30_), .Y(alu_n48) );
  INVX0_LVT alu_U66 ( .A(alu_io_in1[30]), .Y(alu_n47) );
  AO22X1_LVT alu_U65 ( .A1(alu_io_in1[15]), .A2(alu_in2_inv_15_), .A3(alu_n45), 
        .A4(alu_n46), .Y(alu_n331) );
  INVX0_LVT alu_U64 ( .A(alu_in2_inv_15_), .Y(alu_n46) );
  INVX0_LVT alu_U63 ( .A(alu_io_in1[15]), .Y(alu_n45) );
  AO22X1_LVT alu_U61 ( .A1(alu_n441), .A2(alu_n_T_101_50_), .A3(alu_n121), 
        .A4(alu_n_T_101_13_), .Y(alu_n43) );
  OAI21X1_LVT alu_U60 ( .A1(alu_n423), .A2(alu_n324), .A3(alu_n41), .Y(alu_n42) );
  NAND3X0_LVT alu_U59 ( .A1(alu_io_in1[13]), .A2(alu_io_in2[13]), .A3(alu_n122), .Y(alu_n41) );
  NAND4X0_LVT alu_U58 ( .A1(alu_n38), .A2(alu_n115), .A3(alu_n39), .A4(alu_n40), .Y(alu_io_out[38]) );
  NAND2X0_LVT alu_U57 ( .A1(alu_n602), .A2(io_dmem_req_bits_addr[38]), .Y(
        alu_n40) );
  AOI22X1_LVT alu_U56 ( .A1(alu_n_T_101_25_), .A2(alu_n598), .A3(
        alu_n_T_101_38_), .A4(alu_n124), .Y(alu_n39) );
  OA21X1_LVT alu_U55 ( .A1(alu_n605), .A2(alu_n456), .A3(alu_n37), .Y(alu_n38)
         );
  NAND3X0_LVT alu_U54 ( .A1(alu_io_in1[38]), .A2(alu_n603), .A3(alu_io_in2[38]), .Y(alu_n37) );
  AO22X1_LVT alu_U53 ( .A1(alu_io_in1[16]), .A2(alu_in2_inv_16_), .A3(alu_n35), 
        .A4(alu_n36), .Y(alu_n338) );
  INVX0_LVT alu_U52 ( .A(alu_in2_inv_16_), .Y(alu_n36) );
  INVX0_LVT alu_U51 ( .A(alu_io_in1[16]), .Y(alu_n35) );
  AO22X1_LVT alu_U50 ( .A1(alu_io_in1[10]), .A2(alu_in2_inv_10_), .A3(alu_n33), 
        .A4(alu_n34), .Y(alu_n307) );
  INVX0_LVT alu_U49 ( .A(alu_in2_inv_10_), .Y(alu_n34) );
  INVX0_LVT alu_U48 ( .A(alu_io_in1[10]), .Y(alu_n33) );
  AO22X1_LVT alu_U47 ( .A1(alu_io_in1[63]), .A2(alu_in2_inv_63_), .A3(alu_n31), 
        .A4(alu_n32), .Y(alu_n604) );
  INVX0_LVT alu_U46 ( .A(alu_in2_inv_63_), .Y(alu_n32) );
  INVX0_LVT alu_U45 ( .A(alu_io_in1[63]), .Y(alu_n31) );
  AO22X1_LVT alu_U44 ( .A1(alu_io_in1[13]), .A2(alu_in2_inv_13_), .A3(alu_n29), 
        .A4(alu_n30), .Y(alu_n324) );
  INVX0_LVT alu_U43 ( .A(alu_in2_inv_13_), .Y(alu_n30) );
  INVX0_LVT alu_U42 ( .A(alu_io_in1[13]), .Y(alu_n29) );
  AO22X1_LVT alu_U41 ( .A1(alu_io_in1[6]), .A2(alu_in2_inv_6_), .A3(alu_n27), 
        .A4(alu_n28), .Y(alu_n282) );
  INVX0_LVT alu_U40 ( .A(alu_in2_inv_6_), .Y(alu_n28) );
  INVX0_LVT alu_U39 ( .A(alu_io_in1[6]), .Y(alu_n27) );
  NAND4X0_LVT alu_U38 ( .A1(alu_n24), .A2(alu_n115), .A3(alu_n25), .A4(alu_n26), .Y(alu_io_out[37]) );
  NAND2X0_LVT alu_U37 ( .A1(alu_n602), .A2(io_dmem_req_bits_addr[37]), .Y(
        alu_n26) );
  AOI22X1_LVT alu_U36 ( .A1(alu_n_T_101_37_), .A2(alu_n124), .A3(
        alu_n_T_101_26_), .A4(alu_n598), .Y(alu_n25) );
  OA21X1_LVT alu_U35 ( .A1(alu_n605), .A2(alu_n455), .A3(alu_n23), .Y(alu_n24)
         );
  NAND3X0_LVT alu_U34 ( .A1(alu_io_in1[37]), .A2(alu_n603), .A3(alu_io_in2[37]), .Y(alu_n23) );
  AO22X1_LVT alu_U33 ( .A1(alu_io_in1[39]), .A2(alu_in2_inv_39_), .A3(alu_n21), 
        .A4(alu_n22), .Y(alu_n457) );
  INVX0_LVT alu_U32 ( .A(alu_in2_inv_39_), .Y(alu_n22) );
  INVX0_LVT alu_U31 ( .A(alu_io_in1[39]), .Y(alu_n21) );
  AO22X1_LVT alu_U30 ( .A1(alu_io_in1[7]), .A2(alu_in2_inv_7_), .A3(alu_n19), 
        .A4(alu_n20), .Y(alu_n288) );
  INVX0_LVT alu_U29 ( .A(alu_in2_inv_7_), .Y(alu_n20) );
  INVX0_LVT alu_U28 ( .A(alu_io_in1[7]), .Y(alu_n19) );
  AO22X1_LVT alu_U27 ( .A1(alu_io_in1[12]), .A2(alu_in2_inv_12_), .A3(alu_n17), 
        .A4(alu_n18), .Y(alu_n319) );
  INVX0_LVT alu_U26 ( .A(alu_in2_inv_12_), .Y(alu_n18) );
  INVX0_LVT alu_U25 ( .A(alu_io_in1[12]), .Y(alu_n17) );
  NAND4X0_LVT alu_U24 ( .A1(alu_n14), .A2(alu_n115), .A3(alu_n15), .A4(alu_n16), .Y(alu_io_out[36]) );
  NAND2X0_LVT alu_U23 ( .A1(alu_n602), .A2(io_dmem_req_bits_addr[36]), .Y(
        alu_n16) );
  AOI22X1_LVT alu_U22 ( .A1(alu_n_T_101_27_), .A2(alu_n598), .A3(
        alu_n_T_101_36_), .A4(alu_n124), .Y(alu_n15) );
  OA21X1_LVT alu_U21 ( .A1(alu_n605), .A2(alu_n454), .A3(alu_n13), .Y(alu_n14)
         );
  NAND3X0_LVT alu_U20 ( .A1(alu_io_in1[36]), .A2(alu_n603), .A3(alu_io_in2[36]), .Y(alu_n13) );
  AO22X1_LVT alu_U19 ( .A1(alu_io_in1[14]), .A2(alu_in2_inv_14_), .A3(alu_n11), 
        .A4(alu_n12), .Y(alu_n326) );
  INVX0_LVT alu_U18 ( .A(alu_in2_inv_14_), .Y(alu_n12) );
  INVX0_LVT alu_U17 ( .A(alu_io_in1[14]), .Y(alu_n11) );
  NAND4X0_LVT alu_U16 ( .A1(alu_n8), .A2(alu_n115), .A3(alu_n9), .A4(alu_n10), 
        .Y(alu_io_out[35]) );
  NAND3X0_LVT alu_U15 ( .A1(alu_io_in1[35]), .A2(alu_io_in2[35]), .A3(alu_n603), .Y(alu_n10) );
  AOI22X1_LVT alu_U14 ( .A1(alu_n602), .A2(io_dmem_req_bits_addr[35]), .A3(
        alu_n124), .A4(alu_n_T_101_35_), .Y(alu_n9) );
  OA22X1_LVT alu_U13 ( .A1(alu_n605), .A2(alu_n453), .A3(alu_n123), .A4(alu_n7), .Y(alu_n8) );
  INVX0_LVT alu_U12 ( .A(alu_n_T_101_28_), .Y(alu_n7) );
  NAND4X0_LVT alu_U11 ( .A1(alu_n115), .A2(alu_n4), .A3(alu_n5), .A4(alu_n6), 
        .Y(alu_io_out[34]) );
  NAND2X0_LVT alu_U10 ( .A1(io_dmem_req_bits_addr[34]), .A2(alu_n602), .Y(
        alu_n6) );
  AOI22X1_LVT alu_U9 ( .A1(alu_n124), .A2(alu_n_T_101_34_), .A3(alu_n598), 
        .A4(alu_n_T_101_29_), .Y(alu_n5) );
  OA21X1_LVT alu_U8 ( .A1(alu_n605), .A2(alu_n452), .A3(alu_n3), .Y(alu_n4) );
  NAND3X0_LVT alu_U7 ( .A1(alu_io_in1[34]), .A2(alu_io_in2[34]), .A3(alu_n603), 
        .Y(alu_n3) );
  AO22X1_LVT alu_U6 ( .A1(alu_io_in1[25]), .A2(alu_in2_inv_25_), .A3(alu_n1), 
        .A4(alu_n2), .Y(alu_n392) );
  INVX0_LVT alu_U5 ( .A(alu_in2_inv_25_), .Y(alu_n2) );
  INVX0_LVT alu_U4 ( .A(alu_io_in1[25]), .Y(alu_n1) );
  AO221X1_LVT alu_U3 ( .A1(1'b1), .A2(alu_n42), .A3(io_dmem_req_bits_addr[13]), 
        .A4(alu_n434), .A5(alu_n43), .Y(alu_io_out[13]) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U848 ( .A(alu_DP_OP_31J40_124_1870_n442), 
        .B(alu_in2_inv_1_), .CI(alu_io_in1[1]), .S(io_dmem_req_bits_addr[1])
         );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U847 ( .A1(alu_in2_inv_1_), .A2(
        alu_io_in1[1]), .Y(alu_DP_OP_31J40_124_1870_n915) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U846 ( .A1(alu_in2_inv_1_), .A2(
        alu_io_in1[1]), .Y(alu_DP_OP_31J40_124_1870_n916) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U845 ( .A1(alu_DP_OP_31J40_124_1870_n442), .A2(alu_DP_OP_31J40_124_1870_n915), .A3(alu_DP_OP_31J40_124_1870_n916), .Y(
        alu_DP_OP_31J40_124_1870_n917) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U844 ( .A(alu_io_in1[2]), .B(
        alu_in2_inv_2_), .CI(alu_DP_OP_31J40_124_1870_n917), .S(
        io_dmem_req_bits_addr[2]) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U843 ( .A1(alu_io_in1[2]), .A2(
        alu_in2_inv_2_), .Y(alu_DP_OP_31J40_124_1870_n914) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U842 ( .A1(alu_io_in1[2]), .A2(
        alu_in2_inv_2_), .A3(alu_DP_OP_31J40_124_1870_n916), .A4(
        alu_DP_OP_31J40_124_1870_n914), .Y(alu_DP_OP_31J40_124_1870_n913) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U841 ( .A(alu_DP_OP_31J40_124_1870_n906), 
        .B(alu_io_in1[3]), .CI(alu_in2_inv_3_), .S(io_dmem_req_bits_addr[3])
         );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U840 ( .A1(alu_io_in1[3]), .A2(
        alu_in2_inv_3_), .Y(alu_DP_OP_31J40_124_1870_n910) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U839 ( .A1(alu_DP_OP_31J40_124_1870_n906), .A2(alu_DP_OP_31J40_124_1870_n910), .A3(alu_io_in1[3]), .A4(alu_in2_inv_3_), 
        .Y(alu_DP_OP_31J40_124_1870_n912) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U838 ( .A(alu_io_in1[4]), .B(
        alu_in2_inv_4_), .CI(alu_DP_OP_31J40_124_1870_n912), .S(
        io_dmem_req_bits_addr[4]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U837 ( .A1(alu_io_in1[4]), .A2(
        alu_in2_inv_4_), .A3(alu_io_in1[3]), .A4(alu_in2_inv_3_), .Y(
        alu_DP_OP_31J40_124_1870_n907) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U836 ( .A1(alu_io_in1[4]), .A2(
        alu_in2_inv_4_), .Y(alu_DP_OP_31J40_124_1870_n911) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U835 ( .A1(alu_io_in1[4]), .A2(
        alu_in2_inv_4_), .A3(alu_DP_OP_31J40_124_1870_n910), .A4(
        alu_DP_OP_31J40_124_1870_n911), .Y(alu_DP_OP_31J40_124_1870_n902) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U834 ( .A1(alu_DP_OP_31J40_124_1870_n907), .A2(alu_DP_OP_31J40_124_1870_n906), .A3(alu_DP_OP_31J40_124_1870_n902), .Y(
        alu_DP_OP_31J40_124_1870_n909) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U833 ( .A(alu_io_in1[5]), .B(
        alu_in2_inv_5_), .CI(alu_DP_OP_31J40_124_1870_n909), .S(
        io_dmem_req_bits_addr[5]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U832 ( .A1(alu_io_in1[5]), .A2(
        alu_in2_inv_5_), .Y(alu_DP_OP_31J40_124_1870_n904) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U831 ( .A1(
        alu_DP_OP_31J40_124_1870_n909), .A2(alu_io_in1[5]), .A3(
        alu_DP_OP_31J40_124_1870_n909), .A4(alu_in2_inv_5_), .A5(
        alu_DP_OP_31J40_124_1870_n904), .Y(alu_DP_OP_31J40_124_1870_n908) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U830 ( .A(alu_io_in1[6]), .B(
        alu_in2_inv_6_), .CI(alu_DP_OP_31J40_124_1870_n908), .S(
        io_dmem_req_bits_addr[6]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U829 ( .A1(alu_io_in1[6]), .A2(
        alu_in2_inv_6_), .A3(alu_io_in1[5]), .A4(alu_in2_inv_5_), .Y(
        alu_DP_OP_31J40_124_1870_n900) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U828 ( .A1(alu_DP_OP_31J40_124_1870_n906), .A2(alu_DP_OP_31J40_124_1870_n907), .Y(alu_DP_OP_31J40_124_1870_n901) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U827 ( .A1(alu_io_in1[6]), .A2(
        alu_in2_inv_6_), .Y(alu_DP_OP_31J40_124_1870_n905) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U826 ( .A1(alu_io_in1[6]), .A2(
        alu_in2_inv_6_), .A3(alu_DP_OP_31J40_124_1870_n904), .A4(
        alu_DP_OP_31J40_124_1870_n905), .Y(alu_DP_OP_31J40_124_1870_n903) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U825 ( .A1(
        alu_DP_OP_31J40_124_1870_n900), .A2(alu_DP_OP_31J40_124_1870_n901), 
        .A3(alu_DP_OP_31J40_124_1870_n900), .A4(alu_DP_OP_31J40_124_1870_n902), 
        .A5(alu_DP_OP_31J40_124_1870_n903), .Y(alu_DP_OP_31J40_124_1870_n876)
         );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U824 ( .A(alu_io_in1[7]), .B(
        alu_in2_inv_7_), .CI(alu_DP_OP_31J40_124_1870_n876), .S(
        io_dmem_req_bits_addr[7]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U823 ( .A1(alu_io_in1[7]), .A2(
        alu_in2_inv_7_), .Y(alu_DP_OP_31J40_124_1870_n897) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U822 ( .A1(
        alu_DP_OP_31J40_124_1870_n876), .A2(alu_io_in1[7]), .A3(
        alu_DP_OP_31J40_124_1870_n876), .A4(alu_in2_inv_7_), .A5(
        alu_DP_OP_31J40_124_1870_n897), .Y(alu_DP_OP_31J40_124_1870_n899) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U821 ( .A(alu_io_in1[8]), .B(
        alu_in2_inv_8_), .CI(alu_DP_OP_31J40_124_1870_n899), .S(
        io_dmem_req_bits_addr[8]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U820 ( .A1(alu_io_in1[8]), .A2(
        alu_in2_inv_8_), .A3(alu_io_in1[7]), .A4(alu_in2_inv_7_), .Y(
        alu_DP_OP_31J40_124_1870_n894) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U819 ( .A1(alu_io_in1[8]), .A2(
        alu_in2_inv_8_), .Y(alu_DP_OP_31J40_124_1870_n898) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U818 ( .A1(alu_io_in1[8]), .A2(
        alu_in2_inv_8_), .A3(alu_DP_OP_31J40_124_1870_n897), .A4(
        alu_DP_OP_31J40_124_1870_n898), .Y(alu_DP_OP_31J40_124_1870_n893) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U817 ( .A1(alu_DP_OP_31J40_124_1870_n894), .A2(alu_DP_OP_31J40_124_1870_n876), .A3(alu_DP_OP_31J40_124_1870_n893), .Y(
        alu_DP_OP_31J40_124_1870_n896) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U816 ( .A(alu_io_in1[9]), .B(
        alu_in2_inv_9_), .CI(alu_DP_OP_31J40_124_1870_n896), .S(
        io_dmem_req_bits_addr[9]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U815 ( .A1(alu_io_in1[9]), .A2(
        alu_in2_inv_9_), .Y(alu_DP_OP_31J40_124_1870_n890) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U814 ( .A1(alu_DP_OP_31J40_124_1870_n890), .A2(alu_DP_OP_31J40_124_1870_n896), .A3(alu_io_in1[9]), .A4(alu_in2_inv_9_), 
        .Y(alu_DP_OP_31J40_124_1870_n895) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U813 ( .A(alu_io_in1[10]), .B(
        alu_in2_inv_10_), .CI(alu_DP_OP_31J40_124_1870_n895), .S(
        io_dmem_req_bits_addr[10]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U812 ( .A1(alu_io_in1[10]), .A2(
        alu_in2_inv_10_), .A3(alu_io_in1[9]), .A4(alu_in2_inv_9_), .Y(
        alu_DP_OP_31J40_124_1870_n892) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U811 ( .A1(alu_DP_OP_31J40_124_1870_n892), .A2(alu_DP_OP_31J40_124_1870_n894), .Y(alu_DP_OP_31J40_124_1870_n875) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U810 ( .A1(alu_in2_inv_10_), .A2(
        alu_io_in1[10]), .Y(alu_DP_OP_31J40_124_1870_n891) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U809 ( .A1(alu_io_in1[10]), .A2(
        alu_in2_inv_10_), .A3(alu_DP_OP_31J40_124_1870_n890), .A4(
        alu_DP_OP_31J40_124_1870_n891), .A5(alu_DP_OP_31J40_124_1870_n892), 
        .A6(alu_DP_OP_31J40_124_1870_n893), .Y(alu_DP_OP_31J40_124_1870_n879)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U808 ( .A1(alu_DP_OP_31J40_124_1870_n875), .A2(alu_DP_OP_31J40_124_1870_n876), .A3(alu_DP_OP_31J40_124_1870_n879), .Y(
        alu_DP_OP_31J40_124_1870_n886) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U807 ( .A(alu_io_in1[11]), .B(
        alu_in2_inv_11_), .CI(alu_DP_OP_31J40_124_1870_n886), .S(
        io_dmem_req_bits_addr[11]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U806 ( .A1(alu_io_in1[11]), .A2(
        alu_in2_inv_11_), .Y(alu_DP_OP_31J40_124_1870_n887) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U805 ( .A1(alu_DP_OP_31J40_124_1870_n887), .A2(alu_DP_OP_31J40_124_1870_n886), .A3(alu_io_in1[11]), .A4(alu_in2_inv_11_), .Y(alu_DP_OP_31J40_124_1870_n889) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U804 ( .A(alu_io_in1[12]), .B(
        alu_in2_inv_12_), .CI(alu_DP_OP_31J40_124_1870_n889), .S(
        io_dmem_req_bits_addr[12]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U803 ( .A1(alu_io_in1[12]), .A2(
        alu_in2_inv_12_), .A3(alu_io_in1[11]), .A4(alu_in2_inv_11_), .Y(
        alu_DP_OP_31J40_124_1870_n883) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U802 ( .A1(alu_io_in1[12]), .A2(
        alu_in2_inv_12_), .Y(alu_DP_OP_31J40_124_1870_n888) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U801 ( .A1(alu_io_in1[12]), .A2(
        alu_in2_inv_12_), .A3(alu_DP_OP_31J40_124_1870_n887), .A4(
        alu_DP_OP_31J40_124_1870_n888), .Y(alu_DP_OP_31J40_124_1870_n878) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U800 ( .A1(alu_DP_OP_31J40_124_1870_n883), .A2(alu_DP_OP_31J40_124_1870_n886), .A3(alu_DP_OP_31J40_124_1870_n878), .Y(
        alu_DP_OP_31J40_124_1870_n885) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U799 ( .A(alu_io_in1[13]), .B(
        alu_in2_inv_13_), .CI(alu_DP_OP_31J40_124_1870_n885), .S(
        io_dmem_req_bits_addr[13]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U798 ( .A1(alu_io_in1[13]), .A2(
        alu_in2_inv_13_), .Y(alu_DP_OP_31J40_124_1870_n881) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U797 ( .A1(alu_DP_OP_31J40_124_1870_n881), .A2(alu_DP_OP_31J40_124_1870_n885), .A3(alu_io_in1[13]), .A4(alu_in2_inv_13_), .Y(alu_DP_OP_31J40_124_1870_n884) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U796 ( .A(alu_io_in1[14]), .B(
        alu_in2_inv_14_), .CI(alu_DP_OP_31J40_124_1870_n884), .S(
        io_dmem_req_bits_addr[14]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U795 ( .A1(alu_io_in1[14]), .A2(
        alu_in2_inv_14_), .A3(alu_io_in1[13]), .A4(alu_in2_inv_13_), .Y(
        alu_DP_OP_31J40_124_1870_n877) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U794 ( .A1(alu_DP_OP_31J40_124_1870_n877), .A2(alu_DP_OP_31J40_124_1870_n883), .Y(alu_DP_OP_31J40_124_1870_n874) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U793 ( .A1(alu_in2_inv_14_), .A2(
        alu_io_in1[14]), .Y(alu_DP_OP_31J40_124_1870_n882) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U792 ( .A1(alu_io_in1[14]), .A2(
        alu_in2_inv_14_), .A3(alu_DP_OP_31J40_124_1870_n881), .A4(
        alu_DP_OP_31J40_124_1870_n882), .Y(alu_DP_OP_31J40_124_1870_n880) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U791 ( .A1(
        alu_DP_OP_31J40_124_1870_n877), .A2(alu_DP_OP_31J40_124_1870_n878), 
        .A3(alu_DP_OP_31J40_124_1870_n879), .A4(alu_DP_OP_31J40_124_1870_n874), 
        .A5(alu_DP_OP_31J40_124_1870_n880), .Y(alu_DP_OP_31J40_124_1870_n873)
         );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U790 ( .A(alu_DP_OP_31J40_124_1870_n827), 
        .B(alu_io_in1[15]), .CI(alu_in2_inv_15_), .S(io_dmem_req_bits_addr[15]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U789 ( .A1(alu_io_in1[15]), .A2(
        alu_in2_inv_15_), .Y(alu_DP_OP_31J40_124_1870_n870) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U788 ( .A1(alu_DP_OP_31J40_124_1870_n827), .A2(alu_DP_OP_31J40_124_1870_n870), .A3(alu_io_in1[15]), .A4(alu_in2_inv_15_), .Y(alu_DP_OP_31J40_124_1870_n872) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U787 ( .A(alu_io_in1[16]), .B(
        alu_in2_inv_16_), .CI(alu_DP_OP_31J40_124_1870_n872), .S(
        io_dmem_req_bits_addr[16]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U786 ( .A1(alu_io_in1[16]), .A2(
        alu_in2_inv_16_), .A3(alu_io_in1[15]), .A4(alu_in2_inv_15_), .Y(
        alu_DP_OP_31J40_124_1870_n867) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U785 ( .A1(alu_io_in1[16]), .A2(
        alu_in2_inv_16_), .Y(alu_DP_OP_31J40_124_1870_n871) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U784 ( .A1(alu_io_in1[16]), .A2(
        alu_in2_inv_16_), .A3(alu_DP_OP_31J40_124_1870_n870), .A4(
        alu_DP_OP_31J40_124_1870_n871), .Y(alu_DP_OP_31J40_124_1870_n866) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U783 ( .A1(alu_DP_OP_31J40_124_1870_n867), .A2(alu_DP_OP_31J40_124_1870_n827), .A3(alu_DP_OP_31J40_124_1870_n866), .Y(
        alu_DP_OP_31J40_124_1870_n869) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U782 ( .A(alu_io_in1[17]), .B(
        alu_in2_inv_17_), .CI(alu_DP_OP_31J40_124_1870_n869), .S(
        io_dmem_req_bits_addr[17]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U781 ( .A1(alu_io_in1[17]), .A2(
        alu_in2_inv_17_), .Y(alu_DP_OP_31J40_124_1870_n863) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U780 ( .A1(
        alu_DP_OP_31J40_124_1870_n869), .A2(alu_io_in1[17]), .A3(
        alu_DP_OP_31J40_124_1870_n869), .A4(alu_in2_inv_17_), .A5(
        alu_DP_OP_31J40_124_1870_n863), .Y(alu_DP_OP_31J40_124_1870_n868) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U779 ( .A(alu_io_in1[18]), .B(
        alu_in2_inv_18_), .CI(alu_DP_OP_31J40_124_1870_n868), .S(
        io_dmem_req_bits_addr[18]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U778 ( .A1(alu_io_in1[18]), .A2(
        alu_in2_inv_18_), .A3(alu_io_in1[17]), .A4(alu_in2_inv_17_), .Y(
        alu_DP_OP_31J40_124_1870_n865) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U777 ( .A1(alu_DP_OP_31J40_124_1870_n865), .A2(alu_DP_OP_31J40_124_1870_n867), .Y(alu_DP_OP_31J40_124_1870_n855) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U776 ( .A1(alu_in2_inv_18_), .A2(
        alu_io_in1[18]), .Y(alu_DP_OP_31J40_124_1870_n864) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U775 ( .A1(alu_io_in1[18]), .A2(
        alu_in2_inv_18_), .A3(alu_DP_OP_31J40_124_1870_n863), .A4(
        alu_DP_OP_31J40_124_1870_n864), .A5(alu_DP_OP_31J40_124_1870_n865), 
        .A6(alu_DP_OP_31J40_124_1870_n866), .Y(alu_DP_OP_31J40_124_1870_n850)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U774 ( .A1(alu_DP_OP_31J40_124_1870_n827), .A2(alu_DP_OP_31J40_124_1870_n855), .A3(alu_DP_OP_31J40_124_1870_n850), .Y(
        alu_DP_OP_31J40_124_1870_n859) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U773 ( .A(alu_io_in1[19]), .B(
        alu_in2_inv_19_), .CI(alu_DP_OP_31J40_124_1870_n859), .S(
        io_dmem_req_bits_addr[19]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U772 ( .A1(alu_io_in1[19]), .A2(
        alu_in2_inv_19_), .Y(alu_DP_OP_31J40_124_1870_n860) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U771 ( .A1(
        alu_DP_OP_31J40_124_1870_n859), .A2(alu_io_in1[19]), .A3(
        alu_DP_OP_31J40_124_1870_n859), .A4(alu_in2_inv_19_), .A5(
        alu_DP_OP_31J40_124_1870_n860), .Y(alu_DP_OP_31J40_124_1870_n862) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U770 ( .A(alu_io_in1[20]), .B(
        alu_in2_inv_20_), .CI(alu_DP_OP_31J40_124_1870_n862), .S(
        io_dmem_req_bits_addr[20]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U769 ( .A1(alu_io_in1[20]), .A2(
        alu_in2_inv_20_), .A3(alu_io_in1[19]), .A4(alu_in2_inv_19_), .Y(
        alu_DP_OP_31J40_124_1870_n856) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U768 ( .A1(alu_io_in1[20]), .A2(
        alu_in2_inv_20_), .Y(alu_DP_OP_31J40_124_1870_n861) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U767 ( .A1(alu_io_in1[20]), .A2(
        alu_in2_inv_20_), .A3(alu_DP_OP_31J40_124_1870_n860), .A4(
        alu_DP_OP_31J40_124_1870_n861), .Y(alu_DP_OP_31J40_124_1870_n849) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U766 ( .A1(alu_DP_OP_31J40_124_1870_n856), .A2(alu_DP_OP_31J40_124_1870_n859), .A3(alu_DP_OP_31J40_124_1870_n849), .Y(
        alu_DP_OP_31J40_124_1870_n858) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U765 ( .A(alu_io_in1[21]), .B(
        alu_in2_inv_21_), .CI(alu_DP_OP_31J40_124_1870_n858), .S(
        io_dmem_req_bits_addr[21]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U764 ( .A1(alu_io_in1[21]), .A2(
        alu_in2_inv_21_), .Y(alu_DP_OP_31J40_124_1870_n853) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U763 ( .A1(
        alu_DP_OP_31J40_124_1870_n858), .A2(alu_io_in1[21]), .A3(
        alu_DP_OP_31J40_124_1870_n858), .A4(alu_in2_inv_21_), .A5(
        alu_DP_OP_31J40_124_1870_n853), .Y(alu_DP_OP_31J40_124_1870_n857) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U762 ( .A(alu_io_in1[22]), .B(
        alu_in2_inv_22_), .CI(alu_DP_OP_31J40_124_1870_n857), .S(
        io_dmem_req_bits_addr[22]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U761 ( .A1(alu_io_in1[22]), .A2(
        alu_in2_inv_22_), .A3(alu_io_in1[21]), .A4(alu_in2_inv_21_), .Y(
        alu_DP_OP_31J40_124_1870_n848) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U760 ( .A1(alu_DP_OP_31J40_124_1870_n848), .A2(alu_DP_OP_31J40_124_1870_n856), .Y(alu_DP_OP_31J40_124_1870_n851) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U759 ( .A1(alu_DP_OP_31J40_124_1870_n855), .A2(alu_DP_OP_31J40_124_1870_n851), .Y(alu_DP_OP_31J40_124_1870_n828) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U758 ( .A1(alu_in2_inv_22_), .A2(
        alu_io_in1[22]), .Y(alu_DP_OP_31J40_124_1870_n854) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U757 ( .A1(alu_io_in1[22]), .A2(
        alu_in2_inv_22_), .A3(alu_DP_OP_31J40_124_1870_n853), .A4(
        alu_DP_OP_31J40_124_1870_n854), .Y(alu_DP_OP_31J40_124_1870_n852) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U756 ( .A1(
        alu_DP_OP_31J40_124_1870_n848), .A2(alu_DP_OP_31J40_124_1870_n849), 
        .A3(alu_DP_OP_31J40_124_1870_n850), .A4(alu_DP_OP_31J40_124_1870_n851), 
        .A5(alu_DP_OP_31J40_124_1870_n852), .Y(alu_DP_OP_31J40_124_1870_n817)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U755 ( .A1(alu_DP_OP_31J40_124_1870_n828), .A2(alu_DP_OP_31J40_124_1870_n827), .A3(alu_DP_OP_31J40_124_1870_n817), .Y(
        alu_DP_OP_31J40_124_1870_n837) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U754 ( .A(alu_io_in1[23]), .B(
        alu_in2_inv_23_), .CI(alu_DP_OP_31J40_124_1870_n837), .S(
        io_dmem_req_bits_addr[23]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U753 ( .A1(alu_io_in1[23]), .A2(
        alu_in2_inv_23_), .Y(alu_DP_OP_31J40_124_1870_n845) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U752 ( .A1(
        alu_DP_OP_31J40_124_1870_n837), .A2(alu_io_in1[23]), .A3(
        alu_DP_OP_31J40_124_1870_n837), .A4(alu_in2_inv_23_), .A5(
        alu_DP_OP_31J40_124_1870_n845), .Y(alu_DP_OP_31J40_124_1870_n847) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U751 ( .A(alu_io_in1[24]), .B(
        alu_in2_inv_24_), .CI(alu_DP_OP_31J40_124_1870_n847), .S(
        io_dmem_req_bits_addr[24]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U750 ( .A1(alu_io_in1[24]), .A2(
        alu_in2_inv_24_), .A3(alu_io_in1[23]), .A4(alu_in2_inv_23_), .Y(
        alu_DP_OP_31J40_124_1870_n842) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U749 ( .A1(alu_io_in1[24]), .A2(
        alu_in2_inv_24_), .Y(alu_DP_OP_31J40_124_1870_n846) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U748 ( .A1(alu_io_in1[24]), .A2(
        alu_in2_inv_24_), .A3(alu_DP_OP_31J40_124_1870_n845), .A4(
        alu_DP_OP_31J40_124_1870_n846), .Y(alu_DP_OP_31J40_124_1870_n841) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U747 ( .A1(alu_DP_OP_31J40_124_1870_n842), .A2(alu_DP_OP_31J40_124_1870_n837), .A3(alu_DP_OP_31J40_124_1870_n841), .Y(
        alu_DP_OP_31J40_124_1870_n844) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U746 ( .A(alu_io_in1[25]), .B(
        alu_in2_inv_25_), .CI(alu_DP_OP_31J40_124_1870_n844), .S(
        io_dmem_req_bits_addr[25]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U745 ( .A1(alu_io_in1[25]), .A2(
        alu_in2_inv_25_), .Y(alu_DP_OP_31J40_124_1870_n838) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U744 ( .A1(
        alu_DP_OP_31J40_124_1870_n844), .A2(alu_io_in1[25]), .A3(
        alu_DP_OP_31J40_124_1870_n844), .A4(alu_in2_inv_25_), .A5(
        alu_DP_OP_31J40_124_1870_n838), .Y(alu_DP_OP_31J40_124_1870_n843) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U743 ( .A(alu_io_in1[26]), .B(
        alu_in2_inv_26_), .CI(alu_DP_OP_31J40_124_1870_n843), .S(
        io_dmem_req_bits_addr[26]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U742 ( .A1(alu_io_in1[26]), .A2(
        alu_in2_inv_26_), .A3(alu_io_in1[25]), .A4(alu_in2_inv_25_), .Y(
        alu_DP_OP_31J40_124_1870_n840) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U741 ( .A1(alu_DP_OP_31J40_124_1870_n840), .A2(alu_DP_OP_31J40_124_1870_n842), .Y(alu_DP_OP_31J40_124_1870_n829) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U740 ( .A1(alu_in2_inv_26_), .A2(
        alu_io_in1[26]), .Y(alu_DP_OP_31J40_124_1870_n839) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U739 ( .A1(alu_io_in1[26]), .A2(
        alu_in2_inv_26_), .A3(alu_DP_OP_31J40_124_1870_n838), .A4(
        alu_DP_OP_31J40_124_1870_n839), .A5(alu_DP_OP_31J40_124_1870_n840), 
        .A6(alu_DP_OP_31J40_124_1870_n841), .Y(alu_DP_OP_31J40_124_1870_n822)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U738 ( .A1(alu_DP_OP_31J40_124_1870_n829), .A2(alu_DP_OP_31J40_124_1870_n837), .A3(alu_DP_OP_31J40_124_1870_n822), .Y(
        alu_DP_OP_31J40_124_1870_n833) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U737 ( .A(alu_io_in1[27]), .B(
        alu_in2_inv_27_), .CI(alu_DP_OP_31J40_124_1870_n833), .S(
        io_dmem_req_bits_addr[27]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U736 ( .A1(alu_io_in1[27]), .A2(
        alu_in2_inv_27_), .Y(alu_DP_OP_31J40_124_1870_n834) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U735 ( .A1(
        alu_DP_OP_31J40_124_1870_n833), .A2(alu_io_in1[27]), .A3(
        alu_DP_OP_31J40_124_1870_n833), .A4(alu_in2_inv_27_), .A5(
        alu_DP_OP_31J40_124_1870_n834), .Y(alu_DP_OP_31J40_124_1870_n836) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U734 ( .A(alu_io_in1[28]), .B(
        alu_in2_inv_28_), .CI(alu_DP_OP_31J40_124_1870_n836), .S(
        io_dmem_req_bits_addr[28]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U733 ( .A1(alu_io_in1[28]), .A2(
        alu_in2_inv_28_), .A3(alu_io_in1[27]), .A4(alu_in2_inv_27_), .Y(
        alu_DP_OP_31J40_124_1870_n830) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U732 ( .A1(alu_io_in1[28]), .A2(
        alu_in2_inv_28_), .Y(alu_DP_OP_31J40_124_1870_n835) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U731 ( .A1(alu_io_in1[28]), .A2(
        alu_in2_inv_28_), .A3(alu_DP_OP_31J40_124_1870_n834), .A4(
        alu_DP_OP_31J40_124_1870_n835), .Y(alu_DP_OP_31J40_124_1870_n821) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U730 ( .A1(alu_DP_OP_31J40_124_1870_n830), .A2(alu_DP_OP_31J40_124_1870_n833), .A3(alu_DP_OP_31J40_124_1870_n821), .Y(
        alu_DP_OP_31J40_124_1870_n832) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U729 ( .A(alu_io_in1[29]), .B(
        alu_in2_inv_29_), .CI(alu_DP_OP_31J40_124_1870_n832), .S(
        io_dmem_req_bits_addr[29]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U728 ( .A1(alu_io_in1[29]), .A2(
        alu_in2_inv_29_), .Y(alu_DP_OP_31J40_124_1870_n825) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U727 ( .A1(
        alu_DP_OP_31J40_124_1870_n832), .A2(alu_io_in1[29]), .A3(
        alu_DP_OP_31J40_124_1870_n832), .A4(alu_in2_inv_29_), .A5(
        alu_DP_OP_31J40_124_1870_n825), .Y(alu_DP_OP_31J40_124_1870_n831) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U726 ( .A(alu_io_in1[30]), .B(
        alu_in2_inv_30_), .CI(alu_DP_OP_31J40_124_1870_n831), .S(
        io_dmem_req_bits_addr[30]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U725 ( .A1(alu_io_in1[30]), .A2(
        alu_in2_inv_30_), .A3(alu_io_in1[29]), .A4(alu_in2_inv_29_), .Y(
        alu_DP_OP_31J40_124_1870_n820) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U724 ( .A1(alu_DP_OP_31J40_124_1870_n820), .A2(alu_DP_OP_31J40_124_1870_n830), .Y(alu_DP_OP_31J40_124_1870_n823) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U723 ( .A1(alu_DP_OP_31J40_124_1870_n829), .A2(alu_DP_OP_31J40_124_1870_n823), .Y(alu_DP_OP_31J40_124_1870_n816) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U722 ( .A1(alu_DP_OP_31J40_124_1870_n827), .A2(alu_DP_OP_31J40_124_1870_n828), .Y(alu_DP_OP_31J40_124_1870_n818) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U721 ( .A1(alu_in2_inv_30_), .A2(
        alu_io_in1[30]), .Y(alu_DP_OP_31J40_124_1870_n826) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U720 ( .A1(alu_io_in1[30]), .A2(
        alu_in2_inv_30_), .A3(alu_DP_OP_31J40_124_1870_n825), .A4(
        alu_DP_OP_31J40_124_1870_n826), .Y(alu_DP_OP_31J40_124_1870_n824) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U719 ( .A1(
        alu_DP_OP_31J40_124_1870_n820), .A2(alu_DP_OP_31J40_124_1870_n821), 
        .A3(alu_DP_OP_31J40_124_1870_n822), .A4(alu_DP_OP_31J40_124_1870_n823), 
        .A5(alu_DP_OP_31J40_124_1870_n824), .Y(alu_DP_OP_31J40_124_1870_n819)
         );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U718 ( .A1(
        alu_DP_OP_31J40_124_1870_n816), .A2(alu_DP_OP_31J40_124_1870_n817), 
        .A3(alu_DP_OP_31J40_124_1870_n816), .A4(alu_DP_OP_31J40_124_1870_n818), 
        .A5(alu_DP_OP_31J40_124_1870_n819), .Y(alu_DP_OP_31J40_124_1870_n708)
         );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U717 ( .A(alu_io_in1[31]), .B(
        alu_in2_inv_31_), .CI(alu_DP_OP_31J40_124_1870_n708), .S(
        io_dmem_req_bits_addr[31]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U716 ( .A1(alu_io_in1[31]), .A2(
        alu_in2_inv_31_), .Y(alu_DP_OP_31J40_124_1870_n813) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U715 ( .A1(
        alu_DP_OP_31J40_124_1870_n708), .A2(alu_io_in1[31]), .A3(
        alu_DP_OP_31J40_124_1870_n708), .A4(alu_in2_inv_31_), .A5(
        alu_DP_OP_31J40_124_1870_n813), .Y(alu_DP_OP_31J40_124_1870_n815) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U714 ( .A(alu_io_in1[32]), .B(
        alu_in2_inv_32_), .CI(alu_DP_OP_31J40_124_1870_n815), .S(
        io_dmem_req_bits_addr[32]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U713 ( .A1(alu_io_in1[32]), .A2(
        alu_in2_inv_32_), .A3(alu_io_in1[31]), .A4(alu_in2_inv_31_), .Y(
        alu_DP_OP_31J40_124_1870_n810) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U712 ( .A1(alu_io_in1[32]), .A2(
        alu_in2_inv_32_), .Y(alu_DP_OP_31J40_124_1870_n814) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U711 ( .A1(alu_io_in1[32]), .A2(
        alu_in2_inv_32_), .A3(alu_DP_OP_31J40_124_1870_n813), .A4(
        alu_DP_OP_31J40_124_1870_n814), .Y(alu_DP_OP_31J40_124_1870_n809) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U710 ( .A1(alu_DP_OP_31J40_124_1870_n810), .A2(alu_DP_OP_31J40_124_1870_n708), .A3(alu_DP_OP_31J40_124_1870_n809), .Y(
        alu_DP_OP_31J40_124_1870_n812) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U709 ( .A(alu_io_in1[33]), .B(
        alu_in2_inv_33_), .CI(alu_DP_OP_31J40_124_1870_n812), .S(
        io_dmem_req_bits_addr[33]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U708 ( .A1(alu_io_in1[33]), .A2(
        alu_in2_inv_33_), .Y(alu_DP_OP_31J40_124_1870_n806) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U707 ( .A1(alu_DP_OP_31J40_124_1870_n806), .A2(alu_DP_OP_31J40_124_1870_n812), .A3(alu_io_in1[33]), .A4(alu_in2_inv_33_), .Y(alu_DP_OP_31J40_124_1870_n811) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U706 ( .A(alu_io_in1[34]), .B(
        alu_in2_inv_34_), .CI(alu_DP_OP_31J40_124_1870_n811), .S(
        io_dmem_req_bits_addr[34]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U705 ( .A1(alu_io_in1[34]), .A2(
        alu_in2_inv_34_), .A3(alu_io_in1[33]), .A4(alu_in2_inv_33_), .Y(
        alu_DP_OP_31J40_124_1870_n808) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U704 ( .A1(alu_DP_OP_31J40_124_1870_n808), .A2(alu_DP_OP_31J40_124_1870_n810), .Y(alu_DP_OP_31J40_124_1870_n798) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U703 ( .A1(alu_in2_inv_34_), .A2(
        alu_io_in1[34]), .Y(alu_DP_OP_31J40_124_1870_n807) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U702 ( .A1(alu_io_in1[34]), .A2(
        alu_in2_inv_34_), .A3(alu_DP_OP_31J40_124_1870_n806), .A4(
        alu_DP_OP_31J40_124_1870_n807), .A5(alu_DP_OP_31J40_124_1870_n808), 
        .A6(alu_DP_OP_31J40_124_1870_n809), .Y(alu_DP_OP_31J40_124_1870_n793)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U701 ( .A1(alu_DP_OP_31J40_124_1870_n798), .A2(alu_DP_OP_31J40_124_1870_n708), .A3(alu_DP_OP_31J40_124_1870_n793), .Y(
        alu_DP_OP_31J40_124_1870_n802) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U700 ( .A(alu_io_in1[35]), .B(
        alu_in2_inv_35_), .CI(alu_DP_OP_31J40_124_1870_n802), .S(
        io_dmem_req_bits_addr[35]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U699 ( .A1(alu_io_in1[35]), .A2(
        alu_in2_inv_35_), .Y(alu_DP_OP_31J40_124_1870_n803) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U698 ( .A1(alu_DP_OP_31J40_124_1870_n803), .A2(alu_DP_OP_31J40_124_1870_n802), .A3(alu_io_in1[35]), .A4(alu_in2_inv_35_), .Y(alu_DP_OP_31J40_124_1870_n805) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U697 ( .A(alu_io_in1[36]), .B(
        alu_in2_inv_36_), .CI(alu_DP_OP_31J40_124_1870_n805), .S(
        io_dmem_req_bits_addr[36]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U696 ( .A1(alu_io_in1[36]), .A2(
        alu_in2_inv_36_), .A3(alu_io_in1[35]), .A4(alu_in2_inv_35_), .Y(
        alu_DP_OP_31J40_124_1870_n799) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U695 ( .A1(alu_io_in1[36]), .A2(
        alu_in2_inv_36_), .Y(alu_DP_OP_31J40_124_1870_n804) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U694 ( .A1(alu_io_in1[36]), .A2(
        alu_in2_inv_36_), .A3(alu_DP_OP_31J40_124_1870_n803), .A4(
        alu_DP_OP_31J40_124_1870_n804), .Y(alu_DP_OP_31J40_124_1870_n792) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U693 ( .A1(alu_DP_OP_31J40_124_1870_n799), .A2(alu_DP_OP_31J40_124_1870_n802), .A3(alu_DP_OP_31J40_124_1870_n792), .Y(
        alu_DP_OP_31J40_124_1870_n801) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U692 ( .A(alu_io_in1[37]), .B(
        alu_in2_inv_37_), .CI(alu_DP_OP_31J40_124_1870_n801), .S(
        io_dmem_req_bits_addr[37]) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U691 ( .A1(alu_io_in1[37]), .A2(
        alu_in2_inv_37_), .Y(alu_DP_OP_31J40_124_1870_n796) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U690 ( .A1(alu_DP_OP_31J40_124_1870_n796), .A2(alu_DP_OP_31J40_124_1870_n801), .A3(alu_io_in1[37]), .A4(alu_in2_inv_37_), .Y(alu_DP_OP_31J40_124_1870_n800) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U689 ( .A(alu_io_in1[38]), .B(
        alu_in2_inv_38_), .CI(alu_DP_OP_31J40_124_1870_n800), .S(
        io_dmem_req_bits_addr[38]) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U688 ( .A1(alu_io_in1[38]), .A2(
        alu_in2_inv_38_), .A3(alu_io_in1[37]), .A4(alu_in2_inv_37_), .Y(
        alu_DP_OP_31J40_124_1870_n791) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U687 ( .A1(alu_DP_OP_31J40_124_1870_n791), .A2(alu_DP_OP_31J40_124_1870_n799), .Y(alu_DP_OP_31J40_124_1870_n794) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U686 ( .A1(alu_DP_OP_31J40_124_1870_n794), .A2(alu_DP_OP_31J40_124_1870_n798), .Y(alu_DP_OP_31J40_124_1870_n773) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U685 ( .A1(alu_in2_inv_38_), .A2(
        alu_io_in1[38]), .Y(alu_DP_OP_31J40_124_1870_n797) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U684 ( .A1(alu_io_in1[38]), .A2(
        alu_in2_inv_38_), .A3(alu_DP_OP_31J40_124_1870_n796), .A4(
        alu_DP_OP_31J40_124_1870_n797), .Y(alu_DP_OP_31J40_124_1870_n795) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U683 ( .A1(
        alu_DP_OP_31J40_124_1870_n791), .A2(alu_DP_OP_31J40_124_1870_n792), 
        .A3(alu_DP_OP_31J40_124_1870_n793), .A4(alu_DP_OP_31J40_124_1870_n794), 
        .A5(alu_DP_OP_31J40_124_1870_n795), .Y(alu_DP_OP_31J40_124_1870_n767)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U682 ( .A1(alu_DP_OP_31J40_124_1870_n773), .A2(alu_DP_OP_31J40_124_1870_n708), .A3(alu_DP_OP_31J40_124_1870_n767), .Y(
        alu_DP_OP_31J40_124_1870_n781) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U681 ( .A(alu_io_in1[39]), .B(
        alu_in2_inv_39_), .CI(alu_DP_OP_31J40_124_1870_n781), .S(
        alu_io_adder_out_39_) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U680 ( .A1(alu_io_in1[39]), .A2(
        alu_in2_inv_39_), .Y(alu_DP_OP_31J40_124_1870_n789) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U679 ( .A1(alu_DP_OP_31J40_124_1870_n789), .A2(alu_DP_OP_31J40_124_1870_n781), .A3(alu_io_in1[39]), .A4(alu_in2_inv_39_), .Y(alu_DP_OP_31J40_124_1870_n790) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U678 ( .A(alu_io_in1[40]), .B(
        alu_in2_inv_40_), .CI(alu_DP_OP_31J40_124_1870_n790), .S(alu_n630) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U677 ( .A1(alu_io_in1[40]), .A2(
        alu_in2_inv_40_), .A3(alu_io_in1[39]), .A4(alu_in2_inv_39_), .Y(
        alu_DP_OP_31J40_124_1870_n786) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U676 ( .A1(alu_DP_OP_31J40_124_1870_n786), .A2(alu_DP_OP_31J40_124_1870_n781), .A3(alu_DP_OP_31J40_124_1870_n785), .Y(
        alu_DP_OP_31J40_124_1870_n788) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U675 ( .A(alu_io_in1[41]), .B(
        alu_in2_inv_41_), .CI(alu_DP_OP_31J40_124_1870_n788), .S(alu_n629) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U674 ( .A1(alu_io_in1[41]), .A2(
        alu_in2_inv_41_), .Y(alu_DP_OP_31J40_124_1870_n782) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U673 ( .A1(alu_DP_OP_31J40_124_1870_n782), .A2(alu_DP_OP_31J40_124_1870_n788), .A3(alu_io_in1[41]), .A4(alu_in2_inv_41_), .Y(alu_DP_OP_31J40_124_1870_n787) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U672 ( .A(alu_io_in1[42]), .B(
        alu_in2_inv_42_), .CI(alu_DP_OP_31J40_124_1870_n787), .S(alu_n628) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U671 ( .A1(alu_io_in1[42]), .A2(
        alu_in2_inv_42_), .A3(alu_io_in1[41]), .A4(alu_in2_inv_41_), .Y(
        alu_DP_OP_31J40_124_1870_n784) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U670 ( .A1(alu_DP_OP_31J40_124_1870_n784), .A2(alu_DP_OP_31J40_124_1870_n786), .Y(alu_DP_OP_31J40_124_1870_n774) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U669 ( .A1(alu_in2_inv_42_), .A2(
        alu_io_in1[42]), .Y(alu_DP_OP_31J40_124_1870_n783) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U668 ( .A1(alu_io_in1[42]), .A2(
        alu_in2_inv_42_), .A3(alu_DP_OP_31J40_124_1870_n782), .A4(
        alu_DP_OP_31J40_124_1870_n783), .A5(alu_DP_OP_31J40_124_1870_n784), 
        .A6(alu_DP_OP_31J40_124_1870_n785), .Y(alu_DP_OP_31J40_124_1870_n764)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U667 ( .A1(alu_DP_OP_31J40_124_1870_n774), .A2(alu_DP_OP_31J40_124_1870_n781), .A3(alu_DP_OP_31J40_124_1870_n764), .Y(
        alu_DP_OP_31J40_124_1870_n778) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U666 ( .A(alu_io_in1[43]), .B(
        alu_in2_inv_43_), .CI(alu_DP_OP_31J40_124_1870_n778), .S(alu_n627) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U665 ( .A1(alu_io_in1[43]), .A2(
        alu_in2_inv_43_), .Y(alu_DP_OP_31J40_124_1870_n779) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U664 ( .A1(alu_DP_OP_31J40_124_1870_n779), .A2(alu_DP_OP_31J40_124_1870_n778), .A3(alu_io_in1[43]), .A4(alu_in2_inv_43_), .Y(alu_DP_OP_31J40_124_1870_n780) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U663 ( .A(alu_io_in1[44]), .B(
        alu_in2_inv_44_), .CI(alu_DP_OP_31J40_124_1870_n780), .S(alu_n626) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U662 ( .A1(alu_io_in1[44]), .A2(
        alu_in2_inv_44_), .A3(alu_io_in1[43]), .A4(alu_in2_inv_43_), .Y(
        alu_DP_OP_31J40_124_1870_n775) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U661 ( .A1(alu_DP_OP_31J40_124_1870_n775), .A2(alu_DP_OP_31J40_124_1870_n778), .A3(alu_DP_OP_31J40_124_1870_n772), .Y(
        alu_DP_OP_31J40_124_1870_n777) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U660 ( .A(alu_io_in1[45]), .B(
        alu_in2_inv_45_), .CI(alu_DP_OP_31J40_124_1870_n777), .S(alu_n625) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U659 ( .A1(alu_io_in1[45]), .A2(
        alu_in2_inv_45_), .Y(alu_DP_OP_31J40_124_1870_n769) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U658 ( .A1(alu_DP_OP_31J40_124_1870_n769), .A2(alu_DP_OP_31J40_124_1870_n777), .A3(alu_io_in1[45]), .A4(alu_in2_inv_45_), .Y(alu_DP_OP_31J40_124_1870_n776) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U657 ( .A(alu_io_in1[46]), .B(
        alu_in2_inv_46_), .CI(alu_DP_OP_31J40_124_1870_n776), .S(alu_n624) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U656 ( .A1(alu_io_in1[46]), .A2(
        alu_in2_inv_46_), .A3(alu_io_in1[45]), .A4(alu_in2_inv_45_), .Y(
        alu_DP_OP_31J40_124_1870_n771) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U655 ( .A1(alu_DP_OP_31J40_124_1870_n771), .A2(alu_DP_OP_31J40_124_1870_n775), .Y(alu_DP_OP_31J40_124_1870_n765) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U654 ( .A1(alu_DP_OP_31J40_124_1870_n774), .A2(alu_DP_OP_31J40_124_1870_n765), .Y(alu_DP_OP_31J40_124_1870_n766) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U653 ( .A1(alu_DP_OP_31J40_124_1870_n766), .A2(alu_DP_OP_31J40_124_1870_n773), .Y(alu_DP_OP_31J40_124_1870_n706) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U652 ( .A1(alu_in2_inv_46_), .A2(
        alu_io_in1[46]), .Y(alu_DP_OP_31J40_124_1870_n770) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U651 ( .A1(alu_io_in1[46]), .A2(
        alu_in2_inv_46_), .A3(alu_DP_OP_31J40_124_1870_n769), .A4(
        alu_DP_OP_31J40_124_1870_n770), .A5(alu_DP_OP_31J40_124_1870_n771), 
        .A6(alu_DP_OP_31J40_124_1870_n772), .Y(alu_DP_OP_31J40_124_1870_n768)
         );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U650 ( .A1(
        alu_DP_OP_31J40_124_1870_n764), .A2(alu_DP_OP_31J40_124_1870_n765), 
        .A3(alu_DP_OP_31J40_124_1870_n766), .A4(alu_DP_OP_31J40_124_1870_n767), 
        .A5(alu_DP_OP_31J40_124_1870_n768), .Y(alu_DP_OP_31J40_124_1870_n709)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U649 ( .A1(alu_DP_OP_31J40_124_1870_n706), .A2(alu_DP_OP_31J40_124_1870_n708), .A3(alu_DP_OP_31J40_124_1870_n709), .Y(
        alu_DP_OP_31J40_124_1870_n739) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U648 ( .A(alu_io_in1[47]), .B(
        alu_in2_inv_47_), .CI(alu_DP_OP_31J40_124_1870_n739), .S(alu_n623) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U647 ( .A1(alu_io_in1[47]), .A2(
        alu_in2_inv_47_), .Y(alu_DP_OP_31J40_124_1870_n761) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U646 ( .A1(alu_DP_OP_31J40_124_1870_n761), .A2(alu_DP_OP_31J40_124_1870_n739), .A3(alu_io_in1[47]), .A4(alu_in2_inv_47_), .Y(alu_DP_OP_31J40_124_1870_n763) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U645 ( .A(alu_io_in1[48]), .B(
        alu_in2_inv_48_), .CI(alu_DP_OP_31J40_124_1870_n763), .S(alu_n622) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U644 ( .A1(alu_io_in1[48]), .A2(
        alu_in2_inv_48_), .A3(alu_io_in1[47]), .A4(alu_in2_inv_47_), .Y(
        alu_DP_OP_31J40_124_1870_n758) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U643 ( .A1(alu_io_in1[48]), .A2(
        alu_in2_inv_48_), .Y(alu_DP_OP_31J40_124_1870_n762) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U642 ( .A1(alu_io_in1[48]), .A2(
        alu_in2_inv_48_), .A3(alu_DP_OP_31J40_124_1870_n761), .A4(
        alu_DP_OP_31J40_124_1870_n762), .Y(alu_DP_OP_31J40_124_1870_n757) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U641 ( .A1(alu_DP_OP_31J40_124_1870_n758), .A2(alu_DP_OP_31J40_124_1870_n739), .A3(alu_DP_OP_31J40_124_1870_n757), .Y(
        alu_DP_OP_31J40_124_1870_n760) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U640 ( .A(alu_io_in1[49]), .B(
        alu_in2_inv_49_), .CI(alu_DP_OP_31J40_124_1870_n760), .S(alu_n621) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U639 ( .A1(alu_io_in1[49]), .A2(
        alu_in2_inv_49_), .Y(alu_DP_OP_31J40_124_1870_n754) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U638 ( .A1(alu_DP_OP_31J40_124_1870_n754), .A2(alu_DP_OP_31J40_124_1870_n760), .A3(alu_io_in1[49]), .A4(alu_in2_inv_49_), .Y(alu_DP_OP_31J40_124_1870_n759) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U637 ( .A(alu_io_in1[50]), .B(
        alu_in2_inv_50_), .CI(alu_DP_OP_31J40_124_1870_n759), .S(alu_n620) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U636 ( .A1(alu_io_in1[50]), .A2(
        alu_in2_inv_50_), .A3(alu_io_in1[49]), .A4(alu_in2_inv_49_), .Y(
        alu_DP_OP_31J40_124_1870_n756) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U635 ( .A1(alu_DP_OP_31J40_124_1870_n756), .A2(alu_DP_OP_31J40_124_1870_n758), .Y(alu_DP_OP_31J40_124_1870_n747) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U634 ( .A1(alu_in2_inv_50_), .A2(
        alu_io_in1[50]), .Y(alu_DP_OP_31J40_124_1870_n755) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U633 ( .A1(alu_io_in1[50]), .A2(
        alu_in2_inv_50_), .A3(alu_DP_OP_31J40_124_1870_n754), .A4(
        alu_DP_OP_31J40_124_1870_n755), .A5(alu_DP_OP_31J40_124_1870_n756), 
        .A6(alu_DP_OP_31J40_124_1870_n757), .Y(alu_DP_OP_31J40_124_1870_n742)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U632 ( .A1(alu_DP_OP_31J40_124_1870_n747), .A2(alu_DP_OP_31J40_124_1870_n739), .A3(alu_DP_OP_31J40_124_1870_n742), .Y(
        alu_DP_OP_31J40_124_1870_n751) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U631 ( .A(alu_io_in1[51]), .B(
        alu_in2_inv_51_), .CI(alu_DP_OP_31J40_124_1870_n751), .S(alu_n619) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U630 ( .A1(alu_io_in1[51]), .A2(
        alu_in2_inv_51_), .Y(alu_DP_OP_31J40_124_1870_n752) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U629 ( .A1(alu_DP_OP_31J40_124_1870_n752), .A2(alu_DP_OP_31J40_124_1870_n751), .A3(alu_io_in1[51]), .A4(alu_in2_inv_51_), .Y(alu_DP_OP_31J40_124_1870_n753) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U628 ( .A(alu_io_in1[52]), .B(
        alu_in2_inv_52_), .CI(alu_DP_OP_31J40_124_1870_n753), .S(alu_n618) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U627 ( .A1(alu_io_in1[52]), .A2(
        alu_in2_inv_52_), .A3(alu_io_in1[51]), .A4(alu_in2_inv_51_), .Y(
        alu_DP_OP_31J40_124_1870_n748) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U626 ( .A1(alu_DP_OP_31J40_124_1870_n748), .A2(alu_DP_OP_31J40_124_1870_n751), .A3(alu_DP_OP_31J40_124_1870_n741), .Y(
        alu_DP_OP_31J40_124_1870_n750) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U625 ( .A(alu_io_in1[53]), .B(
        alu_in2_inv_53_), .CI(alu_DP_OP_31J40_124_1870_n750), .S(alu_n617) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U624 ( .A1(alu_io_in1[53]), .A2(
        alu_in2_inv_53_), .Y(alu_DP_OP_31J40_124_1870_n745) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U623 ( .A1(alu_DP_OP_31J40_124_1870_n745), .A2(alu_DP_OP_31J40_124_1870_n750), .A3(alu_io_in1[53]), .A4(alu_in2_inv_53_), .Y(alu_DP_OP_31J40_124_1870_n749) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U622 ( .A(alu_io_in1[54]), .B(
        alu_in2_inv_54_), .CI(alu_DP_OP_31J40_124_1870_n749), .S(alu_n616) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U621 ( .A1(alu_io_in1[54]), .A2(
        alu_in2_inv_54_), .A3(alu_io_in1[53]), .A4(alu_in2_inv_53_), .Y(
        alu_DP_OP_31J40_124_1870_n740) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U620 ( .A1(alu_DP_OP_31J40_124_1870_n740), .A2(alu_DP_OP_31J40_124_1870_n748), .Y(alu_DP_OP_31J40_124_1870_n743) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U619 ( .A1(alu_DP_OP_31J40_124_1870_n743), .A2(alu_DP_OP_31J40_124_1870_n747), .Y(alu_DP_OP_31J40_124_1870_n723) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U618 ( .A1(alu_in2_inv_54_), .A2(
        alu_io_in1[54]), .Y(alu_DP_OP_31J40_124_1870_n746) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U617 ( .A1(alu_io_in1[54]), .A2(
        alu_in2_inv_54_), .A3(alu_DP_OP_31J40_124_1870_n745), .A4(
        alu_DP_OP_31J40_124_1870_n746), .Y(alu_DP_OP_31J40_124_1870_n744) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U616 ( .A1(
        alu_DP_OP_31J40_124_1870_n740), .A2(alu_DP_OP_31J40_124_1870_n741), 
        .A3(alu_DP_OP_31J40_124_1870_n742), .A4(alu_DP_OP_31J40_124_1870_n743), 
        .A5(alu_DP_OP_31J40_124_1870_n744), .Y(alu_DP_OP_31J40_124_1870_n711)
         );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U615 ( .A1(alu_DP_OP_31J40_124_1870_n723), .A2(alu_DP_OP_31J40_124_1870_n739), .A3(alu_DP_OP_31J40_124_1870_n711), .Y(
        alu_DP_OP_31J40_124_1870_n730) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U614 ( .A(alu_io_in1[55]), .B(
        alu_in2_inv_55_), .CI(alu_DP_OP_31J40_124_1870_n730), .S(alu_n615) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U613 ( .A1(alu_io_in1[55]), .A2(
        alu_in2_inv_55_), .Y(alu_DP_OP_31J40_124_1870_n737) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U612 ( .A1(alu_DP_OP_31J40_124_1870_n737), .A2(alu_DP_OP_31J40_124_1870_n730), .A3(alu_io_in1[55]), .A4(alu_in2_inv_55_), .Y(alu_DP_OP_31J40_124_1870_n738) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U611 ( .A(alu_io_in1[56]), .B(
        alu_in2_inv_56_), .CI(alu_DP_OP_31J40_124_1870_n738), .S(alu_n614) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U610 ( .A1(alu_io_in1[56]), .A2(
        alu_in2_inv_56_), .A3(alu_io_in1[55]), .A4(alu_in2_inv_55_), .Y(
        alu_DP_OP_31J40_124_1870_n734) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U609 ( .A1(alu_DP_OP_31J40_124_1870_n734), .A2(alu_DP_OP_31J40_124_1870_n730), .A3(alu_DP_OP_31J40_124_1870_n733), .Y(
        alu_DP_OP_31J40_124_1870_n736) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U608 ( .A(alu_io_in1[57]), .B(
        alu_in2_inv_57_), .CI(alu_DP_OP_31J40_124_1870_n736), .S(alu_n613) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U607 ( .A1(alu_io_in1[57]), .A2(
        alu_in2_inv_57_), .Y(alu_DP_OP_31J40_124_1870_n731) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U606 ( .A1(alu_DP_OP_31J40_124_1870_n731), .A2(alu_DP_OP_31J40_124_1870_n736), .A3(alu_io_in1[57]), .A4(alu_in2_inv_57_), .Y(alu_DP_OP_31J40_124_1870_n735) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U605 ( .A(alu_io_in1[58]), .B(
        alu_in2_inv_58_), .CI(alu_DP_OP_31J40_124_1870_n735), .S(alu_n612) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U604 ( .A1(alu_io_in1[58]), .A2(
        alu_in2_inv_58_), .A3(alu_io_in1[57]), .A4(alu_in2_inv_57_), .Y(
        alu_DP_OP_31J40_124_1870_n732) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U603 ( .A1(alu_DP_OP_31J40_124_1870_n732), .A2(alu_DP_OP_31J40_124_1870_n734), .Y(alu_DP_OP_31J40_124_1870_n724) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U602 ( .A1(alu_DP_OP_31J40_124_1870_n724), .A2(alu_DP_OP_31J40_124_1870_n730), .A3(alu_DP_OP_31J40_124_1870_n720), .Y(
        alu_DP_OP_31J40_124_1870_n727) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U601 ( .A(alu_io_in1[59]), .B(
        alu_in2_inv_59_), .CI(alu_DP_OP_31J40_124_1870_n727), .S(alu_n611) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U600 ( .A1(alu_io_in1[59]), .A2(
        alu_in2_inv_59_), .Y(alu_DP_OP_31J40_124_1870_n728) );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U599 ( .A1(
        alu_DP_OP_31J40_124_1870_n727), .A2(alu_io_in1[59]), .A3(
        alu_DP_OP_31J40_124_1870_n727), .A4(alu_in2_inv_59_), .A5(
        alu_DP_OP_31J40_124_1870_n728), .Y(alu_DP_OP_31J40_124_1870_n729) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U598 ( .A(alu_io_in1[60]), .B(
        alu_in2_inv_60_), .CI(alu_DP_OP_31J40_124_1870_n729), .S(alu_n610) );
  OA22X1_LVT alu_DP_OP_31J40_124_1870_U597 ( .A1(alu_io_in1[60]), .A2(
        alu_in2_inv_60_), .A3(alu_io_in1[59]), .A4(alu_in2_inv_59_), .Y(
        alu_DP_OP_31J40_124_1870_n719) );
  AO21X1_LVT alu_DP_OP_31J40_124_1870_U596 ( .A1(alu_DP_OP_31J40_124_1870_n719), .A2(alu_DP_OP_31J40_124_1870_n727), .A3(alu_DP_OP_31J40_124_1870_n718), .Y(
        alu_DP_OP_31J40_124_1870_n726) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U595 ( .A(alu_io_in1[61]), .B(
        alu_in2_inv_61_), .CI(alu_DP_OP_31J40_124_1870_n726), .S(alu_n609) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U594 ( .A1(alu_io_in1[61]), .A2(
        alu_in2_inv_61_), .Y(alu_DP_OP_31J40_124_1870_n716) );
  AO22X1_LVT alu_DP_OP_31J40_124_1870_U593 ( .A1(alu_io_in1[61]), .A2(
        alu_in2_inv_61_), .A3(alu_DP_OP_31J40_124_1870_n726), .A4(
        alu_DP_OP_31J40_124_1870_n716), .Y(alu_DP_OP_31J40_124_1870_n725) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U592 ( .A(alu_io_in1[62]), .B(
        alu_in2_inv_62_), .CI(alu_DP_OP_31J40_124_1870_n725), .S(alu_n608) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U591 ( .A1(alu_io_in1[62]), .A2(
        alu_in2_inv_62_), .Y(alu_DP_OP_31J40_124_1870_n717) );
  AND4X1_LVT alu_DP_OP_31J40_124_1870_U590 ( .A1(alu_DP_OP_31J40_124_1870_n719), .A2(alu_DP_OP_31J40_124_1870_n724), .A3(alu_DP_OP_31J40_124_1870_n716), .A4(
        alu_DP_OP_31J40_124_1870_n717), .Y(alu_DP_OP_31J40_124_1870_n710) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U589 ( .A1(alu_DP_OP_31J40_124_1870_n723), .A2(alu_DP_OP_31J40_124_1870_n710), .Y(alu_DP_OP_31J40_124_1870_n707) );
  NAND2X0_LVT alu_DP_OP_31J40_124_1870_U588 ( .A1(alu_io_in1[62]), .A2(
        alu_in2_inv_62_), .Y(alu_DP_OP_31J40_124_1870_n721) );
  NAND3X0_LVT alu_DP_OP_31J40_124_1870_U587 ( .A1(alu_io_in1[61]), .A2(
        alu_in2_inv_61_), .A3(alu_DP_OP_31J40_124_1870_n717), .Y(
        alu_DP_OP_31J40_124_1870_n722) );
  NAND4X0_LVT alu_DP_OP_31J40_124_1870_U586 ( .A1(
        alu_DP_OP_31J40_124_1870_n719), .A2(alu_DP_OP_31J40_124_1870_n720), 
        .A3(alu_DP_OP_31J40_124_1870_n716), .A4(alu_DP_OP_31J40_124_1870_n717), 
        .Y(alu_DP_OP_31J40_124_1870_n714) );
  NAND3X0_LVT alu_DP_OP_31J40_124_1870_U585 ( .A1(
        alu_DP_OP_31J40_124_1870_n716), .A2(alu_DP_OP_31J40_124_1870_n717), 
        .A3(alu_DP_OP_31J40_124_1870_n718), .Y(alu_DP_OP_31J40_124_1870_n715)
         );
  NAND3X0_LVT alu_DP_OP_31J40_124_1870_U584 ( .A1(
        alu_DP_OP_31J40_124_1870_n713), .A2(alu_DP_OP_31J40_124_1870_n714), 
        .A3(alu_DP_OP_31J40_124_1870_n715), .Y(alu_DP_OP_31J40_124_1870_n712)
         );
  AO221X1_LVT alu_DP_OP_31J40_124_1870_U583 ( .A1(
        alu_DP_OP_31J40_124_1870_n709), .A2(alu_DP_OP_31J40_124_1870_n707), 
        .A3(alu_DP_OP_31J40_124_1870_n710), .A4(alu_DP_OP_31J40_124_1870_n711), 
        .A5(alu_DP_OP_31J40_124_1870_n712), .Y(alu_DP_OP_31J40_124_1870_n705)
         );
  OA222X1_LVT alu_DP_OP_31J40_124_1870_U582 ( .A1(
        alu_DP_OP_31J40_124_1870_n705), .A2(alu_DP_OP_31J40_124_1870_n706), 
        .A3(alu_DP_OP_31J40_124_1870_n705), .A4(alu_DP_OP_31J40_124_1870_n707), 
        .A5(alu_DP_OP_31J40_124_1870_n705), .A6(alu_DP_OP_31J40_124_1870_n708), 
        .Y(alu_DP_OP_31J40_124_1870_n704) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U581 ( .A(alu_DP_OP_31J40_124_1870_n704), 
        .B(alu_io_in1[63]), .CI(alu_in2_inv_63_), .S(alu_n607) );
  AND2X1_LVT alu_DP_OP_31J40_124_1870_U580 ( .A1(alu_DP_OP_31J40_124_1870_n721), .A2(alu_DP_OP_31J40_124_1870_n722), .Y(alu_DP_OP_31J40_124_1870_n713) );
  OA222X1_LVT alu_DP_OP_31J40_124_1870_U579 ( .A1(
        alu_DP_OP_31J40_124_1870_n913), .A2(alu_DP_OP_31J40_124_1870_n442), 
        .A3(alu_DP_OP_31J40_124_1870_n913), .A4(alu_DP_OP_31J40_124_1870_n914), 
        .A5(alu_DP_OP_31J40_124_1870_n913), .A6(alu_DP_OP_31J40_124_1870_n915), 
        .Y(alu_DP_OP_31J40_124_1870_n906) );
  OA222X1_LVT alu_DP_OP_31J40_124_1870_U578 ( .A1(
        alu_DP_OP_31J40_124_1870_n873), .A2(alu_DP_OP_31J40_124_1870_n874), 
        .A3(alu_DP_OP_31J40_124_1870_n873), .A4(alu_DP_OP_31J40_124_1870_n875), 
        .A5(alu_DP_OP_31J40_124_1870_n873), .A6(alu_DP_OP_31J40_124_1870_n876), 
        .Y(alu_DP_OP_31J40_124_1870_n827) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U577 ( .A1(alu_io_in1[56]), .A2(
        alu_in2_inv_56_), .A3(alu_io_in1[56]), .A4(
        alu_DP_OP_31J40_124_1870_n737), .A5(alu_in2_inv_56_), .A6(
        alu_DP_OP_31J40_124_1870_n737), .Y(alu_DP_OP_31J40_124_1870_n733) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U576 ( .A1(alu_io_in1[60]), .A2(
        alu_in2_inv_60_), .A3(alu_io_in1[60]), .A4(
        alu_DP_OP_31J40_124_1870_n728), .A5(alu_in2_inv_60_), .A6(
        alu_DP_OP_31J40_124_1870_n728), .Y(alu_DP_OP_31J40_124_1870_n718) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U575 ( .A1(alu_io_in1[44]), .A2(
        alu_in2_inv_44_), .A3(alu_io_in1[44]), .A4(
        alu_DP_OP_31J40_124_1870_n779), .A5(alu_in2_inv_44_), .A6(
        alu_DP_OP_31J40_124_1870_n779), .Y(alu_DP_OP_31J40_124_1870_n772) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U574 ( .A1(alu_io_in1[40]), .A2(
        alu_in2_inv_40_), .A3(alu_io_in1[40]), .A4(
        alu_DP_OP_31J40_124_1870_n789), .A5(alu_in2_inv_40_), .A6(
        alu_DP_OP_31J40_124_1870_n789), .Y(alu_DP_OP_31J40_124_1870_n785) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U573 ( .A1(
        alu_DP_OP_31J40_124_1870_n703), .A2(alu_DP_OP_31J40_124_1870_n731), 
        .A3(alu_DP_OP_31J40_124_1870_n733), .A4(alu_DP_OP_31J40_124_1870_n732), 
        .A5(alu_io_in1[58]), .A6(alu_in2_inv_58_), .Y(
        alu_DP_OP_31J40_124_1870_n720) );
  OR2X1_LVT alu_DP_OP_31J40_124_1870_U572 ( .A1(alu_io_in1[58]), .A2(
        alu_in2_inv_58_), .Y(alu_DP_OP_31J40_124_1870_n703) );
  AO222X1_LVT alu_DP_OP_31J40_124_1870_U571 ( .A1(alu_io_in1[52]), .A2(
        alu_in2_inv_52_), .A3(alu_io_in1[52]), .A4(
        alu_DP_OP_31J40_124_1870_n752), .A5(alu_in2_inv_52_), .A6(
        alu_DP_OP_31J40_124_1870_n752), .Y(alu_DP_OP_31J40_124_1870_n741) );
  FADDX1_LVT alu_DP_OP_31J40_124_1870_U568 ( .A(alu_io_in1[0]), .B(
        alu_in2_inv_0_), .CI(alu_io_fn[3]), .CO(alu_DP_OP_31J40_124_1870_n442), 
        .S(io_dmem_req_bits_addr[0]) );
  AO22X1_LVT alu_ashr_7_U830 ( .A1(alu_ashr_7_n502), .A2(alu_shin_63_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_62_), .Y(alu_ashr_7_n836) );
  AO22X1_LVT alu_ashr_7_U829 ( .A1(alu_ashr_7_n502), .A2(alu_shin_61_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_60_), .Y(alu_ashr_7_n834) );
  AO22X1_LVT alu_ashr_7_U828 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n836), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n834), .Y(alu_ashr_7_n805) );
  AO22X1_LVT alu_ashr_7_U827 ( .A1(alu_ashr_7_n502), .A2(alu_shin_59_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_58_), .Y(alu_ashr_7_n835) );
  AO22X1_LVT alu_ashr_7_U826 ( .A1(alu_ashr_7_n502), .A2(alu_shin_57_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_56_), .Y(alu_ashr_7_n832) );
  AO22X1_LVT alu_ashr_7_U825 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n835), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n832), .Y(alu_ashr_7_n803) );
  AO22X1_LVT alu_ashr_7_U824 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n805), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n803), .Y(alu_ashr_7_n663) );
  AO22X1_LVT alu_ashr_7_U823 ( .A1(alu_ashr_7_n502), .A2(alu_shin_55_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_54_), .Y(alu_ashr_7_n833) );
  AO22X1_LVT alu_ashr_7_U822 ( .A1(alu_ashr_7_n502), .A2(alu_shin_53_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_52_), .Y(alu_ashr_7_n830) );
  AO22X1_LVT alu_ashr_7_U821 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n833), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n830), .Y(alu_ashr_7_n804) );
  AO22X1_LVT alu_ashr_7_U820 ( .A1(alu_ashr_7_n502), .A2(alu_shin_51_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_50_), .Y(alu_ashr_7_n831) );
  AO22X1_LVT alu_ashr_7_U819 ( .A1(alu_ashr_7_n502), .A2(alu_shin_49_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_48_), .Y(alu_ashr_7_n828) );
  AO22X1_LVT alu_ashr_7_U818 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n831), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n828), .Y(alu_ashr_7_n801) );
  AO22X1_LVT alu_ashr_7_U817 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n804), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n801), .Y(alu_ashr_7_n661) );
  AO22X1_LVT alu_ashr_7_U816 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n663), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n661), .Y(alu_ashr_7_n732) );
  AO22X1_LVT alu_ashr_7_U815 ( .A1(alu_ashr_7_n502), .A2(alu_shin_47_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_46_), .Y(alu_ashr_7_n829) );
  AO22X1_LVT alu_ashr_7_U814 ( .A1(alu_ashr_7_n502), .A2(alu_shin_45_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_44_), .Y(alu_ashr_7_n826) );
  AO22X1_LVT alu_ashr_7_U813 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n829), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n826), .Y(alu_ashr_7_n802) );
  AO22X1_LVT alu_ashr_7_U812 ( .A1(alu_ashr_7_n502), .A2(alu_shin_43_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_42_), .Y(alu_ashr_7_n827) );
  AO22X1_LVT alu_ashr_7_U811 ( .A1(alu_ashr_7_n502), .A2(alu_shin_41_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_40_), .Y(alu_ashr_7_n824) );
  AO22X1_LVT alu_ashr_7_U810 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n827), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n824), .Y(alu_ashr_7_n799) );
  AO22X1_LVT alu_ashr_7_U809 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n802), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n799), .Y(alu_ashr_7_n662) );
  AO22X1_LVT alu_ashr_7_U808 ( .A1(alu_ashr_7_n502), .A2(alu_shin_39_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_38_), .Y(alu_ashr_7_n825) );
  AO22X1_LVT alu_ashr_7_U807 ( .A1(alu_ashr_7_n502), .A2(alu_shin_37_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_36_), .Y(alu_ashr_7_n822) );
  AO22X1_LVT alu_ashr_7_U806 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n825), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n822), .Y(alu_ashr_7_n800) );
  AO22X1_LVT alu_ashr_7_U805 ( .A1(alu_ashr_7_n502), .A2(alu_shin_35_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_34_), .Y(alu_ashr_7_n823) );
  AO22X1_LVT alu_ashr_7_U804 ( .A1(alu_ashr_7_n502), .A2(alu_shin_33_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_32_), .Y(alu_ashr_7_n820) );
  AO22X1_LVT alu_ashr_7_U803 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n823), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n820), .Y(alu_ashr_7_n797) );
  AO22X1_LVT alu_ashr_7_U802 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n800), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n797), .Y(alu_ashr_7_n659) );
  AO22X1_LVT alu_ashr_7_U801 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n662), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n659), .Y(alu_ashr_7_n730) );
  AO22X1_LVT alu_ashr_7_U800 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n732), 
        .A3(alu_ashr_7_n521), .A4(alu_ashr_7_n730), .Y(alu_ashr_7_n615) );
  AO22X1_LVT alu_ashr_7_U799 ( .A1(alu_ashr_7_n502), .A2(alu_shin_31_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_30_), .Y(alu_ashr_7_n821) );
  AO22X1_LVT alu_ashr_7_U798 ( .A1(alu_ashr_7_n502), .A2(alu_shin_29_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_28_), .Y(alu_ashr_7_n818) );
  AO22X1_LVT alu_ashr_7_U797 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n821), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n818), .Y(alu_ashr_7_n798) );
  AO22X1_LVT alu_ashr_7_U796 ( .A1(alu_ashr_7_n502), .A2(alu_shin_27_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_26_), .Y(alu_ashr_7_n819) );
  AO22X1_LVT alu_ashr_7_U795 ( .A1(alu_ashr_7_n502), .A2(alu_shin_25_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_24_), .Y(alu_ashr_7_n816) );
  AO22X1_LVT alu_ashr_7_U794 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n819), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n816), .Y(alu_ashr_7_n795) );
  AO22X1_LVT alu_ashr_7_U793 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n798), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n795), .Y(alu_ashr_7_n660) );
  AO22X1_LVT alu_ashr_7_U792 ( .A1(alu_ashr_7_n502), .A2(alu_shin_23_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_22_), .Y(alu_ashr_7_n817) );
  AO22X1_LVT alu_ashr_7_U791 ( .A1(alu_ashr_7_n502), .A2(alu_shin_21_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_20_), .Y(alu_ashr_7_n814) );
  AO22X1_LVT alu_ashr_7_U790 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n817), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n814), .Y(alu_ashr_7_n796) );
  AO22X1_LVT alu_ashr_7_U789 ( .A1(alu_ashr_7_n502), .A2(alu_shin_19_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_18_), .Y(alu_ashr_7_n815) );
  AO22X1_LVT alu_ashr_7_U788 ( .A1(alu_ashr_7_n502), .A2(alu_shin_17_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_16_), .Y(alu_ashr_7_n812) );
  AO22X1_LVT alu_ashr_7_U787 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n815), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n812), .Y(alu_ashr_7_n793) );
  AO22X1_LVT alu_ashr_7_U786 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n796), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n793), .Y(alu_ashr_7_n532) );
  AO22X1_LVT alu_ashr_7_U785 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n660), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n532), .Y(alu_ashr_7_n731) );
  AO22X1_LVT alu_ashr_7_U784 ( .A1(alu_ashr_7_n502), .A2(alu_shin_15_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_14_), .Y(alu_ashr_7_n813) );
  AO22X1_LVT alu_ashr_7_U783 ( .A1(alu_ashr_7_n502), .A2(alu_shin_13_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_12_), .Y(alu_ashr_7_n810) );
  AO22X1_LVT alu_ashr_7_U782 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n813), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n810), .Y(alu_ashr_7_n794) );
  AO22X1_LVT alu_ashr_7_U781 ( .A1(alu_ashr_7_n502), .A2(alu_shin_11_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_10_), .Y(alu_ashr_7_n811) );
  AO22X1_LVT alu_ashr_7_U780 ( .A1(alu_ashr_7_n502), .A2(alu_shin_9_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_8_), .Y(alu_ashr_7_n632) );
  AO22X1_LVT alu_ashr_7_U779 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n811), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n632), .Y(alu_ashr_7_n578) );
  AO22X1_LVT alu_ashr_7_U778 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n794), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n578), .Y(alu_ashr_7_n533) );
  AO22X1_LVT alu_ashr_7_U777 ( .A1(alu_ashr_7_n502), .A2(alu_shin_7_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_6_), .Y(alu_ashr_7_n633) );
  AO22X1_LVT alu_ashr_7_U776 ( .A1(alu_ashr_7_n502), .A2(alu_shin_5_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_4_), .Y(alu_ashr_7_n630) );
  AO22X1_LVT alu_ashr_7_U775 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n633), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n630), .Y(alu_ashr_7_n579) );
  AO22X1_LVT alu_ashr_7_U774 ( .A1(alu_ashr_7_n502), .A2(alu_shin_3_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_2_), .Y(alu_ashr_7_n631) );
  AO22X1_LVT alu_ashr_7_U773 ( .A1(alu_ashr_7_n502), .A2(alu_shin_1_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_0_), .Y(alu_ashr_7_n841) );
  AO22X1_LVT alu_ashr_7_U772 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n631), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n841), .Y(alu_ashr_7_n840) );
  AO22X1_LVT alu_ashr_7_U771 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n579), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n840), .Y(alu_ashr_7_n839) );
  AO22X1_LVT alu_ashr_7_U770 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n533), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n839), .Y(alu_ashr_7_n838) );
  AO22X1_LVT alu_ashr_7_U769 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n731), 
        .A3(alu_ashr_7_n521), .A4(alu_ashr_7_n838), .Y(alu_ashr_7_n837) );
  AO22X1_LVT alu_ashr_7_U768 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n615), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n837), .Y(alu_n_T_101_0_) );
  AO22X1_LVT alu_ashr_7_U767 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n836), .Y(alu_ashr_7_n762) );
  AO22X1_LVT alu_ashr_7_U766 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n834), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n835), .Y(alu_ashr_7_n760) );
  AO22X1_LVT alu_ashr_7_U765 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n762), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n760), .Y(alu_ashr_7_n714) );
  AO22X1_LVT alu_ashr_7_U764 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n714), .Y(alu_ashr_7_n651) );
  AO22X1_LVT alu_ashr_7_U763 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n832), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n833), .Y(alu_ashr_7_n761) );
  AO22X1_LVT alu_ashr_7_U762 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n830), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n831), .Y(alu_ashr_7_n758) );
  AO22X1_LVT alu_ashr_7_U761 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n761), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n758), .Y(alu_ashr_7_n715) );
  AO22X1_LVT alu_ashr_7_U760 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n828), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n829), .Y(alu_ashr_7_n759) );
  AO22X1_LVT alu_ashr_7_U759 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n826), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n827), .Y(alu_ashr_7_n756) );
  AO22X1_LVT alu_ashr_7_U758 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n759), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n756), .Y(alu_ashr_7_n712) );
  AO22X1_LVT alu_ashr_7_U757 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n715), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n712), .Y(alu_ashr_7_n649) );
  AO22X1_LVT alu_ashr_7_U756 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n651), 
        .A3(alu_ashr_7_n521), .A4(alu_ashr_7_n649), .Y(alu_ashr_7_n587) );
  AO22X1_LVT alu_ashr_7_U755 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n824), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n825), .Y(alu_ashr_7_n757) );
  AO22X1_LVT alu_ashr_7_U754 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n822), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n823), .Y(alu_ashr_7_n754) );
  AO22X1_LVT alu_ashr_7_U753 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n757), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n754), .Y(alu_ashr_7_n713) );
  AO22X1_LVT alu_ashr_7_U752 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n820), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n821), .Y(alu_ashr_7_n755) );
  AO22X1_LVT alu_ashr_7_U751 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n818), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n819), .Y(alu_ashr_7_n752) );
  AO22X1_LVT alu_ashr_7_U750 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n755), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n752), .Y(alu_ashr_7_n710) );
  AO22X1_LVT alu_ashr_7_U749 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n713), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n710), .Y(alu_ashr_7_n650) );
  AO22X1_LVT alu_ashr_7_U748 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n816), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n817), .Y(alu_ashr_7_n753) );
  AO22X1_LVT alu_ashr_7_U747 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n814), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n815), .Y(alu_ashr_7_n750) );
  AO22X1_LVT alu_ashr_7_U746 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n753), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n750), .Y(alu_ashr_7_n711) );
  AO22X1_LVT alu_ashr_7_U745 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n812), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n813), .Y(alu_ashr_7_n751) );
  AO22X1_LVT alu_ashr_7_U744 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n810), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n811), .Y(alu_ashr_7_n548) );
  AO22X1_LVT alu_ashr_7_U743 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n751), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n548), .Y(alu_ashr_7_n627) );
  AO22X1_LVT alu_ashr_7_U742 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n711), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n627), .Y(alu_ashr_7_n809) );
  AO22X1_LVT alu_ashr_7_U741 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n650), 
        .A3(alu_ashr_7_n521), .A4(alu_ashr_7_n809), .Y(alu_ashr_7_n808) );
  AO22X1_LVT alu_ashr_7_U740 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n587), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n808), .Y(alu_n_T_101_10_) );
  AO22X1_LVT alu_ashr_7_U739 ( .A1(alu_ashr_7_n502), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n505), .A4(alu_shin_63_), .Y(alu_ashr_7_n789) );
  AO22X1_LVT alu_ashr_7_U738 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n789), .Y(alu_ashr_7_n747) );
  AO22X1_LVT alu_ashr_7_U737 ( .A1(alu_ashr_7_n502), .A2(alu_shin_62_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_61_), .Y(alu_ashr_7_n790) );
  AO22X1_LVT alu_ashr_7_U736 ( .A1(alu_ashr_7_n502), .A2(alu_shin_60_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_59_), .Y(alu_ashr_7_n787) );
  AO22X1_LVT alu_ashr_7_U735 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n790), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n787), .Y(alu_ashr_7_n745) );
  AO22X1_LVT alu_ashr_7_U734 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n747), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n745), .Y(alu_ashr_7_n707) );
  AO22X1_LVT alu_ashr_7_U733 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n707), .Y(alu_ashr_7_n647) );
  AO22X1_LVT alu_ashr_7_U732 ( .A1(alu_ashr_7_n502), .A2(alu_shin_58_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_57_), .Y(alu_ashr_7_n788) );
  AO22X1_LVT alu_ashr_7_U731 ( .A1(alu_ashr_7_n502), .A2(alu_shin_56_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_55_), .Y(alu_ashr_7_n785) );
  AO22X1_LVT alu_ashr_7_U730 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n788), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n785), .Y(alu_ashr_7_n746) );
  AO22X1_LVT alu_ashr_7_U729 ( .A1(alu_ashr_7_n502), .A2(alu_shin_54_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_53_), .Y(alu_ashr_7_n786) );
  AO22X1_LVT alu_ashr_7_U728 ( .A1(alu_ashr_7_n502), .A2(alu_shin_52_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_51_), .Y(alu_ashr_7_n783) );
  AO22X1_LVT alu_ashr_7_U727 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n786), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n783), .Y(alu_ashr_7_n743) );
  AO22X1_LVT alu_ashr_7_U726 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n746), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n743), .Y(alu_ashr_7_n708) );
  AO22X1_LVT alu_ashr_7_U725 ( .A1(alu_ashr_7_n502), .A2(alu_shin_50_), .A3(
        alu_ashr_7_n505), .A4(alu_shin_49_), .Y(alu_ashr_7_n784) );
  AO22X1_LVT alu_ashr_7_U724 ( .A1(alu_ashr_7_n502), .A2(alu_shin_48_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_47_), .Y(alu_ashr_7_n781) );
  AO22X1_LVT alu_ashr_7_U723 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n784), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n781), .Y(alu_ashr_7_n744) );
  AO22X1_LVT alu_ashr_7_U722 ( .A1(alu_ashr_7_n502), .A2(alu_shin_46_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_45_), .Y(alu_ashr_7_n782) );
  AO22X1_LVT alu_ashr_7_U721 ( .A1(alu_ashr_7_n502), .A2(alu_shin_44_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_43_), .Y(alu_ashr_7_n779) );
  AO22X1_LVT alu_ashr_7_U720 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n782), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n779), .Y(alu_ashr_7_n741) );
  AO22X1_LVT alu_ashr_7_U719 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n744), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n741), .Y(alu_ashr_7_n705) );
  AO22X1_LVT alu_ashr_7_U718 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n708), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n705), .Y(alu_ashr_7_n645) );
  AO22X1_LVT alu_ashr_7_U717 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n647), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n645), .Y(alu_ashr_7_n586) );
  AO22X1_LVT alu_ashr_7_U716 ( .A1(alu_ashr_7_n502), .A2(alu_shin_42_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_41_), .Y(alu_ashr_7_n780) );
  AO22X1_LVT alu_ashr_7_U715 ( .A1(alu_ashr_7_n502), .A2(alu_shin_40_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_39_), .Y(alu_ashr_7_n777) );
  AO22X1_LVT alu_ashr_7_U714 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n780), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n777), .Y(alu_ashr_7_n742) );
  AO22X1_LVT alu_ashr_7_U713 ( .A1(alu_ashr_7_n502), .A2(alu_shin_38_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_37_), .Y(alu_ashr_7_n778) );
  AO22X1_LVT alu_ashr_7_U712 ( .A1(alu_ashr_7_n502), .A2(alu_shin_36_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_35_), .Y(alu_ashr_7_n775) );
  AO22X1_LVT alu_ashr_7_U711 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n778), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n775), .Y(alu_ashr_7_n739) );
  AO22X1_LVT alu_ashr_7_U710 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n742), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n739), .Y(alu_ashr_7_n706) );
  AO22X1_LVT alu_ashr_7_U709 ( .A1(alu_ashr_7_n502), .A2(alu_shin_34_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_33_), .Y(alu_ashr_7_n776) );
  AO22X1_LVT alu_ashr_7_U708 ( .A1(alu_ashr_7_n502), .A2(alu_shin_32_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_31_), .Y(alu_ashr_7_n773) );
  AO22X1_LVT alu_ashr_7_U707 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n776), 
        .A3(alu_ashr_7_n493), .A4(alu_ashr_7_n773), .Y(alu_ashr_7_n740) );
  AO22X1_LVT alu_ashr_7_U706 ( .A1(alu_ashr_7_n502), .A2(alu_shin_30_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_29_), .Y(alu_ashr_7_n774) );
  AO22X1_LVT alu_ashr_7_U705 ( .A1(alu_ashr_7_n502), .A2(alu_shin_28_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_27_), .Y(alu_ashr_7_n771) );
  AO22X1_LVT alu_ashr_7_U704 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n774), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n771), .Y(alu_ashr_7_n737) );
  AO22X1_LVT alu_ashr_7_U703 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n740), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n737), .Y(alu_ashr_7_n703) );
  AO22X1_LVT alu_ashr_7_U702 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n706), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n703), .Y(alu_ashr_7_n646) );
  AO22X1_LVT alu_ashr_7_U701 ( .A1(alu_ashr_7_n502), .A2(alu_shin_26_), .A3(
        alu_ashr_7_n503), .A4(alu_shin_25_), .Y(alu_ashr_7_n772) );
  AO22X1_LVT alu_ashr_7_U700 ( .A1(alu_ashr_7_n502), .A2(alu_shin_24_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_23_), .Y(alu_ashr_7_n769) );
  AO22X1_LVT alu_ashr_7_U699 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n772), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n769), .Y(alu_ashr_7_n738) );
  AO22X1_LVT alu_ashr_7_U698 ( .A1(alu_ashr_7_n502), .A2(alu_shin_22_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_21_), .Y(alu_ashr_7_n770) );
  AO22X1_LVT alu_ashr_7_U697 ( .A1(alu_ashr_7_n502), .A2(alu_shin_20_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_19_), .Y(alu_ashr_7_n767) );
  AO22X1_LVT alu_ashr_7_U696 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n770), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n767), .Y(alu_ashr_7_n735) );
  AO22X1_LVT alu_ashr_7_U695 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n738), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n735), .Y(alu_ashr_7_n704) );
  AO22X1_LVT alu_ashr_7_U694 ( .A1(alu_ashr_7_n502), .A2(alu_shin_18_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_17_), .Y(alu_ashr_7_n768) );
  AO22X1_LVT alu_ashr_7_U693 ( .A1(alu_ashr_7_n502), .A2(alu_shin_16_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_15_), .Y(alu_ashr_7_n765) );
  AO22X1_LVT alu_ashr_7_U692 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n768), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n765), .Y(alu_ashr_7_n736) );
  AO22X1_LVT alu_ashr_7_U691 ( .A1(alu_ashr_7_n502), .A2(alu_shin_14_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_13_), .Y(alu_ashr_7_n766) );
  AO22X1_LVT alu_ashr_7_U690 ( .A1(alu_ashr_7_n502), .A2(alu_shin_12_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_11_), .Y(alu_ashr_7_n699) );
  AO22X1_LVT alu_ashr_7_U689 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n766), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n699), .Y(alu_ashr_7_n540) );
  AO22X1_LVT alu_ashr_7_U688 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n736), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n540), .Y(alu_ashr_7_n596) );
  AO22X1_LVT alu_ashr_7_U687 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n704), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n596), .Y(alu_ashr_7_n807) );
  AO22X1_LVT alu_ashr_7_U686 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n646), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n807), .Y(alu_ashr_7_n806) );
  AO22X1_LVT alu_ashr_7_U685 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n586), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n806), .Y(alu_n_T_101_11_) );
  AO22X1_LVT alu_ashr_7_U684 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n805), .Y(alu_ashr_7_n690) );
  AO22X1_LVT alu_ashr_7_U683 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n690), .Y(alu_ashr_7_n643) );
  AO22X1_LVT alu_ashr_7_U682 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n803), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n804), .Y(alu_ashr_7_n691) );
  AO22X1_LVT alu_ashr_7_U681 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n801), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n802), .Y(alu_ashr_7_n688) );
  AO22X1_LVT alu_ashr_7_U680 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n691), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n688), .Y(alu_ashr_7_n641) );
  AO22X1_LVT alu_ashr_7_U679 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n643), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n641), .Y(alu_ashr_7_n585) );
  AO22X1_LVT alu_ashr_7_U678 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n799), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n800), .Y(alu_ashr_7_n689) );
  AO22X1_LVT alu_ashr_7_U677 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n797), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n798), .Y(alu_ashr_7_n686) );
  AO22X1_LVT alu_ashr_7_U676 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n689), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n686), .Y(alu_ashr_7_n642) );
  AO22X1_LVT alu_ashr_7_U675 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n795), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n796), .Y(alu_ashr_7_n687) );
  AO22X1_LVT alu_ashr_7_U674 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n793), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n794), .Y(alu_ashr_7_n576) );
  AO22X1_LVT alu_ashr_7_U673 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n687), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n576), .Y(alu_ashr_7_n792) );
  AO22X1_LVT alu_ashr_7_U672 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n642), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n792), .Y(alu_ashr_7_n791) );
  AO22X1_LVT alu_ashr_7_U671 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n585), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n791), .Y(alu_n_T_101_12_) );
  AO22X1_LVT alu_ashr_7_U670 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n789), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n790), .Y(alu_ashr_7_n727) );
  AO22X1_LVT alu_ashr_7_U669 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n727), .Y(alu_ashr_7_n683) );
  AO22X1_LVT alu_ashr_7_U668 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n683), .Y(alu_ashr_7_n639) );
  AO22X1_LVT alu_ashr_7_U667 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n787), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n788), .Y(alu_ashr_7_n728) );
  AO22X1_LVT alu_ashr_7_U666 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n785), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n786), .Y(alu_ashr_7_n725) );
  AO22X1_LVT alu_ashr_7_U665 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n728), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n725), .Y(alu_ashr_7_n684) );
  AO22X1_LVT alu_ashr_7_U664 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n783), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n784), .Y(alu_ashr_7_n726) );
  AO22X1_LVT alu_ashr_7_U663 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n781), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n782), .Y(alu_ashr_7_n723) );
  AO22X1_LVT alu_ashr_7_U662 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n726), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n723), .Y(alu_ashr_7_n681) );
  AO22X1_LVT alu_ashr_7_U661 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n684), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n681), .Y(alu_ashr_7_n637) );
  AO22X1_LVT alu_ashr_7_U660 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n639), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n637), .Y(alu_ashr_7_n584) );
  AO22X1_LVT alu_ashr_7_U659 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n779), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n780), .Y(alu_ashr_7_n724) );
  AO22X1_LVT alu_ashr_7_U658 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n777), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n778), .Y(alu_ashr_7_n721) );
  AO22X1_LVT alu_ashr_7_U657 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n724), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n721), .Y(alu_ashr_7_n682) );
  AO22X1_LVT alu_ashr_7_U656 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n775), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n776), .Y(alu_ashr_7_n722) );
  AO22X1_LVT alu_ashr_7_U655 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n773), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n774), .Y(alu_ashr_7_n719) );
  AO22X1_LVT alu_ashr_7_U654 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n722), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n719), .Y(alu_ashr_7_n679) );
  AO22X1_LVT alu_ashr_7_U653 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n682), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n679), .Y(alu_ashr_7_n638) );
  AO22X1_LVT alu_ashr_7_U652 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n771), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n772), .Y(alu_ashr_7_n720) );
  AO22X1_LVT alu_ashr_7_U651 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n769), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n770), .Y(alu_ashr_7_n717) );
  AO22X1_LVT alu_ashr_7_U650 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n720), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n717), .Y(alu_ashr_7_n680) );
  AO22X1_LVT alu_ashr_7_U649 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n767), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n768), .Y(alu_ashr_7_n718) );
  AO22X1_LVT alu_ashr_7_U648 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n765), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n766), .Y(alu_ashr_7_n698) );
  AO22X1_LVT alu_ashr_7_U647 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n718), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n698), .Y(alu_ashr_7_n558) );
  AO22X1_LVT alu_ashr_7_U646 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n680), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n558), .Y(alu_ashr_7_n764) );
  AO22X1_LVT alu_ashr_7_U645 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n638), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n764), .Y(alu_ashr_7_n763) );
  AO22X1_LVT alu_ashr_7_U644 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n584), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n763), .Y(alu_n_T_101_13_) );
  AO22X1_LVT alu_ashr_7_U643 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n762), .Y(alu_ashr_7_n676) );
  AO22X1_LVT alu_ashr_7_U642 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n676), .Y(alu_ashr_7_n623) );
  AO22X1_LVT alu_ashr_7_U641 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n760), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n761), .Y(alu_ashr_7_n677) );
  AO22X1_LVT alu_ashr_7_U640 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n758), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n759), .Y(alu_ashr_7_n674) );
  AO22X1_LVT alu_ashr_7_U639 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n677), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n674), .Y(alu_ashr_7_n621) );
  AO22X1_LVT alu_ashr_7_U638 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n623), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n621), .Y(alu_ashr_7_n583) );
  AO22X1_LVT alu_ashr_7_U637 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n756), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n757), .Y(alu_ashr_7_n675) );
  AO22X1_LVT alu_ashr_7_U636 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n754), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n755), .Y(alu_ashr_7_n672) );
  AO22X1_LVT alu_ashr_7_U635 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n675), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n672), .Y(alu_ashr_7_n622) );
  AO22X1_LVT alu_ashr_7_U634 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n752), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n753), .Y(alu_ashr_7_n673) );
  AO22X1_LVT alu_ashr_7_U633 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n750), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n751), .Y(alu_ashr_7_n546) );
  AO22X1_LVT alu_ashr_7_U632 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n673), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n546), .Y(alu_ashr_7_n749) );
  AO22X1_LVT alu_ashr_7_U631 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n622), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n749), .Y(alu_ashr_7_n748) );
  AO22X1_LVT alu_ashr_7_U630 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n583), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n748), .Y(alu_n_T_101_14_) );
  AO22X1_LVT alu_ashr_7_U629 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n496), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n747), .Y(alu_ashr_7_n669) );
  AO22X1_LVT alu_ashr_7_U628 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n669), .Y(alu_ashr_7_n619) );
  AO22X1_LVT alu_ashr_7_U627 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n745), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n746), .Y(alu_ashr_7_n670) );
  AO22X1_LVT alu_ashr_7_U626 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n743), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n744), .Y(alu_ashr_7_n667) );
  AO22X1_LVT alu_ashr_7_U625 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n670), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n667), .Y(alu_ashr_7_n617) );
  AO22X1_LVT alu_ashr_7_U624 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n619), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n617), .Y(alu_ashr_7_n582) );
  AO22X1_LVT alu_ashr_7_U623 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n741), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n742), .Y(alu_ashr_7_n668) );
  AO22X1_LVT alu_ashr_7_U622 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n739), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n740), .Y(alu_ashr_7_n665) );
  AO22X1_LVT alu_ashr_7_U621 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n668), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n665), .Y(alu_ashr_7_n618) );
  AO22X1_LVT alu_ashr_7_U620 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n737), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n738), .Y(alu_ashr_7_n666) );
  AO22X1_LVT alu_ashr_7_U619 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n735), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n736), .Y(alu_ashr_7_n538) );
  AO22X1_LVT alu_ashr_7_U618 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n666), 
        .A3(alu_ashr_7_n515), .A4(alu_ashr_7_n538), .Y(alu_ashr_7_n734) );
  AO22X1_LVT alu_ashr_7_U617 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n618), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n734), .Y(alu_ashr_7_n733) );
  AO22X1_LVT alu_ashr_7_U616 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n582), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n733), .Y(alu_n_T_101_15_) );
  AO22X1_LVT alu_ashr_7_U615 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n732), .Y(alu_ashr_7_n581) );
  AO22X1_LVT alu_ashr_7_U614 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n730), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n731), .Y(alu_ashr_7_n729) );
  AO22X1_LVT alu_ashr_7_U613 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n581), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n729), .Y(alu_n_T_101_16_) );
  AO22X1_LVT alu_ashr_7_U612 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n727), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n728), .Y(alu_ashr_7_n657) );
  AO22X1_LVT alu_ashr_7_U611 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n725), 
        .A3(alu_ashr_7_n510), .A4(alu_ashr_7_n726), .Y(alu_ashr_7_n655) );
  AO22X1_LVT alu_ashr_7_U610 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n657), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n655), .Y(alu_ashr_7_n700) );
  AO22X1_LVT alu_ashr_7_U609 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n700), .Y(alu_ashr_7_n580) );
  AO22X1_LVT alu_ashr_7_U608 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n723), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n724), .Y(alu_ashr_7_n656) );
  AO22X1_LVT alu_ashr_7_U607 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n721), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n722), .Y(alu_ashr_7_n653) );
  AO22X1_LVT alu_ashr_7_U606 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n656), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n653), .Y(alu_ashr_7_n701) );
  AO22X1_LVT alu_ashr_7_U605 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n719), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n720), .Y(alu_ashr_7_n654) );
  AO22X1_LVT alu_ashr_7_U604 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n717), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n718), .Y(alu_ashr_7_n526) );
  AO22X1_LVT alu_ashr_7_U603 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n654), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n526), .Y(alu_ashr_7_n693) );
  AO22X1_LVT alu_ashr_7_U602 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n701), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n693), .Y(alu_ashr_7_n716) );
  AO22X1_LVT alu_ashr_7_U601 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n580), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n716), .Y(alu_n_T_101_17_) );
  AO22X1_LVT alu_ashr_7_U600 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n714), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n715), .Y(alu_ashr_7_n634) );
  AO22X1_LVT alu_ashr_7_U599 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n634), .Y(alu_ashr_7_n571) );
  AO22X1_LVT alu_ashr_7_U598 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n712), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n713), .Y(alu_ashr_7_n635) );
  AO22X1_LVT alu_ashr_7_U597 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n710), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n711), .Y(alu_ashr_7_n625) );
  AO22X1_LVT alu_ashr_7_U596 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n635), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n625), .Y(alu_ashr_7_n709) );
  AO22X1_LVT alu_ashr_7_U595 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n571), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n709), .Y(alu_n_T_101_18_) );
  AO22X1_LVT alu_ashr_7_U594 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n707), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n708), .Y(alu_ashr_7_n611) );
  AO22X1_LVT alu_ashr_7_U593 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n611), .Y(alu_ashr_7_n570) );
  AO22X1_LVT alu_ashr_7_U592 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n705), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n706), .Y(alu_ashr_7_n612) );
  AO22X1_LVT alu_ashr_7_U591 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n703), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n704), .Y(alu_ashr_7_n594) );
  AO22X1_LVT alu_ashr_7_U590 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n612), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n594), .Y(alu_ashr_7_n702) );
  AO22X1_LVT alu_ashr_7_U589 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n570), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n702), .Y(alu_n_T_101_19_) );
  AO22X1_LVT alu_ashr_7_U588 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n700), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n701), .Y(alu_ashr_7_n614) );
  AO22X1_LVT alu_ashr_7_U587 ( .A1(alu_ashr_7_n502), .A2(alu_shin_10_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_9_), .Y(alu_ashr_7_n601) );
  AO22X1_LVT alu_ashr_7_U586 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n699), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n601), .Y(alu_ashr_7_n560) );
  AO22X1_LVT alu_ashr_7_U585 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n698), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n560), .Y(alu_ashr_7_n527) );
  AO22X1_LVT alu_ashr_7_U584 ( .A1(alu_ashr_7_n502), .A2(alu_shin_8_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_7_), .Y(alu_ashr_7_n602) );
  AO22X1_LVT alu_ashr_7_U583 ( .A1(alu_ashr_7_n502), .A2(alu_shin_6_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_5_), .Y(alu_ashr_7_n599) );
  AO22X1_LVT alu_ashr_7_U582 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n602), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n599), .Y(alu_ashr_7_n561) );
  AO22X1_LVT alu_ashr_7_U581 ( .A1(alu_ashr_7_n502), .A2(alu_shin_4_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_3_), .Y(alu_ashr_7_n600) );
  AO22X1_LVT alu_ashr_7_U580 ( .A1(alu_ashr_7_n502), .A2(alu_shin_2_), .A3(
        alu_ashr_7_n504), .A4(alu_shin_1_), .Y(alu_ashr_7_n697) );
  AO22X1_LVT alu_ashr_7_U579 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n600), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n697), .Y(alu_ashr_7_n696) );
  AO22X1_LVT alu_ashr_7_U578 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n561), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n696), .Y(alu_ashr_7_n695) );
  AO22X1_LVT alu_ashr_7_U577 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n527), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n695), .Y(alu_ashr_7_n694) );
  AO22X1_LVT alu_ashr_7_U576 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n693), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n694), .Y(alu_ashr_7_n692) );
  AO22X1_LVT alu_ashr_7_U575 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n614), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n692), .Y(alu_n_T_101_1_) );
  AO22X1_LVT alu_ashr_7_U574 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n690), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n691), .Y(alu_ashr_7_n609) );
  AO22X1_LVT alu_ashr_7_U573 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n609), .Y(alu_ashr_7_n569) );
  AO22X1_LVT alu_ashr_7_U572 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n688), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n689), .Y(alu_ashr_7_n610) );
  AO22X1_LVT alu_ashr_7_U571 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n686), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n687), .Y(alu_ashr_7_n574) );
  AO22X1_LVT alu_ashr_7_U570 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n610), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n574), .Y(alu_ashr_7_n685) );
  AO22X1_LVT alu_ashr_7_U569 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n569), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n685), .Y(alu_n_T_101_20_) );
  AO22X1_LVT alu_ashr_7_U568 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n683), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n684), .Y(alu_ashr_7_n607) );
  AO22X1_LVT alu_ashr_7_U567 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n607), .Y(alu_ashr_7_n568) );
  AO22X1_LVT alu_ashr_7_U566 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n681), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n682), .Y(alu_ashr_7_n608) );
  AO22X1_LVT alu_ashr_7_U565 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n679), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n680), .Y(alu_ashr_7_n556) );
  AO22X1_LVT alu_ashr_7_U564 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n608), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n556), .Y(alu_ashr_7_n678) );
  AO22X1_LVT alu_ashr_7_U563 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n568), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n678), .Y(alu_n_T_101_21_) );
  AO22X1_LVT alu_ashr_7_U562 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n676), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n677), .Y(alu_ashr_7_n605) );
  AO22X1_LVT alu_ashr_7_U561 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n605), .Y(alu_ashr_7_n567) );
  AO22X1_LVT alu_ashr_7_U560 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n674), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n675), .Y(alu_ashr_7_n606) );
  AO22X1_LVT alu_ashr_7_U559 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n672), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n673), .Y(alu_ashr_7_n544) );
  AO22X1_LVT alu_ashr_7_U558 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n606), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n544), .Y(alu_ashr_7_n671) );
  AO22X1_LVT alu_ashr_7_U557 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n567), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n671), .Y(alu_n_T_101_22_) );
  AO22X1_LVT alu_ashr_7_U556 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n669), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n670), .Y(alu_ashr_7_n603) );
  AO22X1_LVT alu_ashr_7_U555 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n603), .Y(alu_ashr_7_n566) );
  AO22X1_LVT alu_ashr_7_U554 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n667), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n668), .Y(alu_ashr_7_n604) );
  AO22X1_LVT alu_ashr_7_U553 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n665), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n666), .Y(alu_ashr_7_n536) );
  AO22X1_LVT alu_ashr_7_U552 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n604), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n536), .Y(alu_ashr_7_n664) );
  AO22X1_LVT alu_ashr_7_U551 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n566), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n664), .Y(alu_n_T_101_23_) );
  AO22X1_LVT alu_ashr_7_U550 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n663), .Y(alu_ashr_7_n590) );
  AO22X1_LVT alu_ashr_7_U549 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n590), .Y(alu_ashr_7_n565) );
  AO22X1_LVT alu_ashr_7_U548 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n661), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n662), .Y(alu_ashr_7_n591) );
  AO22X1_LVT alu_ashr_7_U547 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n659), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n660), .Y(alu_ashr_7_n530) );
  AO22X1_LVT alu_ashr_7_U546 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n591), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n530), .Y(alu_ashr_7_n658) );
  AO22X1_LVT alu_ashr_7_U545 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n565), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n658), .Y(alu_n_T_101_24_) );
  AO22X1_LVT alu_ashr_7_U544 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n657), .Y(alu_ashr_7_n588) );
  AO22X1_LVT alu_ashr_7_U543 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n588), .Y(alu_ashr_7_n564) );
  AO22X1_LVT alu_ashr_7_U542 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n655), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n656), .Y(alu_ashr_7_n589) );
  AO22X1_LVT alu_ashr_7_U541 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n653), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n654), .Y(alu_ashr_7_n524) );
  AO22X1_LVT alu_ashr_7_U540 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n589), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n524), .Y(alu_ashr_7_n652) );
  AO22X1_LVT alu_ashr_7_U539 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n564), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n652), .Y(alu_n_T_101_25_) );
  AO22X1_LVT alu_ashr_7_U538 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n651), .Y(alu_ashr_7_n563) );
  AO22X1_LVT alu_ashr_7_U537 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n649), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n650), .Y(alu_ashr_7_n648) );
  AO22X1_LVT alu_ashr_7_U536 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n563), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n648), .Y(alu_n_T_101_26_) );
  AO22X1_LVT alu_ashr_7_U535 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n647), .Y(alu_ashr_7_n562) );
  AO22X1_LVT alu_ashr_7_U534 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n645), 
        .A3(alu_ashr_7_n520), .A4(alu_ashr_7_n646), .Y(alu_ashr_7_n644) );
  AO22X1_LVT alu_ashr_7_U533 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n562), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n644), .Y(alu_n_T_101_27_) );
  AO22X1_LVT alu_ashr_7_U532 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n643), .Y(alu_ashr_7_n553) );
  AO22X1_LVT alu_ashr_7_U531 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n641), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n642), .Y(alu_ashr_7_n640) );
  AO22X1_LVT alu_ashr_7_U530 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n553), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n640), .Y(alu_n_T_101_28_) );
  AO22X1_LVT alu_ashr_7_U529 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n639), .Y(alu_ashr_7_n552) );
  AO22X1_LVT alu_ashr_7_U528 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n637), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n638), .Y(alu_ashr_7_n636) );
  AO22X1_LVT alu_ashr_7_U527 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n552), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n636), .Y(alu_n_T_101_29_) );
  AO22X1_LVT alu_ashr_7_U526 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n634), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n635), .Y(alu_ashr_7_n613) );
  AO22X1_LVT alu_ashr_7_U525 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n632), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n633), .Y(alu_ashr_7_n549) );
  AO22X1_LVT alu_ashr_7_U524 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n630), 
        .A3(alu_ashr_7_n508), .A4(alu_ashr_7_n631), .Y(alu_ashr_7_n629) );
  AO22X1_LVT alu_ashr_7_U523 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n549), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n629), .Y(alu_ashr_7_n628) );
  AO22X1_LVT alu_ashr_7_U522 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n627), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n628), .Y(alu_ashr_7_n626) );
  AO22X1_LVT alu_ashr_7_U521 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n625), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n626), .Y(alu_ashr_7_n624) );
  AO22X1_LVT alu_ashr_7_U520 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n613), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n624), .Y(alu_n_T_101_2_) );
  AO22X1_LVT alu_ashr_7_U519 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n623), .Y(alu_ashr_7_n551) );
  AO22X1_LVT alu_ashr_7_U518 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n621), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n622), .Y(alu_ashr_7_n620) );
  AO22X1_LVT alu_ashr_7_U517 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n551), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n620), .Y(alu_n_T_101_30_) );
  AO22X1_LVT alu_ashr_7_U516 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n619), .Y(alu_ashr_7_n550) );
  AO22X1_LVT alu_ashr_7_U515 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n617), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n618), .Y(alu_ashr_7_n616) );
  AO22X1_LVT alu_ashr_7_U514 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n550), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n616), .Y(alu_n_T_101_31_) );
  AO22X1_LVT alu_ashr_7_U513 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n501), .A4(alu_ashr_7_n615), .Y(alu_n_T_101_32_) );
  AO22X1_LVT alu_ashr_7_U512 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n614), .Y(alu_n_T_101_33_) );
  AO22X1_LVT alu_ashr_7_U511 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n613), .Y(alu_n_T_101_34_) );
  AO22X1_LVT alu_ashr_7_U510 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n611), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n612), .Y(alu_ashr_7_n592) );
  AO22X1_LVT alu_ashr_7_U509 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n592), .Y(alu_n_T_101_35_) );
  AO22X1_LVT alu_ashr_7_U508 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n609), 
        .A3(alu_ashr_7_n519), .A4(alu_ashr_7_n610), .Y(alu_ashr_7_n572) );
  AO22X1_LVT alu_ashr_7_U507 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n497), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n572), .Y(alu_n_T_101_36_) );
  AO22X1_LVT alu_ashr_7_U506 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n607), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n608), .Y(alu_ashr_7_n554) );
  AO22X1_LVT alu_ashr_7_U505 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n554), .Y(alu_n_T_101_37_) );
  AO22X1_LVT alu_ashr_7_U504 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n605), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n606), .Y(alu_ashr_7_n542) );
  AO22X1_LVT alu_ashr_7_U503 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n542), .Y(alu_n_T_101_38_) );
  AO22X1_LVT alu_ashr_7_U502 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n603), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n604), .Y(alu_ashr_7_n534) );
  AO22X1_LVT alu_ashr_7_U501 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n534), .Y(alu_n_T_101_39_) );
  AO22X1_LVT alu_ashr_7_U500 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n601), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n602), .Y(alu_ashr_7_n541) );
  AO22X1_LVT alu_ashr_7_U499 ( .A1(alu_ashr_7_n506), .A2(alu_ashr_7_n599), 
        .A3(alu_ashr_7_n507), .A4(alu_ashr_7_n600), .Y(alu_ashr_7_n598) );
  AO22X1_LVT alu_ashr_7_U498 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n541), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n598), .Y(alu_ashr_7_n597) );
  AO22X1_LVT alu_ashr_7_U497 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n596), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n597), .Y(alu_ashr_7_n595) );
  AO22X1_LVT alu_ashr_7_U496 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n594), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n595), .Y(alu_ashr_7_n593) );
  AO22X1_LVT alu_ashr_7_U495 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n592), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n593), .Y(alu_n_T_101_3_) );
  AO22X1_LVT alu_ashr_7_U494 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n590), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n591), .Y(alu_ashr_7_n528) );
  AO22X1_LVT alu_ashr_7_U493 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n528), .Y(alu_n_T_101_40_) );
  AO22X1_LVT alu_ashr_7_U492 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n588), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n589), .Y(alu_ashr_7_n522) );
  AO22X1_LVT alu_ashr_7_U491 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n522), .Y(alu_n_T_101_41_) );
  AO22X1_LVT alu_ashr_7_U490 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n587), .Y(alu_n_T_101_42_) );
  AO22X1_LVT alu_ashr_7_U489 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n586), .Y(alu_n_T_101_43_) );
  AO22X1_LVT alu_ashr_7_U488 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n585), .Y(alu_n_T_101_44_) );
  AO22X1_LVT alu_ashr_7_U487 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n500), .A4(alu_ashr_7_n584), .Y(alu_n_T_101_45_) );
  AO22X1_LVT alu_ashr_7_U486 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n583), .Y(alu_n_T_101_46_) );
  AO22X1_LVT alu_ashr_7_U485 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n582), .Y(alu_n_T_101_47_) );
  AO22X1_LVT alu_ashr_7_U484 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n581), .Y(alu_n_T_101_48_) );
  AO22X1_LVT alu_ashr_7_U483 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n580), .Y(alu_n_T_101_49_) );
  AO22X1_LVT alu_ashr_7_U482 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n578), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n579), .Y(alu_ashr_7_n577) );
  AO22X1_LVT alu_ashr_7_U481 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n576), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n577), .Y(alu_ashr_7_n575) );
  AO22X1_LVT alu_ashr_7_U480 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n574), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n575), .Y(alu_ashr_7_n573) );
  AO22X1_LVT alu_ashr_7_U479 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n572), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n573), .Y(alu_n_T_101_4_) );
  AO22X1_LVT alu_ashr_7_U478 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n571), .Y(alu_n_T_101_50_) );
  AO22X1_LVT alu_ashr_7_U477 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n570), .Y(alu_n_T_101_51_) );
  AO22X1_LVT alu_ashr_7_U476 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n569), .Y(alu_n_T_101_52_) );
  AO22X1_LVT alu_ashr_7_U475 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n568), .Y(alu_n_T_101_53_) );
  AO22X1_LVT alu_ashr_7_U474 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n567), .Y(alu_n_T_101_54_) );
  AO22X1_LVT alu_ashr_7_U473 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n566), .Y(alu_n_T_101_55_) );
  AO22X1_LVT alu_ashr_7_U472 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n565), .Y(alu_n_T_101_56_) );
  AO22X1_LVT alu_ashr_7_U471 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n564), .Y(alu_n_T_101_57_) );
  AO22X1_LVT alu_ashr_7_U470 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n563), .Y(alu_n_T_101_58_) );
  AO22X1_LVT alu_ashr_7_U469 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n562), .Y(alu_n_T_101_59_) );
  AO22X1_LVT alu_ashr_7_U468 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n560), 
        .A3(alu_ashr_7_n511), .A4(alu_ashr_7_n561), .Y(alu_ashr_7_n559) );
  AO22X1_LVT alu_ashr_7_U467 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n558), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n559), .Y(alu_ashr_7_n557) );
  AO22X1_LVT alu_ashr_7_U466 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n556), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n557), .Y(alu_ashr_7_n555) );
  AO22X1_LVT alu_ashr_7_U465 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n554), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n555), .Y(alu_n_T_101_5_) );
  AO22X1_LVT alu_ashr_7_U464 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n498), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n553), .Y(alu_n_T_101_60_) );
  AO22X1_LVT alu_ashr_7_U463 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n552), .Y(alu_n_T_101_61_) );
  AO22X1_LVT alu_ashr_7_U462 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n551), .Y(alu_n_T_101_62_) );
  AO22X1_LVT alu_ashr_7_U461 ( .A1(alu_ashr_7_n499), .A2(alu_n_T_100_64_), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n550), .Y(alu_n_T_101_63_) );
  AO22X1_LVT alu_ashr_7_U460 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n548), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n549), .Y(alu_ashr_7_n547) );
  AO22X1_LVT alu_ashr_7_U459 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n546), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n547), .Y(alu_ashr_7_n545) );
  AO22X1_LVT alu_ashr_7_U458 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n544), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n545), .Y(alu_ashr_7_n543) );
  AO22X1_LVT alu_ashr_7_U457 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n542), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n543), .Y(alu_n_T_101_6_) );
  AO22X1_LVT alu_ashr_7_U456 ( .A1(alu_ashr_7_n509), .A2(alu_ashr_7_n540), 
        .A3(alu_ashr_7_n492), .A4(alu_ashr_7_n541), .Y(alu_ashr_7_n539) );
  AO22X1_LVT alu_ashr_7_U455 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n538), 
        .A3(alu_ashr_7_n516), .A4(alu_ashr_7_n539), .Y(alu_ashr_7_n537) );
  AO22X1_LVT alu_ashr_7_U454 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n536), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n537), .Y(alu_ashr_7_n535) );
  AO22X1_LVT alu_ashr_7_U453 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n534), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n535), .Y(alu_n_T_101_7_) );
  AO22X1_LVT alu_ashr_7_U452 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n532), 
        .A3(alu_ashr_7_n514), .A4(alu_ashr_7_n533), .Y(alu_ashr_7_n531) );
  AO22X1_LVT alu_ashr_7_U451 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n530), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n531), .Y(alu_ashr_7_n529) );
  AO22X1_LVT alu_ashr_7_U450 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n528), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n529), .Y(alu_n_T_101_8_) );
  AO22X1_LVT alu_ashr_7_U449 ( .A1(alu_ashr_7_n512), .A2(alu_ashr_7_n526), 
        .A3(alu_ashr_7_n513), .A4(alu_ashr_7_n527), .Y(alu_ashr_7_n525) );
  AO22X1_LVT alu_ashr_7_U448 ( .A1(alu_ashr_7_n517), .A2(alu_ashr_7_n524), 
        .A3(alu_ashr_7_n518), .A4(alu_ashr_7_n525), .Y(alu_ashr_7_n523) );
  AO22X1_LVT alu_ashr_7_U447 ( .A1(alu_ashr_7_n499), .A2(alu_ashr_7_n522), 
        .A3(alu_ashr_7_n495), .A4(alu_ashr_7_n523), .Y(alu_n_T_101_9_) );
  NBUFFX2_LVT alu_ashr_7_U446 ( .A(alu_n_T_100_64_), .Y(alu_ashr_7_n498) );
  NBUFFX2_LVT alu_ashr_7_U445 ( .A(alu_n_T_100_64_), .Y(alu_ashr_7_n497) );
  NBUFFX2_LVT alu_ashr_7_U444 ( .A(alu_n_T_100_64_), .Y(alu_ashr_7_n496) );
  INVX1_LVT alu_ashr_7_U443 ( .A(alu_ashr_7_n517), .Y(alu_ashr_7_n521) );
  NBUFFX2_LVT alu_ashr_7_U442 ( .A(alu_io_in2[0]), .Y(alu_ashr_7_n502) );
  NBUFFX2_LVT alu_ashr_7_U441 ( .A(alu_io_in2[1]), .Y(alu_ashr_7_n506) );
  NBUFFX2_LVT alu_ashr_7_U440 ( .A(alu_io_in2[2]), .Y(alu_ashr_7_n509) );
  INVX1_LVT alu_ashr_7_U439 ( .A(alu_ashr_7_n512), .Y(alu_ashr_7_n516) );
  INVX1_LVT alu_ashr_7_U438 ( .A(alu_ashr_7_n517), .Y(alu_ashr_7_n519) );
  NBUFFX2_LVT alu_ashr_7_U437 ( .A(alu_io_in2[3]), .Y(alu_ashr_7_n512) );
  NBUFFX2_LVT alu_ashr_7_U436 ( .A(alu_io_in2[4]), .Y(alu_ashr_7_n517) );
  NBUFFX4_LVT alu_ashr_7_U435 ( .A(alu_shamt_5_), .Y(alu_ashr_7_n499) );
  IBUFFX2_LVT alu_ashr_7_U434 ( .A(alu_ashr_7_n517), .Y(alu_ashr_7_n518) );
  IBUFFX2_LVT alu_ashr_7_U433 ( .A(alu_ashr_7_n517), .Y(alu_ashr_7_n520) );
  IBUFFX4_LVT alu_ashr_7_U432 ( .A(alu_ashr_7_n509), .Y(alu_ashr_7_n492) );
  IBUFFX2_LVT alu_ashr_7_U431 ( .A(alu_ashr_7_n509), .Y(alu_ashr_7_n511) );
  IBUFFX2_LVT alu_ashr_7_U430 ( .A(alu_ashr_7_n509), .Y(alu_ashr_7_n510) );
  IBUFFX4_LVT alu_ashr_7_U429 ( .A(alu_ashr_7_n499), .Y(alu_ashr_7_n495) );
  IBUFFX2_LVT alu_ashr_7_U428 ( .A(alu_ashr_7_n499), .Y(alu_ashr_7_n501) );
  IBUFFX2_LVT alu_ashr_7_U427 ( .A(alu_ashr_7_n499), .Y(alu_ashr_7_n500) );
  IBUFFX2_LVT alu_ashr_7_U426 ( .A(alu_ashr_7_n512), .Y(alu_ashr_7_n513) );
  IBUFFX2_LVT alu_ashr_7_U425 ( .A(alu_ashr_7_n512), .Y(alu_ashr_7_n515) );
  IBUFFX2_LVT alu_ashr_7_U424 ( .A(alu_ashr_7_n512), .Y(alu_ashr_7_n514) );
  IBUFFX2_LVT alu_ashr_7_U423 ( .A(alu_ashr_7_n502), .Y(alu_ashr_7_n503) );
  IBUFFX2_LVT alu_ashr_7_U422 ( .A(alu_ashr_7_n502), .Y(alu_ashr_7_n505) );
  IBUFFX2_LVT alu_ashr_7_U421 ( .A(alu_ashr_7_n506), .Y(alu_ashr_7_n507) );
  IBUFFX2_LVT alu_ashr_7_U420 ( .A(alu_ashr_7_n506), .Y(alu_ashr_7_n508) );
  IBUFFX2_LVT alu_ashr_7_U419 ( .A(alu_ashr_7_n506), .Y(alu_ashr_7_n493) );
  IBUFFX2_LVT alu_ashr_7_U418 ( .A(alu_ashr_7_n502), .Y(alu_ashr_7_n504) );
  NAND4X0_LVT div_U1248 ( .A1(div_n755), .A2(div_n993), .A3(div_n992), .A4(
        div_n991), .Y(div_n994) );
  NAND4X0_LVT div_U1247 ( .A1(div_n756), .A2(div_n989), .A3(div_n988), .A4(
        div_n987), .Y(div_n995) );
  NAND4X0_LVT div_U1246 ( .A1(div_n757), .A2(div_n986), .A3(div_n985), .A4(
        div_n984), .Y(div_n996) );
  AO22X1_LVT div_U1245 ( .A1(div_n146), .A2(div_result_41_), .A3(div_n209), 
        .A4(div_result_9_), .Y(div_io_resp_bits_data[9]) );
  AO22X1_LVT div_U1244 ( .A1(div_n146), .A2(div_result_40_), .A3(div_n209), 
        .A4(div_result_8_), .Y(div_io_resp_bits_data[8]) );
  AO22X1_LVT div_U1243 ( .A1(div_n146), .A2(div_result_39_), .A3(div_n209), 
        .A4(div_result_7_), .Y(div_io_resp_bits_data[7]) );
  AO22X1_LVT div_U1242 ( .A1(div_n146), .A2(div_result_38_), .A3(div_n209), 
        .A4(div_result_6_), .Y(div_io_resp_bits_data[6]) );
  AO22X1_LVT div_U1241 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_63_), .Y(div_io_resp_bits_data[63]) );
  AO22X1_LVT div_U1240 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_62_), .Y(div_io_resp_bits_data[62]) );
  AO22X1_LVT div_U1239 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_61_), .Y(div_io_resp_bits_data[61]) );
  AO22X1_LVT div_U1238 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_60_), .Y(div_io_resp_bits_data[60]) );
  AO22X1_LVT div_U1237 ( .A1(div_n146), .A2(div_result_37_), .A3(div_n209), 
        .A4(div_result_5_), .Y(div_io_resp_bits_data[5]) );
  AO22X1_LVT div_U1236 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_59_), .Y(div_io_resp_bits_data[59]) );
  AO22X1_LVT div_U1235 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_58_), .Y(div_io_resp_bits_data[58]) );
  AO22X1_LVT div_U1234 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_57_), .Y(div_io_resp_bits_data[57]) );
  AO22X1_LVT div_U1233 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_56_), .Y(div_io_resp_bits_data[56]) );
  AO22X1_LVT div_U1232 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_55_), .Y(div_io_resp_bits_data[55]) );
  AO22X1_LVT div_U1231 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_54_), .Y(div_io_resp_bits_data[54]) );
  AO22X1_LVT div_U1230 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_53_), .Y(div_io_resp_bits_data[53]) );
  AO22X1_LVT div_U1229 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_52_), .Y(div_io_resp_bits_data[52]) );
  AO22X1_LVT div_U1228 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_51_), .Y(div_io_resp_bits_data[51]) );
  AO22X1_LVT div_U1227 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_50_), .Y(div_io_resp_bits_data[50]) );
  AO22X1_LVT div_U1226 ( .A1(div_n146), .A2(div_result_36_), .A3(div_n209), 
        .A4(div_result_4_), .Y(div_io_resp_bits_data[4]) );
  AO22X1_LVT div_U1225 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_49_), .Y(div_io_resp_bits_data[49]) );
  AO22X1_LVT div_U1224 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_48_), .Y(div_io_resp_bits_data[48]) );
  AO22X1_LVT div_U1223 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_47_), .Y(div_io_resp_bits_data[47]) );
  AO22X1_LVT div_U1222 ( .A1(div_n244), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_46_), .Y(div_io_resp_bits_data[46]) );
  AO22X1_LVT div_U1221 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_45_), .Y(div_io_resp_bits_data[45]) );
  AO22X1_LVT div_U1220 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_44_), .Y(div_io_resp_bits_data[44]) );
  AO22X1_LVT div_U1219 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_43_), .Y(div_io_resp_bits_data[43]) );
  AO22X1_LVT div_U1218 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_42_), .Y(div_io_resp_bits_data[42]) );
  AO22X1_LVT div_U1217 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_41_), .Y(div_io_resp_bits_data[41]) );
  AO22X1_LVT div_U1216 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_40_), .Y(div_io_resp_bits_data[40]) );
  AO22X1_LVT div_U1215 ( .A1(div_n146), .A2(div_result_35_), .A3(div_n209), 
        .A4(div_result_3_), .Y(div_io_resp_bits_data[3]) );
  AO22X1_LVT div_U1214 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_39_), .Y(div_io_resp_bits_data[39]) );
  AO22X1_LVT div_U1213 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_38_), .Y(div_io_resp_bits_data[38]) );
  AO22X1_LVT div_U1212 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_37_), .Y(div_io_resp_bits_data[37]) );
  AO22X1_LVT div_U1211 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_36_), .Y(div_io_resp_bits_data[36]) );
  AO22X1_LVT div_U1210 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n206), .A4(div_result_35_), .Y(div_io_resp_bits_data[35]) );
  AO22X1_LVT div_U1209 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_34_), .Y(div_io_resp_bits_data[34]) );
  AO22X1_LVT div_U1208 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_33_), .Y(div_io_resp_bits_data[33]) );
  AO22X1_LVT div_U1207 ( .A1(div_n156), .A2(div_io_resp_bits_data[31]), .A3(
        div_n242), .A4(div_result_32_), .Y(div_io_resp_bits_data[32]) );
  AO22X1_LVT div_U1206 ( .A1(div_n146), .A2(div_result_62_), .A3(div_n209), 
        .A4(div_result_30_), .Y(div_io_resp_bits_data[30]) );
  AO22X1_LVT div_U1205 ( .A1(div_n146), .A2(div_result_34_), .A3(div_n209), 
        .A4(div_result_2_), .Y(div_io_resp_bits_data[2]) );
  AO22X1_LVT div_U1204 ( .A1(div_n146), .A2(div_result_61_), .A3(div_n209), 
        .A4(div_result_29_), .Y(div_io_resp_bits_data[29]) );
  AO22X1_LVT div_U1203 ( .A1(div_n146), .A2(div_result_60_), .A3(div_n209), 
        .A4(div_result_28_), .Y(div_io_resp_bits_data[28]) );
  AO22X1_LVT div_U1202 ( .A1(div_n146), .A2(div_result_59_), .A3(div_n209), 
        .A4(div_result_27_), .Y(div_io_resp_bits_data[27]) );
  AO22X1_LVT div_U1201 ( .A1(div_n146), .A2(div_result_58_), .A3(div_n209), 
        .A4(div_result_26_), .Y(div_io_resp_bits_data[26]) );
  AO22X1_LVT div_U1200 ( .A1(div_n146), .A2(div_result_57_), .A3(div_n209), 
        .A4(div_result_25_), .Y(div_io_resp_bits_data[25]) );
  AO22X1_LVT div_U1199 ( .A1(div_n146), .A2(div_result_56_), .A3(div_n209), 
        .A4(div_result_24_), .Y(div_io_resp_bits_data[24]) );
  AO22X1_LVT div_U1198 ( .A1(div_n146), .A2(div_result_55_), .A3(div_n209), 
        .A4(div_result_23_), .Y(div_io_resp_bits_data[23]) );
  AO22X1_LVT div_U1197 ( .A1(div_n146), .A2(div_result_53_), .A3(div_n209), 
        .A4(div_result_21_), .Y(div_io_resp_bits_data[21]) );
  AO22X1_LVT div_U1196 ( .A1(div_n146), .A2(div_result_52_), .A3(div_n209), 
        .A4(div_result_20_), .Y(div_io_resp_bits_data[20]) );
  AO22X1_LVT div_U1195 ( .A1(div_n146), .A2(div_result_33_), .A3(div_n209), 
        .A4(div_result_1_), .Y(div_io_resp_bits_data[1]) );
  AO22X1_LVT div_U1194 ( .A1(div_n146), .A2(div_result_51_), .A3(div_n209), 
        .A4(div_result_19_), .Y(div_io_resp_bits_data[19]) );
  AO22X1_LVT div_U1193 ( .A1(div_n146), .A2(div_result_50_), .A3(div_n209), 
        .A4(div_result_18_), .Y(div_io_resp_bits_data[18]) );
  AO22X1_LVT div_U1192 ( .A1(div_n146), .A2(div_result_49_), .A3(div_n209), 
        .A4(div_result_17_), .Y(div_io_resp_bits_data[17]) );
  AO22X1_LVT div_U1191 ( .A1(div_n146), .A2(div_result_48_), .A3(div_n209), 
        .A4(div_result_16_), .Y(div_io_resp_bits_data[16]) );
  AO22X1_LVT div_U1190 ( .A1(div_n146), .A2(div_result_47_), .A3(div_n209), 
        .A4(div_result_15_), .Y(div_io_resp_bits_data[15]) );
  AO22X1_LVT div_U1189 ( .A1(div_n146), .A2(div_result_46_), .A3(div_n209), 
        .A4(div_result_14_), .Y(div_io_resp_bits_data[14]) );
  AO22X1_LVT div_U1188 ( .A1(div_n146), .A2(div_result_45_), .A3(div_n209), 
        .A4(div_result_13_), .Y(div_io_resp_bits_data[13]) );
  AO22X1_LVT div_U1187 ( .A1(div_n146), .A2(div_result_44_), .A3(div_n209), 
        .A4(div_result_12_), .Y(div_io_resp_bits_data[12]) );
  AO22X1_LVT div_U1186 ( .A1(div_n146), .A2(div_result_42_), .A3(div_n209), 
        .A4(div_result_10_), .Y(div_io_resp_bits_data[10]) );
  AO22X1_LVT div_U1185 ( .A1(div_n146), .A2(div_result_32_), .A3(div_n209), 
        .A4(div_result_0_), .Y(div_io_resp_bits_data[0]) );
  NAND2X0_LVT div_U1184 ( .A1(div_n1002), .A2(div_n990), .Y(div_n_T_429[4]) );
  NAND2X0_LVT div_U1183 ( .A1(div_n976), .A2(div_n975), .Y(div_n990) );
  OR3X1_LVT div_U1182 ( .A1(div_n974), .A2(div_n973), .A3(div_n997), .Y(
        div_n975) );
  NAND2X0_LVT div_U1181 ( .A1(div_n969), .A2(div_n968), .Y(div_n_T_272[4]) );
  NAND4X0_LVT div_U1180 ( .A1(div_n961), .A2(div_n960), .A3(div_n959), .A4(
        div_n958), .Y(div_n_T_272[2]) );
  AO221X1_LVT div_U1179 ( .A1(div_n761), .A2(div_n760), .A3(div_n761), .A4(
        div_n962), .A5(div_n957), .Y(div_n958) );
  AO221X1_LVT div_U1178 ( .A1(div_n767), .A2(div_n768), .A3(div_n767), .A4(
        div_n966), .A5(div_n956), .Y(div_n959) );
  AO221X1_LVT div_U1177 ( .A1(div_n764), .A2(div_n765), .A3(div_n764), .A4(
        div_n964), .A5(div_n_T_273_5_), .Y(div_n960) );
  OA21X1_LVT div_U1176 ( .A1(div_n770), .A2(div_n967), .A3(div_n769), .Y(
        div_n961) );
  OR3X1_LVT div_U1175 ( .A1(div_n955), .A2(div_n954), .A3(div_n953), .Y(
        div_n_T_272[1]) );
  AO22X1_LVT div_U1174 ( .A1(div_n969), .A2(div_n952), .A3(div_n763), .A4(
        div_n951), .Y(div_n953) );
  AO221X1_LVT div_U1173 ( .A1(div_n963), .A2(div_n950), .A3(div_n963), .A4(
        div_n949), .A5(div_n948), .Y(div_n954) );
  OR3X1_LVT div_U1172 ( .A1(div_n955), .A2(div_n947), .A3(div_n946), .Y(
        div_n_T_272[0]) );
  AO22X1_LVT div_U1171 ( .A1(div_n969), .A2(div_n945), .A3(div_n963), .A4(
        div_n944), .Y(div_n946) );
  NAND4X0_LVT div_U1170 ( .A1(div_n759), .A2(div_n943), .A3(div_n942), .A4(
        div_n941), .Y(div_n944) );
  NAND2X0_LVT div_U1169 ( .A1(div_n965), .A2(div_n940), .Y(div_n957) );
  NAND4X0_LVT div_U1168 ( .A1(div_n762), .A2(div_n939), .A3(div_n938), .A4(
        div_n937), .Y(div_n945) );
  NAND4X0_LVT div_U1167 ( .A1(div_n936), .A2(div_n935), .A3(div_n934), .A4(
        div_n933), .Y(div_n947) );
  NAND3X0_LVT div_U1166 ( .A1(div_n969), .A2(div_n766), .A3(div_n932), .Y(
        div_n_T_273_5_) );
  OR2X1_LVT div_U1165 ( .A1(div_n930), .A2(div_n929), .Y(div_N521) );
  AO22X1_LVT div_U1164 ( .A1(div_n783), .A2(div_n_T_65[69]), .A3(div_n226), 
        .A4(div_subtractor_61_), .Y(div_n929) );
  AO22X1_LVT div_U1163 ( .A1(div_n157), .A2(div_n_T_442[126]), .A3(div_n931), 
        .A4(div_n_T_51_124_), .Y(div_n930) );
  OR2X1_LVT div_U1162 ( .A1(div_n928), .A2(div_n927), .Y(div_N520) );
  AO22X1_LVT div_U1161 ( .A1(div_n783), .A2(div_n_T_65[68]), .A3(div_n226), 
        .A4(div_subtractor_60_), .Y(div_n927) );
  AO22X1_LVT div_U1160 ( .A1(div_n157), .A2(div_n_T_442[125]), .A3(div_n931), 
        .A4(div_n_T_51_123_), .Y(div_n928) );
  OR2X1_LVT div_U1159 ( .A1(div_n926), .A2(div_n925), .Y(div_N519) );
  AO22X1_LVT div_U1158 ( .A1(div_n783), .A2(div_n_T_65[67]), .A3(div_n226), 
        .A4(div_subtractor_59_), .Y(div_n925) );
  AO22X1_LVT div_U1157 ( .A1(div_n157), .A2(div_n_T_442[124]), .A3(div_n931), 
        .A4(div_n_T_51_122_), .Y(div_n926) );
  OR2X1_LVT div_U1156 ( .A1(div_n924), .A2(div_n923), .Y(div_N518) );
  AO22X1_LVT div_U1155 ( .A1(div_n783), .A2(div_n_T_65[66]), .A3(div_n226), 
        .A4(div_subtractor_58_), .Y(div_n923) );
  AO22X1_LVT div_U1154 ( .A1(div_n157), .A2(div_n_T_442[123]), .A3(div_n931), 
        .A4(div_n_T_51_121_), .Y(div_n924) );
  OR2X1_LVT div_U1153 ( .A1(div_n922), .A2(div_n921), .Y(div_N517) );
  AO22X1_LVT div_U1152 ( .A1(div_n783), .A2(div_n_T_65[65]), .A3(div_n226), 
        .A4(div_subtractor_57_), .Y(div_n921) );
  AO22X1_LVT div_U1151 ( .A1(div_n225), .A2(div_n_T_442[122]), .A3(div_n931), 
        .A4(div_n_T_51_120_), .Y(div_n922) );
  OR2X1_LVT div_U1150 ( .A1(div_n920), .A2(div_n919), .Y(div_N516) );
  AO22X1_LVT div_U1149 ( .A1(div_n783), .A2(div_n_T_65[64]), .A3(div_n226), 
        .A4(div_subtractor_56_), .Y(div_n919) );
  AO22X1_LVT div_U1148 ( .A1(div_n225), .A2(div_n_T_442[121]), .A3(div_n931), 
        .A4(div_n_T_51_119_), .Y(div_n920) );
  OR2X1_LVT div_U1147 ( .A1(div_n918), .A2(div_n917), .Y(div_N515) );
  AO22X1_LVT div_U1146 ( .A1(div_n783), .A2(div_n_T_65[63]), .A3(div_n226), 
        .A4(div_subtractor_55_), .Y(div_n917) );
  AO22X1_LVT div_U1145 ( .A1(div_n225), .A2(div_n_T_442[120]), .A3(div_n931), 
        .A4(div_n_T_51_118_), .Y(div_n918) );
  OR2X1_LVT div_U1144 ( .A1(div_n916), .A2(div_n915), .Y(div_N514) );
  AO22X1_LVT div_U1143 ( .A1(div_n783), .A2(div_n_T_65[62]), .A3(div_n226), 
        .A4(div_subtractor_54_), .Y(div_n915) );
  AO22X1_LVT div_U1142 ( .A1(div_n225), .A2(div_n_T_442[119]), .A3(div_n931), 
        .A4(div_n_T_51_117_), .Y(div_n916) );
  OR2X1_LVT div_U1141 ( .A1(div_n914), .A2(div_n913), .Y(div_N513) );
  AO22X1_LVT div_U1140 ( .A1(div_n783), .A2(div_n_T_65[61]), .A3(div_n226), 
        .A4(div_subtractor_53_), .Y(div_n913) );
  AO22X1_LVT div_U1139 ( .A1(div_n157), .A2(div_n_T_442[118]), .A3(div_n931), 
        .A4(div_n_T_51_116_), .Y(div_n914) );
  OR2X1_LVT div_U1138 ( .A1(div_n912), .A2(div_n911), .Y(div_N512) );
  AO22X1_LVT div_U1137 ( .A1(div_n783), .A2(div_n_T_65[60]), .A3(div_n226), 
        .A4(div_subtractor_52_), .Y(div_n911) );
  AO22X1_LVT div_U1136 ( .A1(div_n225), .A2(div_n_T_442[117]), .A3(div_n931), 
        .A4(div_n_T_51_115_), .Y(div_n912) );
  OR2X1_LVT div_U1135 ( .A1(div_n910), .A2(div_n909), .Y(div_N511) );
  AO22X1_LVT div_U1134 ( .A1(div_n783), .A2(div_n_T_65[59]), .A3(div_n226), 
        .A4(div_subtractor_51_), .Y(div_n909) );
  AO22X1_LVT div_U1133 ( .A1(div_n225), .A2(div_n_T_442[116]), .A3(div_n931), 
        .A4(div_n_T_51_114_), .Y(div_n910) );
  OR2X1_LVT div_U1132 ( .A1(div_n908), .A2(div_n907), .Y(div_N510) );
  AO22X1_LVT div_U1131 ( .A1(div_n783), .A2(div_n_T_65[58]), .A3(div_n226), 
        .A4(div_subtractor_50_), .Y(div_n907) );
  AO22X1_LVT div_U1130 ( .A1(div_n225), .A2(div_n_T_442[115]), .A3(div_n931), 
        .A4(div_n_T_51_113_), .Y(div_n908) );
  OR2X1_LVT div_U1129 ( .A1(div_n906), .A2(div_n905), .Y(div_N509) );
  AO22X1_LVT div_U1128 ( .A1(div_n783), .A2(div_n_T_65[57]), .A3(div_n226), 
        .A4(div_subtractor_49_), .Y(div_n905) );
  AO22X1_LVT div_U1127 ( .A1(div_n225), .A2(div_n_T_442[114]), .A3(div_n931), 
        .A4(div_n_T_51_112_), .Y(div_n906) );
  OR2X1_LVT div_U1126 ( .A1(div_n904), .A2(div_n903), .Y(div_N508) );
  AO22X1_LVT div_U1125 ( .A1(div_n783), .A2(div_n_T_65[56]), .A3(div_n226), 
        .A4(div_subtractor_48_), .Y(div_n903) );
  AO22X1_LVT div_U1124 ( .A1(div_n225), .A2(div_n_T_442[113]), .A3(div_n931), 
        .A4(div_n_T_51_111_), .Y(div_n904) );
  OR2X1_LVT div_U1123 ( .A1(div_n902), .A2(div_n901), .Y(div_N507) );
  AO22X1_LVT div_U1122 ( .A1(div_n783), .A2(div_n_T_65[55]), .A3(div_n226), 
        .A4(div_subtractor_47_), .Y(div_n901) );
  AO22X1_LVT div_U1121 ( .A1(div_n225), .A2(div_n_T_442[112]), .A3(div_n931), 
        .A4(div_n_T_51_110_), .Y(div_n902) );
  OR2X1_LVT div_U1120 ( .A1(div_n900), .A2(div_n899), .Y(div_N506) );
  AO22X1_LVT div_U1119 ( .A1(div_n783), .A2(div_n_T_65[54]), .A3(div_n226), 
        .A4(div_subtractor_46_), .Y(div_n899) );
  AO22X1_LVT div_U1118 ( .A1(div_n157), .A2(div_n_T_442[111]), .A3(div_n931), 
        .A4(div_n_T_51_109_), .Y(div_n900) );
  OR2X1_LVT div_U1117 ( .A1(div_n898), .A2(div_n897), .Y(div_N505) );
  AO22X1_LVT div_U1116 ( .A1(div_n783), .A2(div_n_T_65[53]), .A3(div_n226), 
        .A4(div_subtractor_45_), .Y(div_n897) );
  AO22X1_LVT div_U1115 ( .A1(div_n225), .A2(div_n_T_442[110]), .A3(div_n931), 
        .A4(div_n_T_51_108_), .Y(div_n898) );
  OR2X1_LVT div_U1114 ( .A1(div_n896), .A2(div_n895), .Y(div_N504) );
  AO22X1_LVT div_U1113 ( .A1(div_n783), .A2(div_n_T_65[52]), .A3(div_n226), 
        .A4(div_subtractor_44_), .Y(div_n895) );
  AO22X1_LVT div_U1112 ( .A1(div_n225), .A2(div_n_T_442[109]), .A3(div_n931), 
        .A4(div_n_T_51_107_), .Y(div_n896) );
  OR2X1_LVT div_U1111 ( .A1(div_n894), .A2(div_n893), .Y(div_N503) );
  AO22X1_LVT div_U1110 ( .A1(div_n783), .A2(div_n_T_65[51]), .A3(div_n226), 
        .A4(div_subtractor_43_), .Y(div_n893) );
  AO22X1_LVT div_U1109 ( .A1(div_n225), .A2(div_n_T_442[108]), .A3(div_n931), 
        .A4(div_n_T_51_106_), .Y(div_n894) );
  OR2X1_LVT div_U1108 ( .A1(div_n892), .A2(div_n891), .Y(div_N502) );
  AO22X1_LVT div_U1107 ( .A1(div_n783), .A2(div_n_T_65[50]), .A3(div_n226), 
        .A4(div_subtractor_42_), .Y(div_n891) );
  AO22X1_LVT div_U1106 ( .A1(div_n157), .A2(div_n_T_442[107]), .A3(div_n931), 
        .A4(div_n_T_51_105_), .Y(div_n892) );
  OR2X1_LVT div_U1105 ( .A1(div_n890), .A2(div_n889), .Y(div_N501) );
  AO22X1_LVT div_U1104 ( .A1(div_n783), .A2(div_n_T_65[49]), .A3(div_n226), 
        .A4(div_subtractor_41_), .Y(div_n889) );
  AO22X1_LVT div_U1103 ( .A1(div_n225), .A2(div_n_T_442[106]), .A3(div_n931), 
        .A4(div_n_T_51_104_), .Y(div_n890) );
  OR2X1_LVT div_U1102 ( .A1(div_n888), .A2(div_n887), .Y(div_N500) );
  AO22X1_LVT div_U1101 ( .A1(div_n783), .A2(div_n_T_65[48]), .A3(div_n226), 
        .A4(div_subtractor_40_), .Y(div_n887) );
  AO22X1_LVT div_U1100 ( .A1(div_n225), .A2(div_n_T_442[105]), .A3(div_n931), 
        .A4(div_n_T_51_103_), .Y(div_n888) );
  OR2X1_LVT div_U1099 ( .A1(div_n886), .A2(div_n885), .Y(div_N499) );
  AO22X1_LVT div_U1098 ( .A1(div_n783), .A2(div_n_T_65[47]), .A3(div_n226), 
        .A4(div_subtractor_39_), .Y(div_n885) );
  AO22X1_LVT div_U1097 ( .A1(div_n225), .A2(div_n_T_442[104]), .A3(div_n931), 
        .A4(div_n_T_51_102_), .Y(div_n886) );
  OR2X1_LVT div_U1096 ( .A1(div_n884), .A2(div_n883), .Y(div_N498) );
  AO22X1_LVT div_U1095 ( .A1(div_n783), .A2(div_n_T_65[46]), .A3(div_n226), 
        .A4(div_subtractor_38_), .Y(div_n883) );
  AO22X1_LVT div_U1094 ( .A1(div_n225), .A2(div_n_T_442[103]), .A3(div_n931), 
        .A4(div_n_T_51_101_), .Y(div_n884) );
  OR2X1_LVT div_U1093 ( .A1(div_n882), .A2(div_n881), .Y(div_N497) );
  AO22X1_LVT div_U1092 ( .A1(div_n783), .A2(div_n_T_65[45]), .A3(div_n226), 
        .A4(div_subtractor_37_), .Y(div_n881) );
  AO22X1_LVT div_U1091 ( .A1(div_n157), .A2(div_n_T_442[102]), .A3(div_n931), 
        .A4(div_n_T_51_100_), .Y(div_n882) );
  OR2X1_LVT div_U1090 ( .A1(div_n880), .A2(div_n879), .Y(div_N496) );
  AO22X1_LVT div_U1089 ( .A1(div_n783), .A2(div_n_T_65[44]), .A3(div_n226), 
        .A4(div_subtractor_36_), .Y(div_n879) );
  AO22X1_LVT div_U1088 ( .A1(div_n225), .A2(div_n_T_442[101]), .A3(div_n931), 
        .A4(div_n_T_51_99_), .Y(div_n880) );
  OR2X1_LVT div_U1087 ( .A1(div_n878), .A2(div_n877), .Y(div_N495) );
  AO22X1_LVT div_U1086 ( .A1(div_n783), .A2(div_n_T_65[43]), .A3(div_n226), 
        .A4(div_subtractor_35_), .Y(div_n877) );
  AO22X1_LVT div_U1085 ( .A1(div_n225), .A2(div_n_T_442[100]), .A3(div_n931), 
        .A4(div_n_T_51_98_), .Y(div_n878) );
  OR2X1_LVT div_U1084 ( .A1(div_n876), .A2(div_n875), .Y(div_N494) );
  AO22X1_LVT div_U1083 ( .A1(div_n783), .A2(div_n_T_65[42]), .A3(div_n226), 
        .A4(div_subtractor_34_), .Y(div_n875) );
  AO22X1_LVT div_U1082 ( .A1(div_n157), .A2(div_n_T_442[99]), .A3(div_n931), 
        .A4(div_n_T_51_97_), .Y(div_n876) );
  OR2X1_LVT div_U1081 ( .A1(div_n874), .A2(div_n873), .Y(div_N492) );
  AO22X1_LVT div_U1080 ( .A1(div_n783), .A2(div_n_T_65[41]), .A3(div_n226), 
        .A4(div_subtractor_33_), .Y(div_n873) );
  AO22X1_LVT div_U1079 ( .A1(div_n225), .A2(div_n_T_442[98]), .A3(div_n931), 
        .A4(div_n_T_51_96_), .Y(div_n874) );
  OR2X1_LVT div_U1078 ( .A1(div_n872), .A2(div_n871), .Y(div_N491) );
  AO22X1_LVT div_U1077 ( .A1(div_n783), .A2(div_n_T_65[40]), .A3(div_n226), 
        .A4(div_subtractor_32_), .Y(div_n871) );
  AO22X1_LVT div_U1076 ( .A1(div_n225), .A2(div_n_T_442[97]), .A3(div_n931), 
        .A4(div_n_T_51_95_), .Y(div_n872) );
  OR2X1_LVT div_U1075 ( .A1(div_n870), .A2(div_n869), .Y(div_N490) );
  AO22X1_LVT div_U1074 ( .A1(div_n783), .A2(div_n_T_65[39]), .A3(div_n226), 
        .A4(div_subtractor_31_), .Y(div_n869) );
  AO22X1_LVT div_U1073 ( .A1(div_n157), .A2(div_n_T_442[96]), .A3(div_n931), 
        .A4(div_n_T_51_94_), .Y(div_n870) );
  OR2X1_LVT div_U1072 ( .A1(div_n868), .A2(div_n867), .Y(div_N489) );
  AO22X1_LVT div_U1071 ( .A1(div_n783), .A2(div_n_T_65[38]), .A3(div_n226), 
        .A4(div_subtractor_30_), .Y(div_n867) );
  AO22X1_LVT div_U1070 ( .A1(div_n225), .A2(div_n_T_442[95]), .A3(div_n931), 
        .A4(div_n_T_51_93_), .Y(div_n868) );
  OR2X1_LVT div_U1069 ( .A1(div_n866), .A2(div_n865), .Y(div_N488) );
  AO22X1_LVT div_U1068 ( .A1(div_n783), .A2(div_n_T_65[37]), .A3(div_n226), 
        .A4(div_subtractor_29_), .Y(div_n865) );
  AO22X1_LVT div_U1067 ( .A1(div_n225), .A2(div_n_T_442[94]), .A3(div_n931), 
        .A4(div_n_T_51_92_), .Y(div_n866) );
  OR2X1_LVT div_U1066 ( .A1(div_n864), .A2(div_n863), .Y(div_N487) );
  AO22X1_LVT div_U1065 ( .A1(div_n783), .A2(div_n_T_65[36]), .A3(div_n226), 
        .A4(div_subtractor_28_), .Y(div_n863) );
  AO22X1_LVT div_U1064 ( .A1(div_n157), .A2(div_n_T_442[93]), .A3(div_n931), 
        .A4(div_n_T_51_91_), .Y(div_n864) );
  OR2X1_LVT div_U1063 ( .A1(div_n862), .A2(div_n861), .Y(div_N486) );
  AO22X1_LVT div_U1062 ( .A1(div_n783), .A2(div_n_T_65[35]), .A3(div_n226), 
        .A4(div_subtractor_27_), .Y(div_n861) );
  AO22X1_LVT div_U1061 ( .A1(div_n225), .A2(div_n_T_442[92]), .A3(div_n931), 
        .A4(div_n_T_51_90_), .Y(div_n862) );
  OR2X1_LVT div_U1060 ( .A1(div_n860), .A2(div_n859), .Y(div_N485) );
  AO22X1_LVT div_U1059 ( .A1(div_n783), .A2(div_n_T_65[34]), .A3(div_n226), 
        .A4(div_subtractor_26_), .Y(div_n859) );
  AO22X1_LVT div_U1058 ( .A1(div_n225), .A2(div_n_T_442[91]), .A3(div_n931), 
        .A4(div_n_T_51_89_), .Y(div_n860) );
  OR2X1_LVT div_U1057 ( .A1(div_n858), .A2(div_n857), .Y(div_N484) );
  AO22X1_LVT div_U1056 ( .A1(div_n783), .A2(div_n_T_65[33]), .A3(div_n226), 
        .A4(div_subtractor_25_), .Y(div_n857) );
  AO22X1_LVT div_U1055 ( .A1(div_n157), .A2(div_n_T_442[90]), .A3(div_n931), 
        .A4(div_n_T_51_88_), .Y(div_n858) );
  OR2X1_LVT div_U1054 ( .A1(div_n856), .A2(div_n855), .Y(div_N483) );
  AO22X1_LVT div_U1053 ( .A1(div_n783), .A2(div_n_T_65[32]), .A3(div_n226), 
        .A4(div_subtractor_24_), .Y(div_n855) );
  AO22X1_LVT div_U1052 ( .A1(div_n225), .A2(div_n_T_442[89]), .A3(div_n931), 
        .A4(div_n_T_51_87_), .Y(div_n856) );
  OR2X1_LVT div_U1051 ( .A1(div_n854), .A2(div_n853), .Y(div_N482) );
  AO22X1_LVT div_U1050 ( .A1(div_n783), .A2(div_n_T_65[31]), .A3(div_n226), 
        .A4(div_subtractor_23_), .Y(div_n853) );
  AO22X1_LVT div_U1049 ( .A1(div_n157), .A2(div_n_T_442[88]), .A3(div_n931), 
        .A4(div_n_T_51_86_), .Y(div_n854) );
  OR2X1_LVT div_U1048 ( .A1(div_n852), .A2(div_n851), .Y(div_N481) );
  AO22X1_LVT div_U1047 ( .A1(div_n783), .A2(div_n_T_65[30]), .A3(div_n226), 
        .A4(div_subtractor_22_), .Y(div_n851) );
  AO22X1_LVT div_U1046 ( .A1(div_n225), .A2(div_n_T_442[87]), .A3(div_n931), 
        .A4(div_n_T_51_85_), .Y(div_n852) );
  OR2X1_LVT div_U1045 ( .A1(div_n850), .A2(div_n849), .Y(div_N480) );
  AO22X1_LVT div_U1044 ( .A1(div_n783), .A2(div_n_T_65[29]), .A3(div_n226), 
        .A4(div_subtractor_21_), .Y(div_n849) );
  AO22X1_LVT div_U1043 ( .A1(div_n225), .A2(div_n_T_442[86]), .A3(div_n931), 
        .A4(div_n_T_51_84_), .Y(div_n850) );
  OR2X1_LVT div_U1042 ( .A1(div_n848), .A2(div_n847), .Y(div_N479) );
  AO22X1_LVT div_U1041 ( .A1(div_n783), .A2(div_n_T_65[28]), .A3(div_n226), 
        .A4(div_subtractor_20_), .Y(div_n847) );
  AO22X1_LVT div_U1040 ( .A1(div_n225), .A2(div_n_T_442[85]), .A3(div_n931), 
        .A4(div_n_T_51_83_), .Y(div_n848) );
  OR2X1_LVT div_U1039 ( .A1(div_n846), .A2(div_n845), .Y(div_N478) );
  AO22X1_LVT div_U1038 ( .A1(div_n783), .A2(div_n_T_65[27]), .A3(div_n226), 
        .A4(div_subtractor_19_), .Y(div_n845) );
  AO22X1_LVT div_U1037 ( .A1(div_n225), .A2(div_n_T_442[84]), .A3(div_n931), 
        .A4(div_n_T_51_82_), .Y(div_n846) );
  OR2X1_LVT div_U1036 ( .A1(div_n844), .A2(div_n843), .Y(div_N477) );
  AO22X1_LVT div_U1035 ( .A1(div_n783), .A2(div_n_T_65[26]), .A3(div_n226), 
        .A4(div_subtractor_18_), .Y(div_n843) );
  AO22X1_LVT div_U1034 ( .A1(div_n225), .A2(div_n_T_442[83]), .A3(div_n931), 
        .A4(div_n_T_51_81_), .Y(div_n844) );
  OR2X1_LVT div_U1033 ( .A1(div_n842), .A2(div_n841), .Y(div_N476) );
  AO22X1_LVT div_U1032 ( .A1(div_n783), .A2(div_n_T_65[25]), .A3(div_n226), 
        .A4(div_subtractor_17_), .Y(div_n841) );
  AO22X1_LVT div_U1031 ( .A1(div_n225), .A2(div_n_T_442[82]), .A3(div_n931), 
        .A4(div_n_T_51_80_), .Y(div_n842) );
  OR2X1_LVT div_U1030 ( .A1(div_n840), .A2(div_n839), .Y(div_N475) );
  AO22X1_LVT div_U1029 ( .A1(div_n783), .A2(div_n_T_65[24]), .A3(div_n226), 
        .A4(div_subtractor_16_), .Y(div_n839) );
  AO22X1_LVT div_U1028 ( .A1(div_n225), .A2(div_n_T_442[81]), .A3(div_n931), 
        .A4(div_n_T_51_79_), .Y(div_n840) );
  OR2X1_LVT div_U1027 ( .A1(div_n838), .A2(div_n837), .Y(div_N474) );
  AO22X1_LVT div_U1026 ( .A1(div_n783), .A2(div_n_T_65[23]), .A3(div_n226), 
        .A4(div_subtractor_15_), .Y(div_n837) );
  AO22X1_LVT div_U1025 ( .A1(div_n225), .A2(div_n_T_442[80]), .A3(div_n931), 
        .A4(div_n_T_51_78_), .Y(div_n838) );
  OR2X1_LVT div_U1024 ( .A1(div_n836), .A2(div_n835), .Y(div_N473) );
  AO22X1_LVT div_U1023 ( .A1(div_n783), .A2(div_n_T_65[22]), .A3(div_n226), 
        .A4(div_subtractor_14_), .Y(div_n835) );
  AO22X1_LVT div_U1022 ( .A1(div_n157), .A2(div_n_T_442[79]), .A3(div_n931), 
        .A4(div_n_T_51_77_), .Y(div_n836) );
  OR2X1_LVT div_U1021 ( .A1(div_n834), .A2(div_n833), .Y(div_N472) );
  AO22X1_LVT div_U1020 ( .A1(div_n783), .A2(div_n_T_65[21]), .A3(div_n226), 
        .A4(div_subtractor_13_), .Y(div_n833) );
  AO22X1_LVT div_U1019 ( .A1(div_n225), .A2(div_n_T_442[78]), .A3(div_n931), 
        .A4(div_n_T_51_76_), .Y(div_n834) );
  OR2X1_LVT div_U1018 ( .A1(div_n832), .A2(div_n831), .Y(div_N471) );
  AO22X1_LVT div_U1017 ( .A1(div_n783), .A2(div_n_T_65[20]), .A3(div_n226), 
        .A4(div_subtractor_12_), .Y(div_n831) );
  AO22X1_LVT div_U1016 ( .A1(div_n225), .A2(div_n_T_442[77]), .A3(div_n931), 
        .A4(div_n_T_51_75_), .Y(div_n832) );
  OR2X1_LVT div_U1015 ( .A1(div_n830), .A2(div_n829), .Y(div_N470) );
  AO22X1_LVT div_U1014 ( .A1(div_n783), .A2(div_n_T_65[19]), .A3(div_n226), 
        .A4(div_subtractor_11_), .Y(div_n829) );
  AO22X1_LVT div_U1013 ( .A1(div_n225), .A2(div_n_T_442[76]), .A3(div_n931), 
        .A4(div_n_T_51_74_), .Y(div_n830) );
  OR2X1_LVT div_U1012 ( .A1(div_n828), .A2(div_n827), .Y(div_N469) );
  AO22X1_LVT div_U1011 ( .A1(div_n783), .A2(div_n_T_65[18]), .A3(div_n226), 
        .A4(div_subtractor_10_), .Y(div_n827) );
  AO22X1_LVT div_U1010 ( .A1(div_n225), .A2(div_n_T_442[75]), .A3(div_n931), 
        .A4(div_n_T_51_73_), .Y(div_n828) );
  OR2X1_LVT div_U1009 ( .A1(div_n826), .A2(div_n825), .Y(div_N468) );
  AO22X1_LVT div_U1008 ( .A1(div_n783), .A2(div_n_T_65[17]), .A3(div_n226), 
        .A4(div_subtractor_9_), .Y(div_n825) );
  AO22X1_LVT div_U1007 ( .A1(div_n157), .A2(div_n_T_442[74]), .A3(div_n931), 
        .A4(div_n_T_51_72_), .Y(div_n826) );
  OR2X1_LVT div_U1006 ( .A1(div_n824), .A2(div_n823), .Y(div_N467) );
  AO22X1_LVT div_U1005 ( .A1(div_n783), .A2(div_n_T_65[16]), .A3(div_n226), 
        .A4(div_subtractor_8_), .Y(div_n823) );
  AO22X1_LVT div_U1004 ( .A1(div_n225), .A2(div_n_T_442[73]), .A3(div_n931), 
        .A4(div_n_T_51_71_), .Y(div_n824) );
  OR2X1_LVT div_U1003 ( .A1(div_n822), .A2(div_n821), .Y(div_N466) );
  AO22X1_LVT div_U1002 ( .A1(div_n783), .A2(div_n_T_65[15]), .A3(div_n226), 
        .A4(div_subtractor_7_), .Y(div_n821) );
  AO22X1_LVT div_U1001 ( .A1(div_n225), .A2(div_n_T_442[72]), .A3(div_n931), 
        .A4(div_n_T_51_70_), .Y(div_n822) );
  OR2X1_LVT div_U1000 ( .A1(div_n820), .A2(div_n819), .Y(div_N465) );
  AO22X1_LVT div_U999 ( .A1(div_n783), .A2(div_n_T_65[14]), .A3(div_n226), 
        .A4(div_subtractor_6_), .Y(div_n819) );
  AO22X1_LVT div_U998 ( .A1(div_n225), .A2(div_n_T_442[71]), .A3(div_n931), 
        .A4(div_n_T_51_69_), .Y(div_n820) );
  OR2X1_LVT div_U997 ( .A1(div_n818), .A2(div_n817), .Y(div_N464) );
  AO22X1_LVT div_U996 ( .A1(div_n783), .A2(div_n_T_65[13]), .A3(div_n226), 
        .A4(div_subtractor_5_), .Y(div_n817) );
  AO22X1_LVT div_U995 ( .A1(div_n225), .A2(div_n_T_442[70]), .A3(div_n931), 
        .A4(div_n_T_51_68_), .Y(div_n818) );
  OR2X1_LVT div_U994 ( .A1(div_n816), .A2(div_n815), .Y(div_N463) );
  AO22X1_LVT div_U993 ( .A1(div_n783), .A2(div_n_T_65[12]), .A3(div_n226), 
        .A4(div_subtractor_4_), .Y(div_n815) );
  AO22X1_LVT div_U992 ( .A1(div_n225), .A2(div_n_T_442[69]), .A3(div_n931), 
        .A4(div_n_T_51_67_), .Y(div_n816) );
  OR2X1_LVT div_U991 ( .A1(div_n814), .A2(div_n813), .Y(div_N462) );
  AO22X1_LVT div_U990 ( .A1(div_n783), .A2(div_n_T_65[11]), .A3(div_n226), 
        .A4(div_subtractor_3_), .Y(div_n813) );
  AO22X1_LVT div_U989 ( .A1(div_n225), .A2(div_n_T_442[68]), .A3(div_n931), 
        .A4(div_n_T_51_66_), .Y(div_n814) );
  OR2X1_LVT div_U988 ( .A1(div_n812), .A2(div_n811), .Y(div_N461) );
  AO22X1_LVT div_U987 ( .A1(div_n783), .A2(div_n_T_65[10]), .A3(div_n226), 
        .A4(div_subtractor_2_), .Y(div_n811) );
  AO22X1_LVT div_U986 ( .A1(div_n225), .A2(div_n_T_442[67]), .A3(div_n931), 
        .A4(div_n_T_51_65_), .Y(div_n812) );
  OR2X1_LVT div_U985 ( .A1(div_n810), .A2(div_n809), .Y(div_N460) );
  AO22X1_LVT div_U984 ( .A1(div_n783), .A2(div_n_T_65[9]), .A3(div_n226), .A4(
        div_subtractor_1_), .Y(div_n809) );
  AO22X1_LVT div_U983 ( .A1(div_n157), .A2(div_n_T_442[66]), .A3(
        div_n_T_51_64_), .A4(div_n931), .Y(div_n810) );
  OR2X1_LVT div_U982 ( .A1(div_n808), .A2(div_n807), .Y(div_N459) );
  AO22X1_LVT div_U981 ( .A1(div_n783), .A2(div_n_T_65[8]), .A3(div_n226), .A4(
        div_subtractor_0_), .Y(div_n807) );
  AO22X1_LVT div_U980 ( .A1(div_n225), .A2(div_n_T_442[65]), .A3(div_n931), 
        .A4(div_n301), .Y(div_n808) );
  AO22X1_LVT div_U979 ( .A1(div_n806), .A2(div_n805), .A3(div_n225), .A4(
        div_n170), .Y(div_N299) );
  AO22X1_LVT div_U978 ( .A1(div_n_T_69_8_), .A2(div_n804), .A3(div_n197), .A4(
        div_n803), .Y(div_n806) );
  AO22X1_LVT div_U977 ( .A1(div_n802), .A2(div_n805), .A3(div_n225), .A4(
        div_n169), .Y(div_N298) );
  OA221X1_LVT div_U976 ( .A1(div_n_T_69_7_), .A2(div_n_T_69_6_), .A3(
        div_n_T_69_7_), .A4(div_n778), .A5(div_n804), .Y(div_n802) );
  AO22X1_LVT div_U975 ( .A1(div_n801), .A2(div_n805), .A3(div_n225), .A4(
        div_n168), .Y(div_N297) );
  AO22X1_LVT div_U974 ( .A1(div_n_T_69_6_), .A2(div_n800), .A3(div_n198), .A4(
        div_n778), .Y(div_n801) );
  NAND3X0_LVT div_U973 ( .A1(div_n799), .A2(div_n798), .A3(div_n797), .Y(
        div_N296) );
  NAND3X0_LVT div_U972 ( .A1(div_n235), .A2(div_n787), .A3(div_n784), .Y(
        div_n797) );
  NAND2X0_LVT div_U971 ( .A1(div_n225), .A2(div_n167), .Y(div_n799) );
  AO22X1_LVT div_U970 ( .A1(div_n_T_85_4_), .A2(div_n805), .A3(div_n157), .A4(
        div_n166), .Y(div_N295) );
  NAND2X0_LVT div_U969 ( .A1(div_n230), .A2(div_n200), .Y(div_n805) );
  NAND3X0_LVT div_U968 ( .A1(div_n_T_434_2_), .A2(div_n_T_434_1_), .A3(
        div_n791), .Y(div_n792) );
  AND4X1_LVT div_U967 ( .A1(div_n_T_434_3_), .A2(div_n_T_434_5_), .A3(
        div_n_T_434_4_), .A4(div_n_T_434_0_), .Y(div_n791) );
  NAND3X0_LVT div_U964 ( .A1(div_n_T_69_6_), .A2(div_n_T_69_7_), .A3(div_n778), 
        .Y(div_n804) );
  AO21X1_LVT div_U963 ( .A1(div_n754), .A2(div_divisor_63_), .A3(div_n235), 
        .Y(div_N322) );
  NAND3X0_LVT div_U962 ( .A1(div_n753), .A2(div_n752), .A3(div_n203), .Y(
        div_N282) );
  NAND2X0_LVT div_U961 ( .A1(div_n751), .A2(div_n199), .Y(div_N293) );
  INVX1_LVT div_U960 ( .A(div_n750), .Y(div_n751) );
  NAND3X0_LVT div_U959 ( .A1(div_n749), .A2(div_n277), .A3(div_n_T_51_17_), 
        .Y(div_n991) );
  NAND3X0_LVT div_U958 ( .A1(div_n273), .A2(div_n775), .A3(div_n_T_51_21_), 
        .Y(div_n992) );
  OA22X1_LVT div_U957 ( .A1(div_n181), .A2(div_n_T_51_30_), .A3(div_n748), 
        .A4(div_n739), .Y(div_n993) );
  NAND2X0_LVT div_U956 ( .A1(div_n268), .A2(div_n_T_51_25_), .Y(div_n739) );
  INVX1_LVT div_U955 ( .A(div_n776), .Y(div_n748) );
  AND2X1_LVT div_U954 ( .A1(div_n777), .A2(div_n775), .Y(div_n749) );
  NAND3X0_LVT div_U953 ( .A1(div_n742), .A2(div_n259), .A3(div_n_T_51_33_), 
        .Y(div_n987) );
  NAND3X0_LVT div_U952 ( .A1(div_n255), .A2(div_n741), .A3(div_n_T_51_37_), 
        .Y(div_n988) );
  OA22X1_LVT div_U951 ( .A1(div_n248), .A2(div_n_T_51_46_), .A3(div_n738), 
        .A4(div_n740), .Y(div_n989) );
  INVX1_LVT div_U950 ( .A(div_n771), .Y(div_n740) );
  NAND2X0_LVT div_U949 ( .A1(div_n251), .A2(div_n_T_51_41_), .Y(div_n738) );
  INVX1_LVT div_U948 ( .A(div_n998), .Y(div_n742) );
  INVX1_LVT div_U947 ( .A(div_n999), .Y(div_n741) );
  NAND3X0_LVT div_U946 ( .A1(div_n745), .A2(div_n_T_51_1_), .A3(div_n208), .Y(
        div_n984) );
  NAND3X0_LVT div_U945 ( .A1(div_n291), .A2(div_n744), .A3(div_n_T_51_5_), .Y(
        div_n985) );
  OA22X1_LVT div_U944 ( .A1(div_n283), .A2(div_n_T_51_14_), .A3(div_n743), 
        .A4(div_n737), .Y(div_n986) );
  NAND2X0_LVT div_U943 ( .A1(div_n286), .A2(div_n_T_51_9_), .Y(div_n737) );
  INVX1_LVT div_U942 ( .A(div_n780), .Y(div_n743) );
  AND4X1_LVT div_U941 ( .A1(div_n281), .A2(div_n736), .A3(div_n735), .A4(
        div_n734), .Y(div_n757) );
  NAND2X0_LVT div_U940 ( .A1(div_n780), .A2(div_n_T_51_11_), .Y(div_n734) );
  NAND2X0_LVT div_U939 ( .A1(div_n305), .A2(div_n745), .Y(div_n735) );
  NAND2X0_LVT div_U938 ( .A1(div_n744), .A2(div_n_T_51_7_), .Y(div_n736) );
  NAND3X0_LVT div_U937 ( .A1(div_n241), .A2(div_n_T_51_49_), .A3(div_n747), 
        .Y(div_n981) );
  NAND3X0_LVT div_U936 ( .A1(div_n237), .A2(div_n773), .A3(div_n_T_51_53_), 
        .Y(div_n982) );
  OA22X1_LVT div_U935 ( .A1(div_n229), .A2(div_n_T_51_62_), .A3(div_n733), 
        .A4(div_n746), .Y(div_n983) );
  INVX1_LVT div_U934 ( .A(div_n774), .Y(div_n746) );
  NAND2X0_LVT div_U933 ( .A1(div_n232), .A2(div_n_T_51_57_), .Y(div_n733) );
  OR2X1_LVT div_U932 ( .A1(div_n971), .A2(div_n999), .Y(div_n998) );
  AND2X1_LVT div_U931 ( .A1(div_n747), .A2(div_n732), .Y(div_n1002) );
  AND2X1_LVT div_U930 ( .A1(div_n773), .A2(div_n779), .Y(div_n747) );
  NAND4X0_LVT div_U929 ( .A1(div_n174), .A2(div_n731), .A3(div_n730), .A4(
        div_n729), .Y(div_n951) );
  NAND2X0_LVT div_U928 ( .A1(div_n764), .A2(div_divisor_26_), .Y(div_n729) );
  NAND2X0_LVT div_U927 ( .A1(div_divisor_22_), .A2(div_n728), .Y(div_n730) );
  NAND2X0_LVT div_U926 ( .A1(div_n727), .A2(div_divisor_18_), .Y(div_n731) );
  NAND4X0_LVT div_U925 ( .A1(div_n762), .A2(div_n726), .A3(div_n725), .A4(
        div_n724), .Y(div_n952) );
  NAND2X0_LVT div_U924 ( .A1(div_n766), .A2(div_divisor_34_), .Y(div_n724) );
  NAND2X0_LVT div_U923 ( .A1(div_divisor_38_), .A2(div_n723), .Y(div_n725) );
  OA21X1_LVT div_U922 ( .A1(div_n185), .A2(div_n722), .A3(div_n194), .Y(
        div_n726) );
  NAND4X0_LVT div_U921 ( .A1(div_n177), .A2(div_n721), .A3(div_n720), .A4(
        div_n719), .Y(div_n948) );
  NAND2X0_LVT div_U920 ( .A1(div_n769), .A2(div_n718), .Y(div_n719) );
  INVX1_LVT div_U919 ( .A(div_n179), .Y(div_n718) );
  NAND2X0_LVT div_U918 ( .A1(div_n216), .A2(div_divisor_54_), .Y(div_n720) );
  NAND2X0_LVT div_U917 ( .A1(div_n717), .A2(div_divisor_50_), .Y(div_n721) );
  NAND3X0_LVT div_U916 ( .A1(div_n759), .A2(div_n193), .A3(div_n716), .Y(
        div_n949) );
  OR2X1_LVT div_U915 ( .A1(div_n202), .A2(div_n715), .Y(div_n716) );
  AO22X1_LVT div_U914 ( .A1(div_divisor_6_), .A2(div_n714), .A3(div_n713), 
        .A4(div_n712), .Y(div_n950) );
  INVX1_LVT div_U913 ( .A(div_n205), .Y(div_n712) );
  AO21X1_LVT div_U912 ( .A1(div_n763), .A2(div_n711), .A3(div_n710), .Y(
        div_n955) );
  NAND4X0_LVT div_U911 ( .A1(div_n175), .A2(div_n709), .A3(div_n708), .A4(
        div_n707), .Y(div_n710) );
  NAND2X0_LVT div_U910 ( .A1(div_n769), .A2(div_divisor_59_), .Y(div_n707) );
  NAND2X0_LVT div_U909 ( .A1(div_n216), .A2(div_divisor_55_), .Y(div_n708) );
  NAND2X0_LVT div_U908 ( .A1(div_divisor_51_), .A2(div_n717), .Y(div_n709) );
  NAND4X0_LVT div_U907 ( .A1(div_n176), .A2(div_n706), .A3(div_n705), .A4(
        div_n704), .Y(div_n711) );
  NAND2X0_LVT div_U906 ( .A1(div_n764), .A2(div_divisor_27_), .Y(div_n704) );
  NAND2X0_LVT div_U905 ( .A1(div_divisor_23_), .A2(div_n728), .Y(div_n705) );
  NAND2X0_LVT div_U904 ( .A1(div_n727), .A2(div_divisor_19_), .Y(div_n706) );
  NAND3X0_LVT div_U903 ( .A1(div_n713), .A2(div_n205), .A3(div_divisor_1_), 
        .Y(div_n941) );
  NAND3X0_LVT div_U902 ( .A1(div_divisor_5_), .A2(div_n714), .A3(div_n191), 
        .Y(div_n942) );
  OA22X1_LVT div_U901 ( .A1(div_divisor_14_), .A2(div_n172), .A3(div_n703), 
        .A4(div_n715), .Y(div_n943) );
  INVX1_LVT div_U900 ( .A(div_n761), .Y(div_n715) );
  NAND2X0_LVT div_U899 ( .A1(div_divisor_9_), .A2(div_n202), .Y(div_n703) );
  AND4X1_LVT div_U898 ( .A1(div_n162), .A2(div_n702), .A3(div_n701), .A4(
        div_n700), .Y(div_n759) );
  NAND2X0_LVT div_U897 ( .A1(div_n761), .A2(div_divisor_11_), .Y(div_n700) );
  NAND2X0_LVT div_U896 ( .A1(div_divisor_7_), .A2(div_n714), .Y(div_n701) );
  NAND2X0_LVT div_U895 ( .A1(div_n713), .A2(div_divisor_3_), .Y(div_n702) );
  AND2X1_LVT div_U894 ( .A1(div_n760), .A2(div_n714), .Y(div_n713) );
  INVX1_LVT div_U893 ( .A(div_n962), .Y(div_n714) );
  NOR4X1_LVT div_U892 ( .A1(div_divisor_6_), .A2(div_divisor_7_), .A3(
        div_divisor_5_), .A4(div_divisor_4_), .Y(div_n760) );
  NAND4X0_LVT div_U891 ( .A1(div_n699), .A2(div_n761), .A3(div_n202), .A4(
        div_n165), .Y(div_n962) );
  NOR4X1_LVT div_U890 ( .A1(div_divisor_14_), .A2(div_divisor_13_), .A3(
        div_divisor_15_), .A4(div_divisor_12_), .Y(div_n761) );
  NAND3X0_LVT div_U889 ( .A1(div_n766), .A2(div_divisor_33_), .A3(div_n160), 
        .Y(div_n937) );
  NAND3X0_LVT div_U888 ( .A1(div_divisor_37_), .A2(div_n723), .A3(div_n192), 
        .Y(div_n938) );
  OA22X1_LVT div_U887 ( .A1(div_divisor_46_), .A2(div_n173), .A3(div_n698), 
        .A4(div_n722), .Y(div_n939) );
  INVX1_LVT div_U886 ( .A(div_n767), .Y(div_n722) );
  NAND2X0_LVT div_U885 ( .A1(div_divisor_41_), .A2(div_n185), .Y(div_n698) );
  AND4X1_LVT div_U884 ( .A1(div_n178), .A2(div_n697), .A3(div_n696), .A4(
        div_n695), .Y(div_n762) );
  NAND2X0_LVT div_U883 ( .A1(div_n767), .A2(div_divisor_43_), .Y(div_n695) );
  NAND2X0_LVT div_U882 ( .A1(div_divisor_39_), .A2(div_n723), .Y(div_n696) );
  NAND2X0_LVT div_U881 ( .A1(div_n766), .A2(div_divisor_35_), .Y(div_n697) );
  NAND2X0_LVT div_U880 ( .A1(div_divisor_61_), .A2(div_n177), .Y(div_n933) );
  NAND3X0_LVT div_U879 ( .A1(div_n769), .A2(div_divisor_57_), .A3(div_n179), 
        .Y(div_n934) );
  NAND3X0_LVT div_U878 ( .A1(div_n216), .A2(div_divisor_53_), .A3(div_n195), 
        .Y(div_n935) );
  OA21X1_LVT div_U877 ( .A1(div_n694), .A2(div_n968), .A3(div_n693), .Y(
        div_n936) );
  NAND3X0_LVT div_U876 ( .A1(div_n717), .A2(div_divisor_49_), .A3(div_n159), 
        .Y(div_n693) );
  AND4X1_LVT div_U875 ( .A1(div_n692), .A2(div_n691), .A3(div_n690), .A4(
        div_n689), .Y(div_n694) );
  NAND2X0_LVT div_U874 ( .A1(div_divisor_29_), .A2(div_n174), .Y(div_n689) );
  NAND3X0_LVT div_U873 ( .A1(div_n764), .A2(div_divisor_25_), .A3(div_n196), 
        .Y(div_n690) );
  NAND3X0_LVT div_U872 ( .A1(div_divisor_21_), .A2(div_n728), .A3(div_n190), 
        .Y(div_n691) );
  NAND3X0_LVT div_U871 ( .A1(div_n727), .A2(div_divisor_17_), .A3(div_n161), 
        .Y(div_n692) );
  AND2X1_LVT div_U870 ( .A1(div_n727), .A2(div_n688), .Y(div_n940) );
  NOR4X1_LVT div_U869 ( .A1(div_divisor_18_), .A2(div_divisor_19_), .A3(
        div_divisor_17_), .A4(div_divisor_16_), .Y(div_n688) );
  AND2X1_LVT div_U868 ( .A1(div_n765), .A2(div_n728), .Y(div_n727) );
  INVX1_LVT div_U867 ( .A(div_n964), .Y(div_n728) );
  NOR4X1_LVT div_U866 ( .A1(div_divisor_22_), .A2(div_divisor_20_), .A3(
        div_divisor_23_), .A4(div_divisor_21_), .Y(div_n765) );
  NAND4X0_LVT div_U865 ( .A1(div_n687), .A2(div_n764), .A3(div_n196), .A4(
        div_n164), .Y(div_n964) );
  NOR4X1_LVT div_U864 ( .A1(div_divisor_31_), .A2(div_divisor_30_), .A3(
        div_divisor_29_), .A4(div_divisor_28_), .Y(div_n764) );
  NOR4X1_LVT div_U863 ( .A1(div_divisor_35_), .A2(div_divisor_34_), .A3(
        div_divisor_33_), .A4(div_divisor_32_), .Y(div_n932) );
  AND2X1_LVT div_U862 ( .A1(div_n768), .A2(div_n723), .Y(div_n766) );
  NOR4X1_LVT div_U861 ( .A1(div_divisor_38_), .A2(div_divisor_37_), .A3(
        div_divisor_39_), .A4(div_divisor_36_), .Y(div_n768) );
  NAND4X0_LVT div_U860 ( .A1(div_n686), .A2(div_n767), .A3(div_n185), .A4(
        div_n163), .Y(div_n966) );
  NOR4X1_LVT div_U859 ( .A1(div_divisor_46_), .A2(div_divisor_45_), .A3(
        div_divisor_47_), .A4(div_divisor_44_), .Y(div_n767) );
  NAND2X0_LVT div_U858 ( .A1(div_n717), .A2(div_n685), .Y(div_n956) );
  NOR4X1_LVT div_U857 ( .A1(div_divisor_51_), .A2(div_divisor_50_), .A3(
        div_divisor_49_), .A4(div_divisor_48_), .Y(div_n685) );
  AND2X1_LVT div_U856 ( .A1(div_n216), .A2(div_n770), .Y(div_n717) );
  NOR4X1_LVT div_U855 ( .A1(div_divisor_55_), .A2(div_divisor_54_), .A3(
        div_divisor_53_), .A4(div_divisor_52_), .Y(div_n770) );
  NAND4X0_LVT div_U854 ( .A1(div_n684), .A2(div_n769), .A3(div_n179), .A4(
        div_n180), .Y(div_n967) );
  NOR4X1_LVT div_U853 ( .A1(div_divisor_62_), .A2(div_divisor_61_), .A3(
        div_divisor_63_), .A4(div_divisor_60_), .Y(div_n769) );
  NOR2X0_LVT div_U852 ( .A1(div_divisor_57_), .A2(div_divisor_56_), .Y(
        div_n684) );
  NAND4X0_LVT div_U851 ( .A1(div_n254), .A2(div_n257), .A3(div_n256), .A4(
        div_n255), .Y(div_n971) );
  NAND2X0_LVT div_U850 ( .A1(div_n772), .A2(div_n771), .Y(div_n999) );
  AND4X1_LVT div_U849 ( .A1(div_n248), .A2(div_n246), .A3(div_n249), .A4(
        div_n247), .Y(div_n771) );
  AND4X1_LVT div_U848 ( .A1(div_n188), .A2(div_n251), .A3(div_n250), .A4(
        div_n252), .Y(div_n772) );
  NAND4X0_LVT div_U847 ( .A1(div_n259), .A2(div_n258), .A3(div_n261), .A4(
        div_n260), .Y(div_n970) );
  AND4X1_LVT div_U846 ( .A1(div_n231), .A2(div_n234), .A3(div_n233), .A4(
        div_n232), .Y(div_n683) );
  AND4X1_LVT div_U845 ( .A1(div_n187), .A2(div_n149), .A3(div_n228), .A4(
        div_n229), .Y(div_n774) );
  AND2X1_LVT div_U844 ( .A1(div_n776), .A2(div_n682), .Y(div_n775) );
  AND4X1_LVT div_U843 ( .A1(div_n267), .A2(div_n270), .A3(div_n269), .A4(
        div_n268), .Y(div_n682) );
  AND4X1_LVT div_U842 ( .A1(div_n181), .A2(div_n264), .A3(div_n263), .A4(
        div_n266), .Y(div_n776) );
  NAND4X0_LVT div_U841 ( .A1(div_n277), .A2(div_n278), .A3(div_n152), .A4(
        div_n183), .Y(div_n973) );
  AND4X1_LVT div_U840 ( .A1(div_n272), .A2(div_n275), .A3(div_n274), .A4(
        div_n273), .Y(div_n777) );
  AO22X1_LVT div_U839 ( .A1(div_n157), .A2(div_n171), .A3(div_n805), .A4(
        div_n204), .Y(div_N294) );
  AO222X1_LVT div_U838 ( .A1(div_n783), .A2(div_n_T_65[71]), .A3(div_n931), 
        .A4(div_n_T_51_126_), .A5(div_subtractor_63_), .A6(div_n226), .Y(
        div_N523) );
  AO21X1_LVT div_U837 ( .A1(div_n753), .A2(div_n681), .A3(div_n680), .Y(
        div_N285) );
  OR2X1_LVT div_U836 ( .A1(div_n977), .A2(div_n978), .Y(div_n681) );
  AND2X1_LVT div_U835 ( .A1(div_n224), .A2(div_n154), .Y(div_n977) );
  NAND4X0_LVT div_U834 ( .A1(div_n678), .A2(div_n677), .A3(div_n676), .A4(
        div_n675), .Y(div_N403) );
  NAND2X0_LVT div_U833 ( .A1(div_negated_remainder[9]), .A2(div_n224), .Y(
        div_n675) );
  NAND2X0_LVT div_U832 ( .A1(div_n227), .A2(div_n_T_51_8_), .Y(div_n676) );
  AOI21X1_LVT div_U831 ( .A1(div_n679), .A2(div_n_T_87[9]), .A3(div_n674), .Y(
        div_n677) );
  AO22X1_LVT div_U830 ( .A1(div_n235), .A2(io_fpu_fromint_data[9]), .A3(
        div_n223), .A4(div_n_T_51_17_), .Y(div_n674) );
  NAND2X0_LVT div_U829 ( .A1(div_n157), .A2(div_n_T_442[9]), .Y(div_n678) );
  NAND4X0_LVT div_U828 ( .A1(div_n673), .A2(div_n672), .A3(div_n671), .A4(
        div_n670), .Y(div_N411) );
  NAND2X0_LVT div_U827 ( .A1(div_negated_remainder[17]), .A2(div_n224), .Y(
        div_n670) );
  NAND2X0_LVT div_U826 ( .A1(div_n227), .A2(div_n_T_51_16_), .Y(div_n671) );
  AOI21X1_LVT div_U825 ( .A1(div_n679), .A2(div_n_T_87[17]), .A3(div_n669), 
        .Y(div_n672) );
  AO22X1_LVT div_U824 ( .A1(div_n235), .A2(io_fpu_fromint_data[17]), .A3(
        div_n223), .A4(div_n_T_51_25_), .Y(div_n669) );
  NAND2X0_LVT div_U823 ( .A1(div_n225), .A2(div_n_T_442[17]), .Y(div_n673) );
  NAND4X0_LVT div_U822 ( .A1(div_n668), .A2(div_n667), .A3(div_n666), .A4(
        div_n665), .Y(div_N419) );
  NAND2X0_LVT div_U821 ( .A1(div_negated_remainder[25]), .A2(div_n224), .Y(
        div_n665) );
  NAND2X0_LVT div_U820 ( .A1(div_n227), .A2(div_n_T_51_24_), .Y(div_n666) );
  AOI21X1_LVT div_U819 ( .A1(div_n679), .A2(div_n_T_87[25]), .A3(div_n664), 
        .Y(div_n667) );
  AO22X1_LVT div_U818 ( .A1(div_n235), .A2(io_fpu_fromint_data[25]), .A3(
        div_n223), .A4(div_n_T_51_33_), .Y(div_n664) );
  NAND2X0_LVT div_U817 ( .A1(div_n225), .A2(div_n_T_442[25]), .Y(div_n668) );
  NAND4X0_LVT div_U816 ( .A1(div_n663), .A2(div_n662), .A3(div_n661), .A4(
        div_n660), .Y(div_N427) );
  NAND2X0_LVT div_U815 ( .A1(div_negated_remainder[33]), .A2(div_n224), .Y(
        div_n660) );
  NAND2X0_LVT div_U814 ( .A1(div_n227), .A2(div_n_T_51_32_), .Y(div_n661) );
  AND4X1_LVT div_U813 ( .A1(div_n659), .A2(div_n658), .A3(div_n657), .A4(
        div_n656), .Y(div_n662) );
  NAND2X0_LVT div_U812 ( .A1(div_n655), .A2(io_fpu_fromint_data[33]), .Y(
        div_n656) );
  NAND2X0_LVT div_U811 ( .A1(div_n223), .A2(div_n_T_51_41_), .Y(div_n657) );
  NAND2X0_LVT div_U810 ( .A1(div_n_T_87[33]), .A2(div_n679), .Y(div_n659) );
  NAND2X0_LVT div_U809 ( .A1(div_n_T_442[33]), .A2(div_n225), .Y(div_n663) );
  NAND4X0_LVT div_U808 ( .A1(div_n654), .A2(div_n653), .A3(div_n652), .A4(
        div_n651), .Y(div_N435) );
  NAND2X0_LVT div_U807 ( .A1(div_negated_remainder[41]), .A2(div_n224), .Y(
        div_n651) );
  NAND2X0_LVT div_U806 ( .A1(div_n227), .A2(div_n_T_51_40_), .Y(div_n652) );
  AND4X1_LVT div_U805 ( .A1(div_n650), .A2(div_n658), .A3(div_n649), .A4(
        div_n648), .Y(div_n653) );
  NAND2X0_LVT div_U804 ( .A1(div_n655), .A2(io_fpu_fromint_data[41]), .Y(
        div_n648) );
  NAND2X0_LVT div_U803 ( .A1(div_n223), .A2(div_n_T_51_49_), .Y(div_n649) );
  NAND2X0_LVT div_U802 ( .A1(div_n_T_87[41]), .A2(div_n679), .Y(div_n650) );
  NAND2X0_LVT div_U801 ( .A1(div_n_T_442[41]), .A2(div_n157), .Y(div_n654) );
  NAND4X0_LVT div_U800 ( .A1(div_n647), .A2(div_n646), .A3(div_n645), .A4(
        div_n644), .Y(div_N443) );
  NAND2X0_LVT div_U799 ( .A1(div_negated_remainder[49]), .A2(div_n224), .Y(
        div_n644) );
  NAND2X0_LVT div_U798 ( .A1(div_n227), .A2(div_n_T_51_48_), .Y(div_n645) );
  AND4X1_LVT div_U797 ( .A1(div_n643), .A2(div_n658), .A3(div_n642), .A4(
        div_n641), .Y(div_n646) );
  NAND2X0_LVT div_U796 ( .A1(div_n655), .A2(io_fpu_fromint_data[49]), .Y(
        div_n641) );
  NAND2X0_LVT div_U795 ( .A1(div_n223), .A2(div_n_T_51_57_), .Y(div_n642) );
  NAND2X0_LVT div_U794 ( .A1(div_n_T_87[49]), .A2(div_n679), .Y(div_n643) );
  NAND2X0_LVT div_U793 ( .A1(div_n_T_442[49]), .A2(div_n157), .Y(div_n647) );
  NAND4X0_LVT div_U792 ( .A1(div_n640), .A2(div_n639), .A3(div_n638), .A4(
        div_n637), .Y(div_N451) );
  NAND2X0_LVT div_U791 ( .A1(div_n227), .A2(div_n_T_51_56_), .Y(div_n637) );
  NAND2X0_LVT div_U790 ( .A1(div_n_T_442[57]), .A2(div_n225), .Y(div_n638) );
  AND4X1_LVT div_U789 ( .A1(div_n636), .A2(div_n658), .A3(div_n635), .A4(
        div_n634), .Y(div_n639) );
  NAND2X0_LVT div_U788 ( .A1(div_n655), .A2(io_fpu_fromint_data[57]), .Y(
        div_n634) );
  NAND2X0_LVT div_U787 ( .A1(div_n223), .A2(div_n_T_65[1]), .Y(div_n635) );
  NAND2X0_LVT div_U786 ( .A1(div_n_T_87[57]), .A2(div_n679), .Y(div_n636) );
  NAND2X0_LVT div_U785 ( .A1(div_negated_remainder[57]), .A2(div_n224), .Y(
        div_n640) );
  AO22X1_LVT div_U784 ( .A1(div_n754), .A2(div_subtractor_0_), .A3(n_T_702[0]), 
        .A4(div_n235), .Y(div_N323) );
  AO22X1_LVT div_U783 ( .A1(div_n754), .A2(div_subtractor_1_), .A3(n_T_702[1]), 
        .A4(div_n235), .Y(div_N324) );
  AO22X1_LVT div_U782 ( .A1(n_T_702[2]), .A2(div_n235), .A3(div_subtractor_2_), 
        .A4(div_n754), .Y(div_N325) );
  AO22X1_LVT div_U781 ( .A1(div_n235), .A2(n_T_702[3]), .A3(div_subtractor_3_), 
        .A4(div_n754), .Y(div_N326) );
  AO22X1_LVT div_U780 ( .A1(div_n235), .A2(n_T_702[4]), .A3(div_subtractor_4_), 
        .A4(div_n754), .Y(div_N327) );
  AO22X1_LVT div_U779 ( .A1(div_n235), .A2(n_T_702[5]), .A3(div_subtractor_5_), 
        .A4(div_n754), .Y(div_N328) );
  AO22X1_LVT div_U778 ( .A1(div_n235), .A2(n_T_702[6]), .A3(div_subtractor_6_), 
        .A4(div_n754), .Y(div_N329) );
  AO22X1_LVT div_U777 ( .A1(div_n235), .A2(n_T_702[7]), .A3(div_subtractor_7_), 
        .A4(div_n754), .Y(div_N330) );
  AO22X1_LVT div_U776 ( .A1(div_n235), .A2(n_T_702[8]), .A3(div_subtractor_8_), 
        .A4(div_n754), .Y(div_N331) );
  AO22X1_LVT div_U775 ( .A1(div_n235), .A2(n_T_702[9]), .A3(div_subtractor_9_), 
        .A4(div_n754), .Y(div_N332) );
  AO22X1_LVT div_U774 ( .A1(div_n235), .A2(n_T_702[10]), .A3(
        div_subtractor_10_), .A4(div_n754), .Y(div_N333) );
  AO22X1_LVT div_U773 ( .A1(div_n235), .A2(n_T_702[11]), .A3(
        div_subtractor_11_), .A4(div_n754), .Y(div_N334) );
  AO22X1_LVT div_U772 ( .A1(div_n235), .A2(n_T_702[12]), .A3(
        div_subtractor_12_), .A4(div_n754), .Y(div_N335) );
  AO22X1_LVT div_U771 ( .A1(div_n235), .A2(n_T_702[13]), .A3(
        div_subtractor_13_), .A4(div_n754), .Y(div_N336) );
  AO22X1_LVT div_U770 ( .A1(div_n235), .A2(n_T_702[14]), .A3(
        div_subtractor_14_), .A4(div_n754), .Y(div_N337) );
  AO22X1_LVT div_U769 ( .A1(div_n235), .A2(n_T_702[15]), .A3(
        div_subtractor_15_), .A4(div_n754), .Y(div_N338) );
  AO22X1_LVT div_U768 ( .A1(div_n235), .A2(n_T_702[16]), .A3(
        div_subtractor_16_), .A4(div_n754), .Y(div_N339) );
  AO22X1_LVT div_U767 ( .A1(div_n235), .A2(n_T_702[17]), .A3(
        div_subtractor_17_), .A4(div_n754), .Y(div_N340) );
  AO22X1_LVT div_U766 ( .A1(div_n235), .A2(n_T_702[18]), .A3(
        div_subtractor_18_), .A4(div_n754), .Y(div_N341) );
  AO22X1_LVT div_U765 ( .A1(div_n235), .A2(n_T_702[19]), .A3(
        div_subtractor_19_), .A4(div_n754), .Y(div_N342) );
  AO22X1_LVT div_U764 ( .A1(div_n235), .A2(n_T_702[20]), .A3(
        div_subtractor_20_), .A4(div_n754), .Y(div_N343) );
  AO22X1_LVT div_U763 ( .A1(div_n235), .A2(n_T_702[21]), .A3(
        div_subtractor_21_), .A4(div_n754), .Y(div_N344) );
  AO22X1_LVT div_U762 ( .A1(div_n235), .A2(n_T_702[22]), .A3(
        div_subtractor_22_), .A4(div_n754), .Y(div_N345) );
  AO22X1_LVT div_U761 ( .A1(div_n235), .A2(n_T_702[23]), .A3(
        div_subtractor_23_), .A4(div_n754), .Y(div_N346) );
  AO22X1_LVT div_U760 ( .A1(div_n235), .A2(n_T_702[24]), .A3(
        div_subtractor_24_), .A4(div_n754), .Y(div_N347) );
  AO22X1_LVT div_U759 ( .A1(div_n235), .A2(n_T_702[25]), .A3(
        div_subtractor_25_), .A4(div_n754), .Y(div_N348) );
  AO22X1_LVT div_U758 ( .A1(div_n235), .A2(n_T_702[26]), .A3(
        div_subtractor_26_), .A4(div_n754), .Y(div_N349) );
  AO22X1_LVT div_U757 ( .A1(div_n235), .A2(n_T_702[27]), .A3(
        div_subtractor_27_), .A4(div_n754), .Y(div_N350) );
  AO22X1_LVT div_U756 ( .A1(div_n235), .A2(n_T_702[28]), .A3(
        div_subtractor_28_), .A4(div_n754), .Y(div_N351) );
  AO22X1_LVT div_U755 ( .A1(div_n235), .A2(n_T_702[29]), .A3(
        div_subtractor_29_), .A4(div_n754), .Y(div_N352) );
  AO22X1_LVT div_U754 ( .A1(div_n235), .A2(n_T_702[30]), .A3(
        div_subtractor_30_), .A4(div_n754), .Y(div_N353) );
  AO22X1_LVT div_U753 ( .A1(div_n235), .A2(n_T_702[31]), .A3(
        div_subtractor_31_), .A4(div_n754), .Y(div_N354) );
  NAND3X0_LVT div_U752 ( .A1(div_n632), .A2(div_n633), .A3(div_n631), .Y(
        div_N356) );
  NAND2X0_LVT div_U751 ( .A1(n_T_702[33]), .A2(div_n655), .Y(div_n631) );
  NAND2X0_LVT div_U750 ( .A1(div_subtractor_33_), .A2(div_n754), .Y(div_n632)
         );
  NAND3X0_LVT div_U749 ( .A1(div_n630), .A2(div_n633), .A3(div_n629), .Y(
        div_N357) );
  NAND2X0_LVT div_U748 ( .A1(n_T_702[34]), .A2(div_n655), .Y(div_n629) );
  NAND2X0_LVT div_U747 ( .A1(div_subtractor_34_), .A2(div_n754), .Y(div_n630)
         );
  NAND3X0_LVT div_U746 ( .A1(div_n628), .A2(div_n633), .A3(div_n627), .Y(
        div_N359) );
  NAND2X0_LVT div_U745 ( .A1(n_T_702[36]), .A2(div_n655), .Y(div_n627) );
  NAND2X0_LVT div_U744 ( .A1(div_subtractor_36_), .A2(div_n754), .Y(div_n628)
         );
  NAND3X0_LVT div_U743 ( .A1(div_n626), .A2(div_n633), .A3(div_n625), .Y(
        div_N360) );
  NAND2X0_LVT div_U742 ( .A1(n_T_702[37]), .A2(div_n655), .Y(div_n625) );
  NAND2X0_LVT div_U741 ( .A1(div_subtractor_37_), .A2(div_n754), .Y(div_n626)
         );
  NAND3X0_LVT div_U740 ( .A1(div_n624), .A2(div_n633), .A3(div_n623), .Y(
        div_N361) );
  NAND2X0_LVT div_U739 ( .A1(n_T_702[38]), .A2(div_n655), .Y(div_n623) );
  NAND2X0_LVT div_U738 ( .A1(div_subtractor_38_), .A2(div_n754), .Y(div_n624)
         );
  NAND3X0_LVT div_U737 ( .A1(div_n622), .A2(div_n633), .A3(div_n621), .Y(
        div_N362) );
  NAND2X0_LVT div_U736 ( .A1(n_T_702[39]), .A2(div_n655), .Y(div_n621) );
  NAND2X0_LVT div_U735 ( .A1(div_subtractor_39_), .A2(div_n754), .Y(div_n622)
         );
  NAND3X0_LVT div_U734 ( .A1(div_n620), .A2(div_n633), .A3(div_n619), .Y(
        div_N365) );
  NAND2X0_LVT div_U733 ( .A1(n_T_702[42]), .A2(div_n655), .Y(div_n619) );
  NAND2X0_LVT div_U732 ( .A1(div_subtractor_42_), .A2(div_n754), .Y(div_n620)
         );
  NAND3X0_LVT div_U731 ( .A1(div_n618), .A2(div_n633), .A3(div_n617), .Y(
        div_N368) );
  NAND2X0_LVT div_U730 ( .A1(n_T_702[45]), .A2(div_n655), .Y(div_n617) );
  NAND2X0_LVT div_U729 ( .A1(div_subtractor_45_), .A2(div_n754), .Y(div_n618)
         );
  AO22X1_LVT div_U728 ( .A1(div_n235), .A2(div_n616), .A3(div_subtractor_64_), 
        .A4(div_n754), .Y(div_N387) );
  NAND4X0_LVT div_U727 ( .A1(div_n612), .A2(div_n611), .A3(div_n610), .A4(
        div_n609), .Y(div_N457) );
  NAND2X0_LVT div_U726 ( .A1(div_n_T_442[63]), .A2(div_n225), .Y(div_n609) );
  NAND2X0_LVT div_U725 ( .A1(div_n227), .A2(div_n_T_51_62_), .Y(div_n610) );
  AND4X1_LVT div_U724 ( .A1(div_n608), .A2(div_n607), .A3(div_n606), .A4(
        div_n658), .Y(div_n611) );
  NAND2X0_LVT div_U723 ( .A1(div_n655), .A2(io_fpu_fromint_data[63]), .Y(
        div_n606) );
  NAND2X0_LVT div_U722 ( .A1(div_n_T_87[63]), .A2(div_n679), .Y(div_n607) );
  NAND2X0_LVT div_U721 ( .A1(div_n_T_65[7]), .A2(div_n223), .Y(div_n608) );
  NAND2X0_LVT div_U720 ( .A1(div_negated_remainder[63]), .A2(div_n224), .Y(
        div_n612) );
  OA21X1_LVT div_U719 ( .A1(div_n300), .A2(div_n_T_69_4_), .A3(div_n_T_71_39_), 
        .Y(div_n788) );
  AO21X1_LVT div_U718 ( .A1(div_negated_remainder[62]), .A2(div_n224), .A3(
        div_n604), .Y(div_N456) );
  AO21X1_LVT div_U717 ( .A1(div_n225), .A2(div_n_T_442[62]), .A3(div_n603), 
        .Y(div_n604) );
  AO21X1_LVT div_U716 ( .A1(div_n227), .A2(div_n_T_51_61_), .A3(div_n602), .Y(
        div_n603) );
  NAND4X0_LVT div_U715 ( .A1(div_n601), .A2(div_n658), .A3(div_n600), .A4(
        div_n599), .Y(div_n602) );
  NAND2X0_LVT div_U714 ( .A1(div_n655), .A2(io_fpu_fromint_data[62]), .Y(
        div_n599) );
  NAND2X0_LVT div_U713 ( .A1(div_n_T_87[62]), .A2(div_n679), .Y(div_n600) );
  NAND2X0_LVT div_U712 ( .A1(div_n_T_65[6]), .A2(div_n223), .Y(div_n601) );
  MUX21X1_LVT div_U711 ( .A1(div_n302), .A2(div_n_T_51_64_), .S0(div_n308), 
        .Y(div_result_0_) );
  MUX21X1_LVT div_U710 ( .A1(div_n_T_51_1_), .A2(div_n_T_51_65_), .S0(div_n308), .Y(div_result_1_) );
  MUX21X1_LVT div_U709 ( .A1(div_n304), .A2(div_n_T_51_66_), .S0(div_n308), 
        .Y(div_result_2_) );
  MUX21X1_LVT div_U708 ( .A1(div_n305), .A2(div_n_T_51_67_), .S0(div_n308), 
        .Y(div_result_3_) );
  MUX21X1_LVT div_U707 ( .A1(div_n_T_51_4_), .A2(div_n_T_51_68_), .S0(div_n308), .Y(div_result_4_) );
  MUX21X1_LVT div_U706 ( .A1(div_n_T_51_5_), .A2(div_n_T_51_69_), .S0(div_n308), .Y(div_result_5_) );
  MUX21X1_LVT div_U705 ( .A1(div_n_T_51_6_), .A2(div_n_T_51_70_), .S0(
        div_resHi), .Y(div_result_6_) );
  MUX21X1_LVT div_U704 ( .A1(div_n_T_51_7_), .A2(div_n_T_51_71_), .S0(div_n308), .Y(div_result_7_) );
  MUX21X1_LVT div_U703 ( .A1(div_n_T_51_8_), .A2(div_n_T_51_72_), .S0(
        div_resHi), .Y(div_result_8_) );
  NAND4X0_LVT div_U702 ( .A1(div_n598), .A2(div_n597), .A3(div_n596), .A4(
        div_n595), .Y(div_N402) );
  NAND2X0_LVT div_U701 ( .A1(div_negated_remainder[8]), .A2(div_n224), .Y(
        div_n595) );
  NAND2X0_LVT div_U700 ( .A1(div_n227), .A2(div_n_T_51_7_), .Y(div_n596) );
  AOI21X1_LVT div_U699 ( .A1(div_n679), .A2(div_n_T_87[8]), .A3(div_n594), .Y(
        div_n597) );
  AO22X1_LVT div_U698 ( .A1(div_n235), .A2(io_fpu_fromint_data[8]), .A3(
        div_n223), .A4(div_n_T_51_16_), .Y(div_n594) );
  NAND2X0_LVT div_U697 ( .A1(div_n225), .A2(div_n_T_442[8]), .Y(div_n598) );
  NAND4X0_LVT div_U696 ( .A1(div_n593), .A2(div_n592), .A3(div_n591), .A4(
        div_n590), .Y(div_N401) );
  NAND2X0_LVT div_U695 ( .A1(div_negated_remainder[7]), .A2(div_n224), .Y(
        div_n590) );
  NAND2X0_LVT div_U694 ( .A1(div_n227), .A2(div_n_T_51_6_), .Y(div_n591) );
  AOI21X1_LVT div_U693 ( .A1(div_n679), .A2(div_n_T_87[7]), .A3(div_n589), .Y(
        div_n592) );
  AO22X1_LVT div_U692 ( .A1(io_fpu_fromint_data[7]), .A2(div_n235), .A3(
        div_n223), .A4(div_n_T_51_15_), .Y(div_n589) );
  NAND2X0_LVT div_U691 ( .A1(div_n157), .A2(div_n_T_442[7]), .Y(div_n593) );
  NAND4X0_LVT div_U690 ( .A1(div_n588), .A2(div_n587), .A3(div_n586), .A4(
        div_n585), .Y(div_N400) );
  NAND2X0_LVT div_U689 ( .A1(div_negated_remainder[6]), .A2(div_n224), .Y(
        div_n585) );
  NAND2X0_LVT div_U688 ( .A1(div_n227), .A2(div_n_T_51_5_), .Y(div_n586) );
  AOI21X1_LVT div_U687 ( .A1(div_n679), .A2(div_n_T_87[6]), .A3(div_n584), .Y(
        div_n587) );
  AO22X1_LVT div_U686 ( .A1(io_fpu_fromint_data[6]), .A2(div_n235), .A3(
        div_n223), .A4(div_n_T_51_14_), .Y(div_n584) );
  NAND2X0_LVT div_U685 ( .A1(div_n225), .A2(div_n_T_442[6]), .Y(div_n588) );
  NAND4X0_LVT div_U684 ( .A1(div_n583), .A2(div_n582), .A3(div_n581), .A4(
        div_n580), .Y(div_N399) );
  NAND2X0_LVT div_U683 ( .A1(div_negated_remainder[5]), .A2(div_n224), .Y(
        div_n580) );
  NAND2X0_LVT div_U682 ( .A1(div_n227), .A2(div_n_T_51_4_), .Y(div_n581) );
  AOI21X1_LVT div_U681 ( .A1(div_n679), .A2(div_n_T_87[5]), .A3(div_n579), .Y(
        div_n582) );
  AO22X1_LVT div_U680 ( .A1(io_fpu_fromint_data[5]), .A2(div_n235), .A3(
        div_n223), .A4(div_n_T_51_13_), .Y(div_n579) );
  NAND2X0_LVT div_U679 ( .A1(div_n225), .A2(div_n_T_442[5]), .Y(div_n583) );
  NAND4X0_LVT div_U678 ( .A1(div_n578), .A2(div_n577), .A3(div_n576), .A4(
        div_n575), .Y(div_N397) );
  NAND2X0_LVT div_U677 ( .A1(div_n_T_87[3]), .A2(div_n679), .Y(div_n575) );
  NAND2X0_LVT div_U676 ( .A1(div_n227), .A2(div_n304), .Y(div_n576) );
  AOI21X1_LVT div_U675 ( .A1(div_n_T_51_11_), .A2(div_n223), .A3(div_n574), 
        .Y(div_n577) );
  AO22X1_LVT div_U674 ( .A1(div_n235), .A2(io_fpu_fromint_data[3]), .A3(
        div_negated_remainder[3]), .A4(div_n224), .Y(div_n574) );
  NAND2X0_LVT div_U673 ( .A1(div_n225), .A2(div_n_T_442[3]), .Y(div_n578) );
  MUX21X1_LVT div_U672 ( .A1(div_n_T_51_9_), .A2(div_n_T_51_73_), .S0(div_n308), .Y(div_result_9_) );
  MUX21X1_LVT div_U671 ( .A1(div_n_T_51_10_), .A2(div_n_T_51_74_), .S0(
        div_resHi), .Y(div_result_10_) );
  MUX21X1_LVT div_U670 ( .A1(div_n_T_51_11_), .A2(div_n_T_51_75_), .S0(
        div_resHi), .Y(div_result_11_) );
  MUX21X1_LVT div_U669 ( .A1(div_n_T_51_12_), .A2(div_n_T_51_76_), .S0(
        div_n308), .Y(div_result_12_) );
  MUX21X1_LVT div_U668 ( .A1(div_n_T_51_13_), .A2(div_n_T_51_77_), .S0(
        div_n308), .Y(div_result_13_) );
  MUX21X1_LVT div_U667 ( .A1(div_n_T_51_15_), .A2(div_n_T_51_79_), .S0(
        div_n308), .Y(div_result_15_) );
  NAND4X0_LVT div_U666 ( .A1(div_n573), .A2(div_n572), .A3(div_n571), .A4(
        div_n570), .Y(div_N409) );
  NAND2X0_LVT div_U665 ( .A1(div_negated_remainder[15]), .A2(div_n224), .Y(
        div_n570) );
  NAND2X0_LVT div_U664 ( .A1(div_n227), .A2(div_n_T_51_14_), .Y(div_n571) );
  AOI21X1_LVT div_U663 ( .A1(div_n679), .A2(div_n_T_87[15]), .A3(div_n569), 
        .Y(div_n572) );
  AO22X1_LVT div_U662 ( .A1(div_n235), .A2(io_fpu_fromint_data[15]), .A3(
        div_n223), .A4(div_n_T_51_23_), .Y(div_n569) );
  NAND2X0_LVT div_U661 ( .A1(div_n157), .A2(div_n_T_442[15]), .Y(div_n573) );
  NAND4X0_LVT div_U660 ( .A1(div_n568), .A2(div_n567), .A3(div_n566), .A4(
        div_n565), .Y(div_N408) );
  NAND2X0_LVT div_U659 ( .A1(div_negated_remainder[14]), .A2(div_n224), .Y(
        div_n565) );
  NAND2X0_LVT div_U658 ( .A1(div_n227), .A2(div_n_T_51_13_), .Y(div_n566) );
  AOI21X1_LVT div_U657 ( .A1(div_n679), .A2(div_n_T_87[14]), .A3(div_n564), 
        .Y(div_n567) );
  AO22X1_LVT div_U656 ( .A1(div_n235), .A2(io_fpu_fromint_data[14]), .A3(
        div_n223), .A4(div_n_T_51_22_), .Y(div_n564) );
  NAND2X0_LVT div_U655 ( .A1(div_n225), .A2(div_n_T_442[14]), .Y(div_n568) );
  NAND4X0_LVT div_U654 ( .A1(div_n563), .A2(div_n562), .A3(div_n561), .A4(
        div_n560), .Y(div_N407) );
  NAND2X0_LVT div_U653 ( .A1(div_negated_remainder[13]), .A2(div_n224), .Y(
        div_n560) );
  NAND2X0_LVT div_U652 ( .A1(div_n227), .A2(div_n_T_51_12_), .Y(div_n561) );
  AOI21X1_LVT div_U651 ( .A1(div_n679), .A2(div_n_T_87[13]), .A3(div_n559), 
        .Y(div_n562) );
  AO22X1_LVT div_U650 ( .A1(div_n235), .A2(io_fpu_fromint_data[13]), .A3(
        div_n223), .A4(div_n_T_51_21_), .Y(div_n559) );
  NAND2X0_LVT div_U649 ( .A1(div_n225), .A2(div_n_T_442[13]), .Y(div_n563) );
  NAND4X0_LVT div_U648 ( .A1(div_n558), .A2(div_n557), .A3(div_n556), .A4(
        div_n555), .Y(div_N405) );
  NAND2X0_LVT div_U647 ( .A1(div_negated_remainder[11]), .A2(div_n224), .Y(
        div_n555) );
  NAND2X0_LVT div_U646 ( .A1(div_n227), .A2(div_n_T_51_10_), .Y(div_n556) );
  AOI21X1_LVT div_U645 ( .A1(div_n679), .A2(div_n_T_87[11]), .A3(div_n554), 
        .Y(div_n557) );
  AO22X1_LVT div_U644 ( .A1(div_n235), .A2(io_fpu_fromint_data[11]), .A3(
        div_n223), .A4(div_n_T_51_19_), .Y(div_n554) );
  NAND2X0_LVT div_U643 ( .A1(div_n225), .A2(div_n_T_442[11]), .Y(div_n558) );
  NAND4X0_LVT div_U642 ( .A1(div_n553), .A2(div_n552), .A3(div_n551), .A4(
        div_n550), .Y(div_N404) );
  NAND2X0_LVT div_U641 ( .A1(div_negated_remainder[10]), .A2(div_n224), .Y(
        div_n550) );
  NAND2X0_LVT div_U640 ( .A1(div_n227), .A2(div_n_T_51_9_), .Y(div_n551) );
  AOI21X1_LVT div_U639 ( .A1(div_n679), .A2(div_n_T_87[10]), .A3(div_n549), 
        .Y(div_n552) );
  AO22X1_LVT div_U638 ( .A1(div_n235), .A2(io_fpu_fromint_data[10]), .A3(
        div_n223), .A4(div_n_T_51_18_), .Y(div_n549) );
  NAND2X0_LVT div_U637 ( .A1(div_n225), .A2(div_n_T_442[10]), .Y(div_n553) );
  MUX21X1_LVT div_U636 ( .A1(div_n_T_51_17_), .A2(div_n_T_51_81_), .S0(
        div_n308), .Y(div_result_17_) );
  MUX21X1_LVT div_U635 ( .A1(div_n_T_51_18_), .A2(div_n_T_51_82_), .S0(
        div_n308), .Y(div_result_18_) );
  MUX21X1_LVT div_U634 ( .A1(div_n_T_51_19_), .A2(div_n_T_51_83_), .S0(
        div_n308), .Y(div_result_19_) );
  MUX21X1_LVT div_U633 ( .A1(div_n_T_51_20_), .A2(div_n_T_51_84_), .S0(
        div_resHi), .Y(div_result_20_) );
  MUX21X1_LVT div_U632 ( .A1(div_n_T_51_21_), .A2(div_n_T_51_85_), .S0(
        div_n308), .Y(div_result_21_) );
  MUX21X1_LVT div_U631 ( .A1(div_n_T_51_22_), .A2(div_n_T_51_86_), .S0(
        div_resHi), .Y(div_result_22_) );
  MUX21X1_LVT div_U630 ( .A1(div_n_T_51_23_), .A2(div_n_T_51_87_), .S0(
        div_resHi), .Y(div_result_23_) );
  NAND4X0_LVT div_U629 ( .A1(div_n548), .A2(div_n547), .A3(div_n546), .A4(
        div_n545), .Y(div_N417) );
  NAND2X0_LVT div_U628 ( .A1(div_negated_remainder[23]), .A2(div_n224), .Y(
        div_n545) );
  NAND2X0_LVT div_U627 ( .A1(div_n227), .A2(div_n_T_51_22_), .Y(div_n546) );
  AOI21X1_LVT div_U626 ( .A1(div_n679), .A2(div_n_T_87[23]), .A3(div_n544), 
        .Y(div_n547) );
  AO22X1_LVT div_U625 ( .A1(div_n235), .A2(io_fpu_fromint_data[23]), .A3(
        div_n223), .A4(div_n_T_51_31_), .Y(div_n544) );
  NAND2X0_LVT div_U624 ( .A1(div_n225), .A2(div_n_T_442[23]), .Y(div_n548) );
  NAND4X0_LVT div_U623 ( .A1(div_n543), .A2(div_n542), .A3(div_n541), .A4(
        div_n540), .Y(div_N416) );
  NAND2X0_LVT div_U622 ( .A1(div_negated_remainder[22]), .A2(div_n224), .Y(
        div_n540) );
  NAND2X0_LVT div_U621 ( .A1(div_n227), .A2(div_n_T_51_21_), .Y(div_n541) );
  AOI21X1_LVT div_U620 ( .A1(div_n679), .A2(div_n_T_87[22]), .A3(div_n539), 
        .Y(div_n542) );
  AO22X1_LVT div_U619 ( .A1(div_n235), .A2(io_fpu_fromint_data[22]), .A3(
        div_n223), .A4(div_n_T_51_30_), .Y(div_n539) );
  NAND2X0_LVT div_U618 ( .A1(div_n225), .A2(div_n_T_442[22]), .Y(div_n543) );
  NAND4X0_LVT div_U617 ( .A1(div_n538), .A2(div_n537), .A3(div_n536), .A4(
        div_n535), .Y(div_N415) );
  NAND2X0_LVT div_U616 ( .A1(div_negated_remainder[21]), .A2(div_n224), .Y(
        div_n535) );
  NAND2X0_LVT div_U615 ( .A1(div_n227), .A2(div_n_T_51_20_), .Y(div_n536) );
  AOI21X1_LVT div_U614 ( .A1(div_n679), .A2(div_n_T_87[21]), .A3(div_n534), 
        .Y(div_n537) );
  AO22X1_LVT div_U613 ( .A1(div_n235), .A2(io_fpu_fromint_data[21]), .A3(
        div_n223), .A4(div_n_T_51_29_), .Y(div_n534) );
  NAND2X0_LVT div_U612 ( .A1(div_n225), .A2(div_n_T_442[21]), .Y(div_n538) );
  NAND4X0_LVT div_U611 ( .A1(div_n533), .A2(div_n532), .A3(div_n531), .A4(
        div_n530), .Y(div_N414) );
  NAND2X0_LVT div_U610 ( .A1(div_negated_remainder[20]), .A2(div_n224), .Y(
        div_n530) );
  NAND2X0_LVT div_U609 ( .A1(div_n227), .A2(div_n_T_51_19_), .Y(div_n531) );
  AOI21X1_LVT div_U608 ( .A1(div_n679), .A2(div_n_T_87[20]), .A3(div_n529), 
        .Y(div_n532) );
  AO22X1_LVT div_U607 ( .A1(div_n235), .A2(io_fpu_fromint_data[20]), .A3(
        div_n223), .A4(div_n_T_51_28_), .Y(div_n529) );
  NAND2X0_LVT div_U606 ( .A1(div_n225), .A2(div_n_T_442[20]), .Y(div_n533) );
  NAND4X0_LVT div_U605 ( .A1(div_n528), .A2(div_n527), .A3(div_n526), .A4(
        div_n525), .Y(div_N413) );
  NAND2X0_LVT div_U604 ( .A1(div_negated_remainder[19]), .A2(div_n224), .Y(
        div_n525) );
  NAND2X0_LVT div_U603 ( .A1(div_n227), .A2(div_n_T_51_18_), .Y(div_n526) );
  AOI21X1_LVT div_U602 ( .A1(div_n679), .A2(div_n_T_87[19]), .A3(div_n524), 
        .Y(div_n527) );
  AO22X1_LVT div_U601 ( .A1(div_n235), .A2(io_fpu_fromint_data[19]), .A3(
        div_n223), .A4(div_n_T_51_27_), .Y(div_n524) );
  NAND2X0_LVT div_U600 ( .A1(div_n225), .A2(div_n_T_442[19]), .Y(div_n528) );
  NAND4X0_LVT div_U599 ( .A1(div_n523), .A2(div_n522), .A3(div_n521), .A4(
        div_n520), .Y(div_N412) );
  NAND2X0_LVT div_U598 ( .A1(div_negated_remainder[18]), .A2(div_n224), .Y(
        div_n520) );
  NAND2X0_LVT div_U597 ( .A1(div_n227), .A2(div_n_T_51_17_), .Y(div_n521) );
  AOI21X1_LVT div_U596 ( .A1(div_n679), .A2(div_n_T_87[18]), .A3(div_n519), 
        .Y(div_n522) );
  AO22X1_LVT div_U595 ( .A1(div_n235), .A2(io_fpu_fromint_data[18]), .A3(
        div_n223), .A4(div_n_T_51_26_), .Y(div_n519) );
  NAND2X0_LVT div_U594 ( .A1(div_n225), .A2(div_n_T_442[18]), .Y(div_n523) );
  MUX21X1_LVT div_U593 ( .A1(div_n_T_51_25_), .A2(div_n_T_51_89_), .S0(
        div_n308), .Y(div_result_25_) );
  MUX21X1_LVT div_U592 ( .A1(div_n_T_51_26_), .A2(div_n_T_51_90_), .S0(
        div_n308), .Y(div_result_26_) );
  MUX21X1_LVT div_U591 ( .A1(div_n_T_51_27_), .A2(div_n_T_51_91_), .S0(
        div_n308), .Y(div_result_27_) );
  MUX21X1_LVT div_U590 ( .A1(div_n_T_51_28_), .A2(div_n_T_51_92_), .S0(
        div_n308), .Y(div_result_28_) );
  MUX21X1_LVT div_U589 ( .A1(div_n_T_51_29_), .A2(div_n_T_51_93_), .S0(
        div_n308), .Y(div_result_29_) );
  NAND4X0_LVT div_U588 ( .A1(div_n518), .A2(div_n517), .A3(div_n516), .A4(
        div_n515), .Y(div_N425) );
  NAND2X0_LVT div_U587 ( .A1(div_negated_remainder[31]), .A2(div_n224), .Y(
        div_n515) );
  NAND2X0_LVT div_U586 ( .A1(div_n227), .A2(div_n_T_51_30_), .Y(div_n516) );
  AOI21X1_LVT div_U585 ( .A1(div_n679), .A2(div_n_T_87[31]), .A3(div_n514), 
        .Y(div_n517) );
  AO22X1_LVT div_U584 ( .A1(div_n235), .A2(io_fpu_fromint_data[31]), .A3(
        div_n223), .A4(div_n_T_51_39_), .Y(div_n514) );
  NAND2X0_LVT div_U583 ( .A1(div_n225), .A2(div_n_T_442[31]), .Y(div_n518) );
  NAND4X0_LVT div_U582 ( .A1(div_n513), .A2(div_n512), .A3(div_n511), .A4(
        div_n510), .Y(div_N424) );
  NAND2X0_LVT div_U581 ( .A1(div_negated_remainder[30]), .A2(div_n224), .Y(
        div_n510) );
  NAND2X0_LVT div_U580 ( .A1(div_n227), .A2(div_n_T_51_29_), .Y(div_n511) );
  AOI21X1_LVT div_U579 ( .A1(div_n679), .A2(div_n_T_87[30]), .A3(div_n509), 
        .Y(div_n512) );
  AO22X1_LVT div_U578 ( .A1(div_n235), .A2(io_fpu_fromint_data[30]), .A3(
        div_n223), .A4(div_n_T_51_38_), .Y(div_n509) );
  NAND2X0_LVT div_U577 ( .A1(div_n225), .A2(div_n_T_442[30]), .Y(div_n513) );
  NAND4X0_LVT div_U576 ( .A1(div_n508), .A2(div_n507), .A3(div_n506), .A4(
        div_n505), .Y(div_N423) );
  NAND2X0_LVT div_U575 ( .A1(div_negated_remainder[29]), .A2(div_n224), .Y(
        div_n505) );
  NAND2X0_LVT div_U574 ( .A1(div_n227), .A2(div_n_T_51_28_), .Y(div_n506) );
  AOI21X1_LVT div_U573 ( .A1(div_n679), .A2(div_n_T_87[29]), .A3(div_n504), 
        .Y(div_n507) );
  AO22X1_LVT div_U572 ( .A1(div_n235), .A2(io_fpu_fromint_data[29]), .A3(
        div_n223), .A4(div_n_T_51_37_), .Y(div_n504) );
  NAND2X0_LVT div_U571 ( .A1(div_n225), .A2(div_n_T_442[29]), .Y(div_n508) );
  NAND4X0_LVT div_U570 ( .A1(div_n503), .A2(div_n502), .A3(div_n501), .A4(
        div_n500), .Y(div_N422) );
  NAND2X0_LVT div_U569 ( .A1(div_negated_remainder[28]), .A2(div_n224), .Y(
        div_n500) );
  NAND2X0_LVT div_U568 ( .A1(div_n227), .A2(div_n_T_51_27_), .Y(div_n501) );
  AOI21X1_LVT div_U567 ( .A1(div_n679), .A2(div_n_T_87[28]), .A3(div_n499), 
        .Y(div_n502) );
  AO22X1_LVT div_U566 ( .A1(div_n235), .A2(io_fpu_fromint_data[28]), .A3(
        div_n223), .A4(div_n_T_51_36_), .Y(div_n499) );
  NAND2X0_LVT div_U565 ( .A1(div_n225), .A2(div_n_T_442[28]), .Y(div_n503) );
  NAND4X0_LVT div_U564 ( .A1(div_n498), .A2(div_n497), .A3(div_n496), .A4(
        div_n495), .Y(div_N421) );
  NAND2X0_LVT div_U563 ( .A1(div_negated_remainder[27]), .A2(div_n224), .Y(
        div_n495) );
  NAND2X0_LVT div_U562 ( .A1(div_n227), .A2(div_n_T_51_26_), .Y(div_n496) );
  AOI21X1_LVT div_U561 ( .A1(div_n679), .A2(div_n_T_87[27]), .A3(div_n494), 
        .Y(div_n497) );
  AO22X1_LVT div_U560 ( .A1(div_n235), .A2(io_fpu_fromint_data[27]), .A3(
        div_n223), .A4(div_n_T_51_35_), .Y(div_n494) );
  NAND2X0_LVT div_U559 ( .A1(div_n225), .A2(div_n_T_442[27]), .Y(div_n498) );
  NAND4X0_LVT div_U558 ( .A1(div_n493), .A2(div_n492), .A3(div_n491), .A4(
        div_n490), .Y(div_N420) );
  NAND2X0_LVT div_U557 ( .A1(div_negated_remainder[26]), .A2(div_n224), .Y(
        div_n490) );
  NAND2X0_LVT div_U556 ( .A1(div_n227), .A2(div_n_T_51_25_), .Y(div_n491) );
  AOI21X1_LVT div_U555 ( .A1(div_n679), .A2(div_n_T_87[26]), .A3(div_n489), 
        .Y(div_n492) );
  AO22X1_LVT div_U554 ( .A1(div_n235), .A2(io_fpu_fromint_data[26]), .A3(
        div_n223), .A4(div_n_T_51_34_), .Y(div_n489) );
  NAND2X0_LVT div_U553 ( .A1(div_n225), .A2(div_n_T_442[26]), .Y(div_n493) );
  MUX21X1_LVT div_U552 ( .A1(div_n_T_51_35_), .A2(div_n_T_51_99_), .S0(
        div_n308), .Y(div_result_35_) );
  NAND4X0_LVT div_U551 ( .A1(div_n488), .A2(div_n487), .A3(div_n486), .A4(
        div_n485), .Y(div_N433) );
  NAND2X0_LVT div_U550 ( .A1(div_negated_remainder[39]), .A2(div_n224), .Y(
        div_n485) );
  NAND2X0_LVT div_U549 ( .A1(div_n227), .A2(div_n_T_51_38_), .Y(div_n486) );
  AND4X1_LVT div_U548 ( .A1(div_n484), .A2(div_n658), .A3(div_n483), .A4(
        div_n482), .Y(div_n487) );
  NAND2X0_LVT div_U547 ( .A1(div_n655), .A2(io_fpu_fromint_data[39]), .Y(
        div_n482) );
  NAND2X0_LVT div_U546 ( .A1(div_n223), .A2(div_n_T_51_47_), .Y(div_n483) );
  NAND2X0_LVT div_U545 ( .A1(div_n_T_87[39]), .A2(div_n679), .Y(div_n484) );
  NAND2X0_LVT div_U544 ( .A1(div_n_T_442[39]), .A2(div_n225), .Y(div_n488) );
  NAND4X0_LVT div_U543 ( .A1(div_n481), .A2(div_n480), .A3(div_n479), .A4(
        div_n478), .Y(div_N432) );
  NAND2X0_LVT div_U542 ( .A1(div_negated_remainder[38]), .A2(div_n224), .Y(
        div_n478) );
  NAND2X0_LVT div_U541 ( .A1(div_n227), .A2(div_n_T_51_37_), .Y(div_n479) );
  AND4X1_LVT div_U540 ( .A1(div_n477), .A2(div_n658), .A3(div_n476), .A4(
        div_n475), .Y(div_n480) );
  NAND2X0_LVT div_U539 ( .A1(div_n655), .A2(io_fpu_fromint_data[38]), .Y(
        div_n475) );
  NAND2X0_LVT div_U538 ( .A1(div_n223), .A2(div_n_T_51_46_), .Y(div_n476) );
  NAND2X0_LVT div_U537 ( .A1(div_n_T_87[38]), .A2(div_n679), .Y(div_n477) );
  NAND2X0_LVT div_U536 ( .A1(div_n_T_442[38]), .A2(div_n225), .Y(div_n481) );
  NAND4X0_LVT div_U535 ( .A1(div_n474), .A2(div_n473), .A3(div_n472), .A4(
        div_n471), .Y(div_N431) );
  NAND2X0_LVT div_U534 ( .A1(div_negated_remainder[37]), .A2(div_n224), .Y(
        div_n471) );
  NAND2X0_LVT div_U533 ( .A1(div_n227), .A2(div_n_T_51_36_), .Y(div_n472) );
  AND4X1_LVT div_U532 ( .A1(div_n470), .A2(div_n658), .A3(div_n469), .A4(
        div_n468), .Y(div_n473) );
  NAND2X0_LVT div_U531 ( .A1(div_n655), .A2(io_fpu_fromint_data[37]), .Y(
        div_n468) );
  NAND2X0_LVT div_U530 ( .A1(div_n223), .A2(div_n_T_51_45_), .Y(div_n469) );
  NAND2X0_LVT div_U529 ( .A1(div_n_T_87[37]), .A2(div_n679), .Y(div_n470) );
  NAND2X0_LVT div_U528 ( .A1(div_n_T_442[37]), .A2(div_n157), .Y(div_n474) );
  NAND4X0_LVT div_U527 ( .A1(div_n467), .A2(div_n466), .A3(div_n465), .A4(
        div_n464), .Y(div_N430) );
  NAND2X0_LVT div_U526 ( .A1(div_negated_remainder[36]), .A2(div_n224), .Y(
        div_n464) );
  NAND2X0_LVT div_U525 ( .A1(div_n227), .A2(div_n_T_51_35_), .Y(div_n465) );
  AND4X1_LVT div_U524 ( .A1(div_n463), .A2(div_n658), .A3(div_n462), .A4(
        div_n461), .Y(div_n466) );
  NAND2X0_LVT div_U523 ( .A1(div_n655), .A2(io_fpu_fromint_data[36]), .Y(
        div_n461) );
  NAND2X0_LVT div_U522 ( .A1(div_n223), .A2(div_n_T_51_44_), .Y(div_n462) );
  NAND2X0_LVT div_U521 ( .A1(div_n_T_87[36]), .A2(div_n679), .Y(div_n463) );
  NAND2X0_LVT div_U520 ( .A1(div_n_T_442[36]), .A2(div_n225), .Y(div_n467) );
  NAND4X0_LVT div_U519 ( .A1(div_n460), .A2(div_n459), .A3(div_n458), .A4(
        div_n457), .Y(div_N429) );
  NAND2X0_LVT div_U518 ( .A1(div_negated_remainder[35]), .A2(div_n224), .Y(
        div_n457) );
  NAND2X0_LVT div_U517 ( .A1(div_n227), .A2(div_n_T_51_34_), .Y(div_n458) );
  AND4X1_LVT div_U516 ( .A1(div_n456), .A2(div_n658), .A3(div_n455), .A4(
        div_n454), .Y(div_n459) );
  NAND2X0_LVT div_U515 ( .A1(div_n655), .A2(io_fpu_fromint_data[35]), .Y(
        div_n454) );
  NAND2X0_LVT div_U514 ( .A1(div_n223), .A2(div_n_T_51_43_), .Y(div_n455) );
  NAND2X0_LVT div_U513 ( .A1(div_n_T_87[35]), .A2(div_n679), .Y(div_n456) );
  NAND2X0_LVT div_U512 ( .A1(div_n_T_442[35]), .A2(div_n157), .Y(div_n460) );
  NAND4X0_LVT div_U511 ( .A1(div_n453), .A2(div_n452), .A3(div_n451), .A4(
        div_n450), .Y(div_N428) );
  NAND2X0_LVT div_U510 ( .A1(div_negated_remainder[34]), .A2(div_n224), .Y(
        div_n450) );
  NAND2X0_LVT div_U509 ( .A1(div_n227), .A2(div_n_T_51_33_), .Y(div_n451) );
  AND4X1_LVT div_U508 ( .A1(div_n449), .A2(div_n658), .A3(div_n448), .A4(
        div_n447), .Y(div_n452) );
  NAND2X0_LVT div_U507 ( .A1(div_n655), .A2(io_fpu_fromint_data[34]), .Y(
        div_n447) );
  NAND2X0_LVT div_U506 ( .A1(div_n223), .A2(div_n_T_51_42_), .Y(div_n448) );
  NAND2X0_LVT div_U505 ( .A1(div_n_T_87[34]), .A2(div_n679), .Y(div_n449) );
  NAND2X0_LVT div_U504 ( .A1(div_n_T_442[34]), .A2(div_n225), .Y(div_n453) );
  NAND4X0_LVT div_U503 ( .A1(div_n446), .A2(div_n445), .A3(div_n444), .A4(
        div_n443), .Y(div_N441) );
  NAND2X0_LVT div_U502 ( .A1(div_negated_remainder[47]), .A2(div_n224), .Y(
        div_n443) );
  NAND2X0_LVT div_U501 ( .A1(div_n227), .A2(div_n_T_51_46_), .Y(div_n444) );
  AND4X1_LVT div_U500 ( .A1(div_n442), .A2(div_n658), .A3(div_n441), .A4(
        div_n440), .Y(div_n445) );
  NAND2X0_LVT div_U499 ( .A1(div_n655), .A2(io_fpu_fromint_data[47]), .Y(
        div_n440) );
  NAND2X0_LVT div_U498 ( .A1(div_n223), .A2(div_n_T_51_55_), .Y(div_n441) );
  NAND2X0_LVT div_U497 ( .A1(div_n_T_87[47]), .A2(div_n679), .Y(div_n442) );
  NAND2X0_LVT div_U496 ( .A1(div_n_T_442[47]), .A2(div_n225), .Y(div_n446) );
  NAND4X0_LVT div_U495 ( .A1(div_n439), .A2(div_n438), .A3(div_n437), .A4(
        div_n436), .Y(div_N440) );
  NAND2X0_LVT div_U494 ( .A1(div_negated_remainder[46]), .A2(div_n224), .Y(
        div_n436) );
  NAND2X0_LVT div_U493 ( .A1(div_n227), .A2(div_n_T_51_45_), .Y(div_n437) );
  AND4X1_LVT div_U492 ( .A1(div_n435), .A2(div_n658), .A3(div_n434), .A4(
        div_n433), .Y(div_n438) );
  NAND2X0_LVT div_U491 ( .A1(div_n655), .A2(io_fpu_fromint_data[46]), .Y(
        div_n433) );
  NAND2X0_LVT div_U490 ( .A1(div_n223), .A2(div_n_T_51_54_), .Y(div_n434) );
  NAND2X0_LVT div_U489 ( .A1(div_n_T_87[46]), .A2(div_n679), .Y(div_n435) );
  NAND2X0_LVT div_U488 ( .A1(div_n_T_442[46]), .A2(div_n225), .Y(div_n439) );
  NAND4X0_LVT div_U487 ( .A1(div_n432), .A2(div_n431), .A3(div_n430), .A4(
        div_n429), .Y(div_N439) );
  NAND2X0_LVT div_U486 ( .A1(div_negated_remainder[45]), .A2(div_n224), .Y(
        div_n429) );
  NAND2X0_LVT div_U485 ( .A1(div_n227), .A2(div_n_T_51_44_), .Y(div_n430) );
  AND4X1_LVT div_U484 ( .A1(div_n428), .A2(div_n658), .A3(div_n427), .A4(
        div_n426), .Y(div_n431) );
  NAND2X0_LVT div_U483 ( .A1(div_n655), .A2(io_fpu_fromint_data[45]), .Y(
        div_n426) );
  NAND2X0_LVT div_U482 ( .A1(div_n223), .A2(div_n_T_51_53_), .Y(div_n427) );
  NAND2X0_LVT div_U481 ( .A1(div_n_T_87[45]), .A2(div_n679), .Y(div_n428) );
  NAND2X0_LVT div_U480 ( .A1(div_n_T_442[45]), .A2(div_n225), .Y(div_n432) );
  NAND4X0_LVT div_U479 ( .A1(div_n425), .A2(div_n424), .A3(div_n423), .A4(
        div_n422), .Y(div_N438) );
  NAND2X0_LVT div_U478 ( .A1(div_negated_remainder[44]), .A2(div_n224), .Y(
        div_n422) );
  NAND2X0_LVT div_U477 ( .A1(div_n227), .A2(div_n_T_51_43_), .Y(div_n423) );
  AND4X1_LVT div_U476 ( .A1(div_n421), .A2(div_n658), .A3(div_n420), .A4(
        div_n419), .Y(div_n424) );
  NAND2X0_LVT div_U475 ( .A1(div_n655), .A2(io_fpu_fromint_data[44]), .Y(
        div_n419) );
  NAND2X0_LVT div_U474 ( .A1(div_n223), .A2(div_n_T_51_52_), .Y(div_n420) );
  NAND2X0_LVT div_U473 ( .A1(div_n_T_87[44]), .A2(div_n679), .Y(div_n421) );
  NAND2X0_LVT div_U472 ( .A1(div_n_T_442[44]), .A2(div_n225), .Y(div_n425) );
  NAND4X0_LVT div_U471 ( .A1(div_n418), .A2(div_n417), .A3(div_n416), .A4(
        div_n415), .Y(div_N437) );
  NAND2X0_LVT div_U470 ( .A1(div_negated_remainder[43]), .A2(div_n224), .Y(
        div_n415) );
  NAND2X0_LVT div_U469 ( .A1(div_n227), .A2(div_n_T_51_42_), .Y(div_n416) );
  AND4X1_LVT div_U468 ( .A1(div_n414), .A2(div_n658), .A3(div_n413), .A4(
        div_n412), .Y(div_n417) );
  NAND2X0_LVT div_U467 ( .A1(div_n655), .A2(io_fpu_fromint_data[43]), .Y(
        div_n412) );
  NAND2X0_LVT div_U466 ( .A1(div_n223), .A2(div_n_T_51_51_), .Y(div_n413) );
  NAND2X0_LVT div_U465 ( .A1(div_n_T_87[43]), .A2(div_n679), .Y(div_n414) );
  NAND2X0_LVT div_U464 ( .A1(div_n_T_442[43]), .A2(div_n225), .Y(div_n418) );
  NAND4X0_LVT div_U463 ( .A1(div_n411), .A2(div_n410), .A3(div_n409), .A4(
        div_n408), .Y(div_N436) );
  NAND2X0_LVT div_U462 ( .A1(div_negated_remainder[42]), .A2(div_n224), .Y(
        div_n408) );
  NAND2X0_LVT div_U461 ( .A1(div_n227), .A2(div_n_T_51_41_), .Y(div_n409) );
  AND4X1_LVT div_U460 ( .A1(div_n407), .A2(div_n658), .A3(div_n406), .A4(
        div_n405), .Y(div_n410) );
  NAND2X0_LVT div_U459 ( .A1(div_n655), .A2(io_fpu_fromint_data[42]), .Y(
        div_n405) );
  NAND2X0_LVT div_U458 ( .A1(div_n223), .A2(div_n_T_51_50_), .Y(div_n406) );
  NAND2X0_LVT div_U457 ( .A1(div_n_T_87[42]), .A2(div_n679), .Y(div_n407) );
  NAND2X0_LVT div_U456 ( .A1(div_n_T_442[42]), .A2(div_n225), .Y(div_n411) );
  NAND4X0_LVT div_U455 ( .A1(div_n404), .A2(div_n403), .A3(div_n402), .A4(
        div_n401), .Y(div_N449) );
  NAND2X0_LVT div_U454 ( .A1(div_negated_remainder[55]), .A2(div_n224), .Y(
        div_n401) );
  NAND2X0_LVT div_U453 ( .A1(div_n227), .A2(div_n_T_51_54_), .Y(div_n402) );
  AND4X1_LVT div_U452 ( .A1(div_n400), .A2(div_n658), .A3(div_n399), .A4(
        div_n398), .Y(div_n403) );
  NAND2X0_LVT div_U451 ( .A1(div_n655), .A2(io_fpu_fromint_data[55]), .Y(
        div_n398) );
  NAND2X0_LVT div_U450 ( .A1(div_n223), .A2(div_n_T_51_63_), .Y(div_n399) );
  NAND2X0_LVT div_U449 ( .A1(div_n_T_87[55]), .A2(div_n679), .Y(div_n400) );
  NAND2X0_LVT div_U448 ( .A1(div_n_T_442[55]), .A2(div_n157), .Y(div_n404) );
  NAND4X0_LVT div_U447 ( .A1(div_n397), .A2(div_n396), .A3(div_n395), .A4(
        div_n394), .Y(div_N448) );
  NAND2X0_LVT div_U446 ( .A1(div_negated_remainder[54]), .A2(div_n224), .Y(
        div_n394) );
  NAND2X0_LVT div_U445 ( .A1(div_n227), .A2(div_n_T_51_53_), .Y(div_n395) );
  AND4X1_LVT div_U444 ( .A1(div_n393), .A2(div_n658), .A3(div_n392), .A4(
        div_n391), .Y(div_n396) );
  NAND2X0_LVT div_U443 ( .A1(div_n655), .A2(io_fpu_fromint_data[54]), .Y(
        div_n391) );
  NAND2X0_LVT div_U442 ( .A1(div_n223), .A2(div_n_T_51_62_), .Y(div_n392) );
  NAND2X0_LVT div_U441 ( .A1(div_n_T_87[54]), .A2(div_n679), .Y(div_n393) );
  NAND2X0_LVT div_U440 ( .A1(div_n_T_442[54]), .A2(div_n157), .Y(div_n397) );
  NAND4X0_LVT div_U439 ( .A1(div_n390), .A2(div_n389), .A3(div_n388), .A4(
        div_n387), .Y(div_N447) );
  NAND2X0_LVT div_U438 ( .A1(div_negated_remainder[53]), .A2(div_n224), .Y(
        div_n387) );
  NAND2X0_LVT div_U437 ( .A1(div_n227), .A2(div_n_T_51_52_), .Y(div_n388) );
  AND4X1_LVT div_U436 ( .A1(div_n386), .A2(div_n658), .A3(div_n385), .A4(
        div_n384), .Y(div_n389) );
  NAND2X0_LVT div_U435 ( .A1(div_n655), .A2(io_fpu_fromint_data[53]), .Y(
        div_n384) );
  NAND2X0_LVT div_U434 ( .A1(div_n223), .A2(div_n_T_51_61_), .Y(div_n385) );
  NAND2X0_LVT div_U433 ( .A1(div_n_T_87[53]), .A2(div_n679), .Y(div_n386) );
  NAND2X0_LVT div_U432 ( .A1(div_n_T_442[53]), .A2(div_n225), .Y(div_n390) );
  NAND4X0_LVT div_U431 ( .A1(div_n383), .A2(div_n382), .A3(div_n381), .A4(
        div_n380), .Y(div_N445) );
  NAND2X0_LVT div_U430 ( .A1(div_negated_remainder[51]), .A2(div_n224), .Y(
        div_n380) );
  NAND2X0_LVT div_U429 ( .A1(div_n227), .A2(div_n_T_51_50_), .Y(div_n381) );
  AND4X1_LVT div_U428 ( .A1(div_n379), .A2(div_n658), .A3(div_n378), .A4(
        div_n377), .Y(div_n382) );
  NAND2X0_LVT div_U427 ( .A1(div_n655), .A2(io_fpu_fromint_data[51]), .Y(
        div_n377) );
  NAND2X0_LVT div_U426 ( .A1(div_n223), .A2(div_n_T_51_59_), .Y(div_n378) );
  NAND2X0_LVT div_U425 ( .A1(div_n_T_87[51]), .A2(div_n679), .Y(div_n379) );
  NAND2X0_LVT div_U424 ( .A1(div_n_T_442[51]), .A2(div_n225), .Y(div_n383) );
  NAND4X0_LVT div_U423 ( .A1(div_n376), .A2(div_n375), .A3(div_n374), .A4(
        div_n373), .Y(div_N444) );
  NAND2X0_LVT div_U422 ( .A1(div_negated_remainder[50]), .A2(div_n224), .Y(
        div_n373) );
  NAND2X0_LVT div_U421 ( .A1(div_n227), .A2(div_n_T_51_49_), .Y(div_n374) );
  AND4X1_LVT div_U420 ( .A1(div_n372), .A2(div_n658), .A3(div_n371), .A4(
        div_n370), .Y(div_n375) );
  NAND2X0_LVT div_U419 ( .A1(div_n655), .A2(io_fpu_fromint_data[50]), .Y(
        div_n370) );
  NAND2X0_LVT div_U418 ( .A1(div_n223), .A2(div_n_T_51_58_), .Y(div_n371) );
  NAND2X0_LVT div_U417 ( .A1(div_n_T_87[50]), .A2(div_n679), .Y(div_n372) );
  NAND2X0_LVT div_U416 ( .A1(div_n_T_442[50]), .A2(div_n225), .Y(div_n376) );
  NAND4X0_LVT div_U415 ( .A1(div_n369), .A2(div_n368), .A3(div_n367), .A4(
        div_n366), .Y(div_N455) );
  NAND2X0_LVT div_U414 ( .A1(div_n_T_442[61]), .A2(div_n225), .Y(div_n366) );
  NAND2X0_LVT div_U413 ( .A1(div_n227), .A2(div_n_T_51_60_), .Y(div_n367) );
  AND4X1_LVT div_U412 ( .A1(div_n365), .A2(div_n658), .A3(div_n364), .A4(
        div_n363), .Y(div_n368) );
  NAND2X0_LVT div_U411 ( .A1(div_n655), .A2(io_fpu_fromint_data[61]), .Y(
        div_n363) );
  NAND2X0_LVT div_U410 ( .A1(div_n_T_87[61]), .A2(div_n679), .Y(div_n364) );
  NAND2X0_LVT div_U409 ( .A1(div_n_T_65[5]), .A2(div_n223), .Y(div_n365) );
  NAND2X0_LVT div_U408 ( .A1(div_negated_remainder[61]), .A2(div_n224), .Y(
        div_n369) );
  NAND4X0_LVT div_U407 ( .A1(div_n362), .A2(div_n361), .A3(div_n360), .A4(
        div_n359), .Y(div_N454) );
  NAND2X0_LVT div_U406 ( .A1(div_n_T_442[60]), .A2(div_n225), .Y(div_n359) );
  NAND2X0_LVT div_U405 ( .A1(div_n227), .A2(div_n_T_51_59_), .Y(div_n360) );
  AND4X1_LVT div_U404 ( .A1(div_n358), .A2(div_n658), .A3(div_n357), .A4(
        div_n356), .Y(div_n361) );
  NAND2X0_LVT div_U403 ( .A1(div_n655), .A2(io_fpu_fromint_data[60]), .Y(
        div_n356) );
  NAND2X0_LVT div_U402 ( .A1(div_n_T_87[60]), .A2(div_n679), .Y(div_n357) );
  NAND2X0_LVT div_U401 ( .A1(div_n_T_65[4]), .A2(div_n223), .Y(div_n358) );
  NAND2X0_LVT div_U400 ( .A1(div_negated_remainder[60]), .A2(div_n224), .Y(
        div_n362) );
  NAND4X0_LVT div_U399 ( .A1(div_n355), .A2(div_n354), .A3(div_n353), .A4(
        div_n352), .Y(div_N453) );
  NAND2X0_LVT div_U398 ( .A1(div_n_T_442[59]), .A2(div_n157), .Y(div_n352) );
  NAND2X0_LVT div_U397 ( .A1(div_n227), .A2(div_n_T_51_58_), .Y(div_n353) );
  AND4X1_LVT div_U396 ( .A1(div_n351), .A2(div_n658), .A3(div_n350), .A4(
        div_n349), .Y(div_n354) );
  NAND2X0_LVT div_U395 ( .A1(div_n655), .A2(io_fpu_fromint_data[59]), .Y(
        div_n349) );
  NAND2X0_LVT div_U394 ( .A1(div_n_T_87[59]), .A2(div_n679), .Y(div_n350) );
  NAND2X0_LVT div_U393 ( .A1(div_n_T_65[3]), .A2(div_n223), .Y(div_n351) );
  NAND2X0_LVT div_U392 ( .A1(div_negated_remainder[59]), .A2(div_n224), .Y(
        div_n355) );
  NAND4X0_LVT div_U391 ( .A1(div_n348), .A2(div_n347), .A3(div_n346), .A4(
        div_n345), .Y(div_N452) );
  NAND2X0_LVT div_U390 ( .A1(div_n227), .A2(div_n_T_51_57_), .Y(div_n345) );
  NAND2X0_LVT div_U389 ( .A1(div_n_T_442[58]), .A2(div_n225), .Y(div_n346) );
  AND4X1_LVT div_U388 ( .A1(div_n341), .A2(div_n658), .A3(div_n340), .A4(
        div_n339), .Y(div_n347) );
  NAND2X0_LVT div_U387 ( .A1(div_n655), .A2(io_fpu_fromint_data[58]), .Y(
        div_n339) );
  NAND2X0_LVT div_U386 ( .A1(div_n223), .A2(div_n_T_65[2]), .Y(div_n340) );
  AND3X1_LVT div_U385 ( .A1(div_n235), .A2(div_n787), .A3(div_n336), .Y(
        div_n337) );
  NAND2X0_LVT div_U384 ( .A1(div_n_T_87[58]), .A2(div_n679), .Y(div_n341) );
  NAND2X0_LVT div_U383 ( .A1(div_negated_remainder[58]), .A2(div_n224), .Y(
        div_n348) );
  AO22X1_LVT div_U382 ( .A1(div_isHi), .A2(div_n335), .A3(div_n308), .A4(
        div_n979), .Y(div_n794) );
  INVX1_LVT div_U381 ( .A(div_n752), .Y(div_n335) );
  NOR2X0_LVT div_U380 ( .A1(div_n782), .A2(div_n978), .Y(div_n752) );
  AO21X1_LVT div_U379 ( .A1(div_n783), .A2(div_n334), .A3(div_n679), .Y(
        div_n978) );
  AND4X1_LVT div_U378 ( .A1(div_n236), .A2(div_n239), .A3(div_n238), .A4(
        div_n237), .Y(div_n779) );
  AND4X1_LVT div_U377 ( .A1(div_n182), .A2(div_n243), .A3(div_n240), .A4(
        div_n241), .Y(div_n732) );
  AND4X1_LVT div_U376 ( .A1(div_n290), .A2(div_n293), .A3(div_n292), .A4(
        div_n291), .Y(div_n781) );
  NAND2X0_LVT div_U375 ( .A1(div_n332), .A2(div_n780), .Y(div_n1000) );
  AND4X1_LVT div_U374 ( .A1(div_n283), .A2(div_n281), .A3(div_n284), .A4(
        div_n282), .Y(div_n780) );
  AND4X1_LVT div_U373 ( .A1(div_n147), .A2(div_n186), .A3(div_n153), .A4(
        div_n286), .Y(div_n332) );
  INVX1_LVT div_U372 ( .A(div_n790), .Y(div_n334) );
  AO222X1_LVT div_U371 ( .A1(div_n783), .A2(div_n_T_65[70]), .A3(
        div_subtractor_62_), .A4(div_n226), .A5(div_n_T_51_125_), .A6(div_n931), .Y(div_N522) );
  NAND3X0_LVT div_U370 ( .A1(div_n778), .A2(div_n614), .A3(div_n613), .Y(
        div_n790) );
  NOR2X0_LVT div_U369 ( .A1(div_n_T_69_9_), .A2(div_n_T_69_8_), .Y(div_n613)
         );
  INVX1_LVT div_U368 ( .A(div_n800), .Y(div_n778) );
  OR2X1_LVT div_U367 ( .A1(div_n210), .A2(div_n795), .Y(div_n800) );
  NAND2X0_LVT div_U366 ( .A1(div_n_T_69_4_), .A2(div_n300), .Y(div_n795) );
  NAND2X0_LVT div_U365 ( .A1(div_n792), .A2(div_subtractor_64_), .Y(div_n344)
         );
  NAND3X0_LVT div_U364 ( .A1(div_n330), .A2(div_n329), .A3(div_n328), .Y(
        div_N284) );
  AO21X1_LVT div_U363 ( .A1(div_n203), .A2(div_n230), .A3(div_n327), .Y(
        div_n328) );
  OR3X1_LVT div_U362 ( .A1(reset), .A2(div_n199), .A3(div_n326), .Y(div_n329)
         );
  OA21X1_LVT div_U361 ( .A1(div_n325), .A2(div_n616), .A3(alu_io_fn[2]), .Y(
        div_n326) );
  AND2X1_LVT div_U360 ( .A1(div_n324), .A2(div_n323), .Y(div_n616) );
  MUX21X1_LVT div_U359 ( .A1(div_n785), .A2(div_n786), .S0(alu_io_fn[2]), .Y(
        div_n323) );
  NAND2X0_LVT div_U358 ( .A1(div_n680), .A2(div_n212), .Y(div_n330) );
  AND2X1_LVT div_U357 ( .A1(div_n753), .A2(div_n782), .Y(div_n680) );
  AND3X1_LVT div_U356 ( .A1(div_n322), .A2(div_n_T_69_9_), .A3(div_n343), .Y(
        div_n782) );
  INVX1_LVT div_U355 ( .A(div_n321), .Y(div_n322) );
  NAND3X0_LVT div_U354 ( .A1(div_n319), .A2(div_n199), .A3(div_n309), .Y(
        div_n320) );
  NAND2X0_LVT div_U353 ( .A1(div_io_resp_ready), .A2(div_io_resp_valid), .Y(
        div_n319) );
  AND2X1_LVT div_U352 ( .A1(div_n184), .A2(div_n154), .Y(div_io_resp_valid) );
  NAND2X0_LVT div_U351 ( .A1(div_n318), .A2(div_n317), .Y(div_n793) );
  MUX21X1_LVT div_U350 ( .A1(div_n316), .A2(div_n315), .S0(div_n314), .Y(
        div_n317) );
  NAND3X0_LVT div_U349 ( .A1(div_n324), .A2(div_n786), .A3(div_n785), .Y(
        div_n314) );
  NAND2X0_LVT div_U348 ( .A1(div_n325), .A2(div_n235), .Y(div_n315) );
  AND2X1_LVT div_U347 ( .A1(div_n313), .A2(div_n336), .Y(div_n325) );
  AO21X1_LVT div_U346 ( .A1(div_n784), .A2(div_n785), .A3(div_n786), .Y(
        div_n336) );
  MUX21X1_LVT div_U345 ( .A1(io_fpu_fromint_data[31]), .A2(
        io_fpu_fromint_data[63]), .S0(alu_io_dw), .Y(div_n313) );
  OA22X1_LVT div_U344 ( .A1(div_n222), .A2(io_fpu_fromint_data[63]), .A3(
        div_n312), .A4(io_fpu_fromint_data[31]), .Y(div_n316) );
  AND2X1_LVT div_U343 ( .A1(div_n235), .A2(div_n787), .Y(div_n615) );
  NAND3X0_LVT div_U342 ( .A1(div_n311), .A2(div_neg_out), .A3(div_n199), .Y(
        div_n318) );
  AND3X1_LVT div_U341 ( .A1(div_n219), .A2(div_n220), .A3(div_n217), .Y(
        div_io_req_ready) );
  NAND4X0_LVT div_U340 ( .A1(div_n310), .A2(div_n342), .A3(div_n150), .A4(
        div_n189), .Y(div_n311) );
  INVX1_LVT div_U339 ( .A(div_n980), .Y(div_n342) );
  OR3X1_LVT div_U338 ( .A1(div_n_T_69_8_), .A2(div_n331), .A3(div_n789), .Y(
        div_n321) );
  OR2X1_LVT div_U337 ( .A1(div_n_T_69_6_), .A2(div_n_T_69_7_), .Y(div_n331) );
  NAND3X0_LVT div_U336 ( .A1(div_n204), .A2(div_n148), .A3(div_n210), .Y(
        div_n789) );
  AND2X1_LVT div_U335 ( .A1(div_n184), .A2(div_n217), .Y(div_n750) );
  NAND3X0_LVT div_U334 ( .A1(div_n800), .A2(div_n805), .A3(div_n221), .Y(
        div_n798) );
  NAND2X0_LVT div_U333 ( .A1(div_n210), .A2(div_n795), .Y(div_n221) );
  NAND3X0_LVT div_U332 ( .A1(div_n211), .A2(div_n216), .A3(div_n218), .Y(
        div_n_T_272[3]) );
  NAND2X0_LVT div_U331 ( .A1(div_n969), .A2(div_n966), .Y(div_n218) );
  NAND3X0_LVT div_U330 ( .A1(div_n158), .A2(div_n773), .A3(div_n215), .Y(
        div_n_T_429[3]) );
  NAND2X0_LVT div_U329 ( .A1(div_n1002), .A2(div_n999), .Y(div_n215) );
  NAND3X0_LVT div_U328 ( .A1(div_n213), .A2(div_n151), .A3(div_n214), .Y(
        div_n_T_429[0]) );
  NAND2X0_LVT div_U327 ( .A1(div_n1001), .A2(div_n996), .Y(div_n214) );
  AOI22X1_LVT div_U326 ( .A1(div_n1002), .A2(div_n995), .A3(div_n1003), .A4(
        div_n994), .Y(div_n213) );
  AOI22X1_LVT div_U325 ( .A1(div_n965), .A2(div_n964), .A3(div_n963), .A4(
        div_n962), .Y(div_n211) );
  NAND2X0_LVT div_U324 ( .A1(div_n783), .A2(div_n338), .Y(div_n201) );
  NBUFFX2_LVT div_U323 ( .A(div_n_T_51_4_), .Y(div_n306) );
  NBUFFX2_LVT div_U322 ( .A(div_n_T_51_1_), .Y(div_n303) );
  NBUFFX2_LVT div_U321 ( .A(div_n_T_51_3_), .Y(div_n305) );
  NBUFFX2_LVT div_U320 ( .A(div_n_T_51_0_), .Y(div_n302) );
  INVX1_LVT div_U319 ( .A(div_n783), .Y(div_n230) );
  AOI22X1_LVT div_U318 ( .A1(div_n976), .A2(div_n997), .A3(div_n1001), .A4(
        div_n1000), .Y(div_n158) );
  NBUFFX2_LVT div_U317 ( .A(div_n_T_51_6_), .Y(div_n307) );
  AND4X1_LVT div_U316 ( .A1(div_n758), .A2(div_n983), .A3(div_n982), .A4(
        div_n981), .Y(div_n151) );
  INVX1_LVT div_U315 ( .A(div_n_T_273_5_), .Y(div_n965) );
  INVX1_LVT div_U314 ( .A(div_n_T_430_5_), .Y(div_n976) );
  INVX1_LVT div_U313 ( .A(div_n990), .Y(div_n1003) );
  INVX1_LVT div_U312 ( .A(div_n804), .Y(div_n803) );
  NOR4X1_LVT div_U311 ( .A1(div_n978), .A2(div_n977), .A3(div_n235), .A4(
        div_n782), .Y(div_n979) );
  NAND2X0_LVT div_U310 ( .A1(n9422), .A2(div_io_req_ready), .Y(div_n199) );
  AND2X1_LVT div_U309 ( .A1(div_n750), .A2(div_n150), .Y(div_n343) );
  NAND2X0_LVT div_U308 ( .A1(div_n150), .A2(div_n219), .Y(div_n203) );
  XOR2X2_LVT div_U307 ( .A1(div_n300), .A2(div_n_T_69_4_), .Y(div_n_T_85_4_)
         );
  INVX1_LVT div_U306 ( .A(div_n206), .Y(div_n244) );
  NAND2X0_LVT div_U305 ( .A1(div_n220), .A2(div_n244), .Y(div_n209) );
  NBUFFX2_LVT div_U304 ( .A(div_resHi), .Y(div_n308) );
  MUX21X1_LVT div_U303 ( .A1(div_n_T_51_50_), .A2(div_n_T_51_114_), .S0(
        div_n308), .Y(div_result_50_) );
  MUX21X1_LVT div_U302 ( .A1(div_n_T_51_61_), .A2(div_n_T_51_125_), .S0(
        div_n308), .Y(div_result_61_) );
  MUX21X1_LVT div_U301 ( .A1(div_n_T_51_55_), .A2(div_n_T_51_119_), .S0(
        div_n308), .Y(div_result_55_) );
  MUX21X1_LVT div_U300 ( .A1(div_n_T_51_59_), .A2(div_n_T_51_123_), .S0(
        div_n308), .Y(div_result_59_) );
  MUX21X1_LVT div_U299 ( .A1(div_n_T_51_63_), .A2(div_n_T_51_127_), .S0(
        div_n308), .Y(div_result_63_) );
  MUX21X1_LVT div_U298 ( .A1(div_n_T_51_31_), .A2(div_n_T_51_95_), .S0(
        div_n308), .Y(div_result_31_) );
  AO22X1_LVT div_U297 ( .A1(div_n146), .A2(div_result_63_), .A3(div_n209), 
        .A4(div_result_31_), .Y(div_io_resp_bits_data[31]) );
  MUX21X1_LVT div_U296 ( .A1(div_n_T_51_62_), .A2(div_n_T_51_126_), .S0(
        div_n308), .Y(div_result_62_) );
  MUX21X1_LVT div_U295 ( .A1(div_n_T_51_30_), .A2(div_n_T_51_94_), .S0(
        div_n308), .Y(div_result_30_) );
  MUX21X1_LVT div_U294 ( .A1(div_n_T_51_54_), .A2(div_n_T_51_118_), .S0(
        div_n308), .Y(div_result_54_) );
  MUX21X1_LVT div_U293 ( .A1(div_n_T_51_32_), .A2(div_n_T_51_96_), .S0(
        div_n308), .Y(div_result_32_) );
  MUX21X1_LVT div_U292 ( .A1(div_n_T_51_36_), .A2(div_n_T_51_100_), .S0(
        div_n308), .Y(div_result_36_) );
  MUX21X1_LVT div_U291 ( .A1(div_n_T_51_60_), .A2(div_n_T_51_124_), .S0(
        div_n308), .Y(div_result_60_) );
  MUX21X1_LVT div_U290 ( .A1(div_n_T_51_43_), .A2(div_n_T_51_107_), .S0(
        div_n308), .Y(div_result_43_) );
  MUX21X1_LVT div_U289 ( .A1(div_n_T_51_34_), .A2(div_n_T_51_98_), .S0(
        div_n308), .Y(div_result_34_) );
  INVX1_LVT div_U288 ( .A(div_n208), .Y(div_n304) );
  MUX21X1_LVT div_U287 ( .A1(div_n_T_51_44_), .A2(div_n_T_51_108_), .S0(
        div_n308), .Y(div_result_44_) );
  MUX21X1_LVT div_U286 ( .A1(div_n_T_51_41_), .A2(div_n_T_51_105_), .S0(
        div_n308), .Y(div_result_41_) );
  MUX21X1_LVT div_U285 ( .A1(div_n_T_51_38_), .A2(div_n_T_51_102_), .S0(
        div_n308), .Y(div_result_38_) );
  MUX21X1_LVT div_U284 ( .A1(div_n_T_51_39_), .A2(div_n_T_51_103_), .S0(
        div_n308), .Y(div_result_39_) );
  MUX21X1_LVT div_U283 ( .A1(div_n_T_51_45_), .A2(div_n_T_51_109_), .S0(
        div_n308), .Y(div_result_45_) );
  INVX1_LVT div_U282 ( .A(div_n156), .Y(div_n242) );
  MUX21X1_LVT div_U281 ( .A1(div_n_T_51_42_), .A2(div_n_T_51_106_), .S0(
        div_n308), .Y(div_result_42_) );
  MUX21X1_LVT div_U280 ( .A1(div_n_T_51_53_), .A2(div_n_T_51_117_), .S0(
        div_n308), .Y(div_result_53_) );
  MUX21X1_LVT div_U279 ( .A1(div_n_T_51_52_), .A2(div_n_T_51_116_), .S0(
        div_n308), .Y(div_result_52_) );
  MUX21X1_LVT div_U278 ( .A1(div_n_T_51_49_), .A2(div_n_T_51_113_), .S0(
        div_n308), .Y(div_result_49_) );
  MUX21X1_LVT div_U277 ( .A1(div_n_T_51_40_), .A2(div_n_T_51_104_), .S0(
        div_n308), .Y(div_result_40_) );
  MUX21X1_LVT div_U276 ( .A1(div_n_T_51_46_), .A2(div_n_T_51_110_), .S0(
        div_n308), .Y(div_result_46_) );
  MUX21X1_LVT div_U275 ( .A1(div_n_T_51_14_), .A2(div_n_T_51_78_), .S0(
        div_n308), .Y(div_result_14_) );
  MUX21X1_LVT div_U274 ( .A1(div_n_T_51_58_), .A2(div_n_T_51_122_), .S0(
        div_n308), .Y(div_result_58_) );
  MUX21X1_LVT div_U273 ( .A1(div_n_T_51_57_), .A2(div_n_T_51_121_), .S0(
        div_n308), .Y(div_result_57_) );
  MUX21X1_LVT div_U272 ( .A1(div_n_T_51_47_), .A2(div_n_T_51_111_), .S0(
        div_n308), .Y(div_result_47_) );
  MUX21X1_LVT div_U271 ( .A1(div_n_T_51_48_), .A2(div_n_T_51_112_), .S0(
        div_n308), .Y(div_result_48_) );
  MUX21X1_LVT div_U270 ( .A1(div_n_T_51_37_), .A2(div_n_T_51_101_), .S0(
        div_n308), .Y(div_result_37_) );
  MUX21X1_LVT div_U269 ( .A1(div_n_T_51_33_), .A2(div_n_T_51_97_), .S0(
        div_n308), .Y(div_result_33_) );
  MUX21X1_LVT div_U268 ( .A1(div_n_T_51_56_), .A2(div_n_T_51_120_), .S0(
        div_n308), .Y(div_result_56_) );
  MUX21X1_LVT div_U267 ( .A1(div_n_T_51_51_), .A2(div_n_T_51_115_), .S0(
        div_n308), .Y(div_result_51_) );
  MUX21X1_LVT div_U266 ( .A1(div_n_T_51_24_), .A2(div_n_T_51_88_), .S0(
        div_n308), .Y(div_result_24_) );
  MUX21X1_LVT div_U265 ( .A1(div_n_T_51_16_), .A2(div_n_T_51_80_), .S0(
        div_n308), .Y(div_result_16_) );
  INVX1_LVT div_U264 ( .A(div_n199), .Y(div_n235) );
  INVX1_LVT div_U263 ( .A(div_n203), .Y(div_n224) );
  AND2X1_LVT div_U262 ( .A1(div_n750), .A2(div_n220), .Y(div_n783) );
  AND2X1_LVT div_U261 ( .A1(div_n774), .A2(div_n683), .Y(div_n773) );
  OR2X1_LVT div_U260 ( .A1(div_n_T_69_9_), .A2(div_n321), .Y(div_n980) );
  AND2X1_LVT div_U259 ( .A1(div_n333), .A2(div_n783), .Y(div_n679) );
  AND2X1_LVT div_U258 ( .A1(div_n224), .A2(div_n217), .Y(div_n754) );
  NBUFFX2_LVT div_U257 ( .A(div_n_T_59_8_), .Y(div_n301) );
  INVX1_LVT div_U256 ( .A(div_n775), .Y(div_n997) );
  OR3X1_LVT div_U255 ( .A1(div_n970), .A2(div_n972), .A3(div_n998), .Y(
        div_n_T_430_5_) );
  NBUFFX2_LVT div_U254 ( .A(div_n157), .Y(div_n225) );
  INVX1_LVT div_U253 ( .A(div_n_T_434_2_), .Y(div_n167) );
  INVX1_LVT div_U252 ( .A(div_n_T_434_1_), .Y(div_n166) );
  INVX1_LVT div_U251 ( .A(div_n_T_434_0_), .Y(div_n171) );
  OAI21X1_LVT div_U250 ( .A1(div_n980), .A2(div_n344), .A3(div_n343), .Y(
        div_n200) );
  INVX1_LVT div_U249 ( .A(div_n200), .Y(div_n227) );
  INVX1_LVT div_U248 ( .A(div_n201), .Y(div_n223) );
  AND2X1_LVT div_U247 ( .A1(div_n789), .A2(div_n605), .Y(div_n_T_85_5_) );
  AND2X1_LVT div_U246 ( .A1(div_n235), .A2(alu_io_dw), .Y(div_n655) );
  AND2X1_LVT div_U245 ( .A1(div_subtractor_64_), .A2(div_n227), .Y(div_n931)
         );
  INVX1_LVT div_U244 ( .A(div_n207), .Y(div_n226) );
  NBUFFX2_LVT div_U243 ( .A(div_net34705), .Y(div_n245) );
  NBUFFX2_LVT div_U242 ( .A(div_net34705), .Y(div_n262) );
  NBUFFX2_LVT div_U241 ( .A(div_net34705), .Y(div_n253) );
  NBUFFX2_LVT div_U240 ( .A(div_net34705), .Y(div_n265) );
  NBUFFX2_LVT div_U239 ( .A(div_net34705), .Y(div_n271) );
  NBUFFX2_LVT div_U238 ( .A(div_net34705), .Y(div_n276) );
  NBUFFX2_LVT div_U237 ( .A(div_net34705), .Y(div_n279) );
  NBUFFX2_LVT div_U236 ( .A(div_net34705), .Y(div_n280) );
  NBUFFX2_LVT div_U235 ( .A(div_net34705), .Y(div_n285) );
  NBUFFX2_LVT div_U234 ( .A(div_net34705), .Y(div_n287) );
  NBUFFX2_LVT div_U233 ( .A(div_net34705), .Y(div_n288) );
  NBUFFX2_LVT div_U232 ( .A(div_net34684), .Y(div_n298) );
  NBUFFX2_LVT div_U231 ( .A(div_net34684), .Y(div_n295) );
  NBUFFX2_LVT div_U230 ( .A(div_net34684), .Y(div_n297) );
  NBUFFX2_LVT div_U229 ( .A(div_net34684), .Y(div_n294) );
  NBUFFX2_LVT div_U228 ( .A(div_net34684), .Y(div_n289) );
  NBUFFX2_LVT div_U227 ( .A(div_net34684), .Y(div_n299) );
  NOR2X1_LVT div_U226 ( .A1(div_divisor_27_), .A2(div_divisor_25_), .Y(
        div_n687) );
  NOR2X1_LVT div_U225 ( .A1(div_divisor_11_), .A2(div_divisor_9_), .Y(div_n699) );
  NOR2X1_LVT div_U224 ( .A1(div_divisor_43_), .A2(div_divisor_41_), .Y(
        div_n686) );
  INVX0_LVT div_U223 ( .A(div_n331), .Y(div_n614) );
  INVX0_LVT div_U222 ( .A(div_n788), .Y(div_n605) );
  INVX0_LVT div_U221 ( .A(div_n777), .Y(div_n974) );
  INVX0_LVT div_U220 ( .A(div_n967), .Y(div_n216) );
  INVX0_LVT div_U219 ( .A(div_n966), .Y(div_n723) );
  INVX0_LVT div_U218 ( .A(div_n615), .Y(div_n312) );
  INVX0_LVT div_U217 ( .A(div_n1002), .Y(div_n972) );
  MUX21X1_LVT div_U216 ( .A1(n_T_702[31]), .A2(n_T_702[63]), .S0(alu_io_dw), 
        .Y(div_n324) );
  INVX0_LVT div_U215 ( .A(div_n956), .Y(div_n969) );
  NOR4X0_LVT div_U214 ( .A1(div_n974), .A2(div_n973), .A3(div_n997), .A4(
        div_n_T_430_5_), .Y(div_n1001) );
  NOR2X1_LVT div_U213 ( .A1(div_n_T_273_5_), .A2(div_n940), .Y(div_n763) );
  INVX0_LVT div_U212 ( .A(div_n338), .Y(div_n333) );
  INVX0_LVT div_U211 ( .A(div_n763), .Y(div_n968) );
  INVX0_LVT div_U210 ( .A(div_n957), .Y(div_n963) );
  NOR2X1_LVT div_U209 ( .A1(div_n320), .A2(div_io_kill), .Y(div_n753) );
  INVX0_LVT div_U208 ( .A(div_n753), .Y(div_n327) );
  INVX0_LVT div_U207 ( .A(div_subtractor_64_), .Y(div_n310) );
  INVX0_LVT div_U206 ( .A(div_n_T_434_3_), .Y(div_n168) );
  INVX0_LVT div_U205 ( .A(div_n_T_434_4_), .Y(div_n169) );
  INVX0_LVT div_U204 ( .A(div_n_T_434_5_), .Y(div_n170) );
  INVX1_LVT div_U203 ( .A(reset), .Y(div_n309) );
  INVX1_LVT div_U202 ( .A(alu_io_fn[2]), .Y(div_n784) );
  INVX1_LVT div_U201 ( .A(alu_io_dw), .Y(div_n787) );
  INVX1_LVT div_U200 ( .A(alu_io_fn[0]), .Y(div_n786) );
  INVX1_LVT div_U199 ( .A(alu_io_fn[1]), .Y(div_n785) );
  INVX1_LVT div_U198 ( .A(div_n1000), .Y(div_n744) );
  INVX1_LVT div_U197 ( .A(div_n655), .Y(div_n222) );
  NAND2X4_LVT div_U196 ( .A1(io_fpu_fromint_data[31]), .A2(div_n337), .Y(
        div_n658) );
  NAND2X4_LVT div_U195 ( .A1(div_n616), .A2(div_n615), .Y(div_n633) );
  HADDX1_LVT div_U194 ( .A0(div_n141), .B0(div_n155), .SO(div_n_T_97_6_) );
  NAND2X0_LVT div_U193 ( .A1(div_n_T_69_8_), .A2(div_n803), .Y(div_n141) );
  NAND3X0_LVT div_U192 ( .A1(div_n140), .A2(div_n633), .A3(div_n139), .Y(
        div_N382) );
  NAND2X0_LVT div_U191 ( .A1(div_subtractor_59_), .A2(div_n754), .Y(div_n140)
         );
  NAND2X0_LVT div_U190 ( .A1(div_n655), .A2(n_T_702[59]), .Y(div_n139) );
  NAND3X0_LVT div_U189 ( .A1(div_n137), .A2(div_n633), .A3(div_n138), .Y(
        div_N371) );
  NAND2X0_LVT div_U188 ( .A1(div_n655), .A2(n_T_702[48]), .Y(div_n138) );
  NAND2X0_LVT div_U187 ( .A1(div_subtractor_48_), .A2(div_n754), .Y(div_n137)
         );
  AO22X1_LVT div_U186 ( .A1(div_n224), .A2(div_negated_remainder[52]), .A3(
        div_n225), .A4(div_n_T_442[52]), .Y(div_n136) );
  AO22X1_LVT div_U184 ( .A1(div_n_T_51_60_), .A2(div_n223), .A3(
        io_fpu_fromint_data[52]), .A4(div_n655), .Y(div_n133) );
  INVX0_LVT div_U183 ( .A(div_n658), .Y(div_n132) );
  AND2X1_LVT div_U182 ( .A1(div_n781), .A2(div_n131), .Y(div_n745) );
  INVX0_LVT div_U181 ( .A(div_n1000), .Y(div_n131) );
  NAND3X0_LVT div_U180 ( .A1(div_n129), .A2(div_n633), .A3(div_n130), .Y(
        div_N379) );
  NAND2X0_LVT div_U179 ( .A1(div_n655), .A2(n_T_702[56]), .Y(div_n130) );
  NAND2X0_LVT div_U178 ( .A1(div_subtractor_56_), .A2(div_n754), .Y(div_n129)
         );
  NAND3X0_LVT div_U177 ( .A1(div_n127), .A2(div_n633), .A3(div_n128), .Y(
        div_N375) );
  NAND2X0_LVT div_U176 ( .A1(div_n655), .A2(n_T_702[52]), .Y(div_n128) );
  NAND2X0_LVT div_U175 ( .A1(div_subtractor_52_), .A2(div_n754), .Y(div_n127)
         );
  NAND3X0_LVT div_U174 ( .A1(div_n125), .A2(div_n633), .A3(div_n126), .Y(
        div_N358) );
  NAND2X0_LVT div_U173 ( .A1(div_n655), .A2(n_T_702[35]), .Y(div_n126) );
  NAND2X0_LVT div_U172 ( .A1(div_subtractor_35_), .A2(div_n754), .Y(div_n125)
         );
  AO22X1_LVT div_U171 ( .A1(div_n224), .A2(div_negated_remainder[32]), .A3(
        div_n225), .A4(div_n_T_442[32]), .Y(div_n124) );
  AO22X1_LVT div_U169 ( .A1(div_n_T_51_40_), .A2(div_n223), .A3(
        io_fpu_fromint_data[32]), .A4(div_n655), .Y(div_n121) );
  INVX0_LVT div_U168 ( .A(div_n658), .Y(div_n120) );
  AO22X1_LVT div_U166 ( .A1(div_n679), .A2(div_n_T_87[1]), .A3(div_n302), .A4(
        div_n227), .Y(div_n118) );
  AO222X1_LVT div_U165 ( .A1(div_n223), .A2(div_n_T_51_9_), .A3(div_n235), 
        .A4(io_fpu_fromint_data[1]), .A5(div_negated_remainder[1]), .A6(
        div_n224), .Y(div_n117) );
  NAND3X0_LVT div_U164 ( .A1(div_n115), .A2(div_n633), .A3(div_n116), .Y(
        div_N374) );
  NAND2X0_LVT div_U163 ( .A1(div_n655), .A2(n_T_702[51]), .Y(div_n116) );
  NAND2X0_LVT div_U162 ( .A1(div_subtractor_51_), .A2(div_n754), .Y(div_n115)
         );
  NAND3X0_LVT div_U161 ( .A1(div_n113), .A2(div_n633), .A3(div_n114), .Y(
        div_N367) );
  NAND2X0_LVT div_U160 ( .A1(div_n655), .A2(n_T_702[44]), .Y(div_n114) );
  NAND2X0_LVT div_U159 ( .A1(div_subtractor_44_), .A2(div_n754), .Y(div_n113)
         );
  NAND3X0_LVT div_U158 ( .A1(div_n111), .A2(div_n633), .A3(div_n112), .Y(
        div_N355) );
  NAND2X0_LVT div_U157 ( .A1(div_n655), .A2(n_T_702[32]), .Y(div_n112) );
  NAND2X0_LVT div_U156 ( .A1(div_subtractor_32_), .A2(div_n754), .Y(div_n111)
         );
  AND3X1_LVT div_U155 ( .A1(div_n342), .A2(div_n343), .A3(div_n110), .Y(
        div_n157) );
  INVX0_LVT div_U154 ( .A(div_n344), .Y(div_n110) );
  NAND3X0_LVT div_U153 ( .A1(div_n108), .A2(div_n207), .A3(div_n109), .Y(
        div_N394) );
  AOI22X1_LVT div_U152 ( .A1(div_n_T_87[0]), .A2(div_n679), .A3(div_n157), 
        .A4(div_n_T_442[0]), .Y(div_n109) );
  AOI222X1_LVT div_U151 ( .A1(div_n_T_51_8_), .A2(div_n223), .A3(div_n224), 
        .A4(div_result_0_), .A5(io_fpu_fromint_data[0]), .A6(div_n235), .Y(
        div_n108) );
  AO22X1_LVT div_U149 ( .A1(div_n679), .A2(div_n_T_87[4]), .A3(div_n305), .A4(
        div_n227), .Y(div_n106) );
  AO222X1_LVT div_U148 ( .A1(div_n_T_51_12_), .A2(div_n223), .A3(div_n224), 
        .A4(div_negated_remainder[4]), .A5(io_fpu_fromint_data[4]), .A6(
        div_n235), .Y(div_n105) );
  NAND3X0_LVT div_U147 ( .A1(div_n104), .A2(div_n633), .A3(div_n103), .Y(
        div_N385) );
  NAND2X0_LVT div_U146 ( .A1(div_subtractor_62_), .A2(div_n754), .Y(div_n104)
         );
  NAND2X0_LVT div_U145 ( .A1(div_n655), .A2(n_T_702[62]), .Y(div_n103) );
  NAND3X0_LVT div_U144 ( .A1(div_n101), .A2(div_n633), .A3(div_n102), .Y(
        div_N366) );
  NAND2X0_LVT div_U143 ( .A1(div_n655), .A2(n_T_702[43]), .Y(div_n102) );
  NAND2X0_LVT div_U142 ( .A1(div_subtractor_43_), .A2(div_n754), .Y(div_n101)
         );
  AO22X1_LVT div_U141 ( .A1(div_n209), .A2(div_result_11_), .A3(div_result_43_), .A4(div_n146), .Y(div_io_resp_bits_data[11]) );
  AO21X1_LVT div_U140 ( .A1(div_n_T_442[16]), .A2(div_n225), .A3(div_n100), 
        .Y(div_N410) );
  AO22X1_LVT div_U138 ( .A1(div_n679), .A2(div_n_T_87[16]), .A3(div_n224), 
        .A4(div_negated_remainder[16]), .Y(div_n98) );
  AO22X1_LVT div_U137 ( .A1(div_n_T_51_24_), .A2(div_n223), .A3(
        io_fpu_fromint_data[16]), .A4(div_n235), .Y(div_n97) );
  NAND3X0_LVT div_U136 ( .A1(div_n95), .A2(div_n633), .A3(div_n96), .Y(
        div_N384) );
  NAND2X0_LVT div_U135 ( .A1(div_n655), .A2(n_T_702[61]), .Y(div_n96) );
  NAND2X0_LVT div_U134 ( .A1(div_subtractor_61_), .A2(div_n754), .Y(div_n95)
         );
  AO22X1_LVT div_U132 ( .A1(div_n679), .A2(div_n_T_87[2]), .A3(div_n_T_51_1_), 
        .A4(div_n227), .Y(div_n93) );
  AO222X1_LVT div_U131 ( .A1(div_n90), .A2(div_n91), .A3(
        div_negated_remainder[2]), .A4(div_n224), .A5(div_n235), .A6(
        io_fpu_fromint_data[2]), .Y(div_n92) );
  INVX0_LVT div_U130 ( .A(div_n201), .Y(div_n91) );
  INVX0_LVT div_U129 ( .A(div_n286), .Y(div_n90) );
  AO22X1_LVT div_U127 ( .A1(div_n224), .A2(div_negated_remainder[24]), .A3(
        div_n_T_51_23_), .A4(div_n227), .Y(div_n88) );
  AO222X1_LVT div_U126 ( .A1(div_n_T_51_32_), .A2(div_n223), .A3(div_n679), 
        .A4(div_n_T_87[24]), .A5(io_fpu_fromint_data[24]), .A6(div_n235), .Y(
        div_n87) );
  NAND3X0_LVT div_U125 ( .A1(div_n85), .A2(div_n633), .A3(div_n86), .Y(
        div_N383) );
  NAND2X0_LVT div_U124 ( .A1(div_n655), .A2(n_T_702[60]), .Y(div_n86) );
  NAND2X0_LVT div_U123 ( .A1(div_subtractor_60_), .A2(div_n754), .Y(div_n85)
         );
  NAND3X0_LVT div_U121 ( .A1(div_n82), .A2(div_n633), .A3(div_n83), .Y(
        div_N386) );
  NAND2X0_LVT div_U120 ( .A1(div_n655), .A2(n_T_702[63]), .Y(div_n83) );
  NAND2X0_LVT div_U119 ( .A1(div_subtractor_63_), .A2(div_n754), .Y(div_n82)
         );
  AO22X1_LVT div_U118 ( .A1(div_n224), .A2(div_negated_remainder[40]), .A3(
        div_n225), .A4(div_n_T_442[40]), .Y(div_n81) );
  AO22X1_LVT div_U116 ( .A1(div_n_T_51_48_), .A2(div_n223), .A3(
        io_fpu_fromint_data[40]), .A4(div_n655), .Y(div_n78) );
  INVX0_LVT div_U115 ( .A(div_n658), .Y(div_n77) );
  AO222X1_LVT div_U114 ( .A1(div_n783), .A2(div_n76), .A3(div_n157), .A4(
        div_n_T_442[64]), .A5(div_n227), .A6(div_n_T_51_63_), .Y(div_N458) );
  AND3X1_LVT div_U113 ( .A1(div_n204), .A2(div_neg_out), .A3(div_n75), .Y(
        div_n76) );
  AND4X1_LVT div_U112 ( .A1(div_n_T_69_4_), .A2(div_n613), .A3(div_n_T_71_39_), 
        .A4(div_n614), .Y(div_n75) );
  AO22X1_LVT div_U110 ( .A1(div_n224), .A2(div_negated_remainder[12]), .A3(
        div_n_T_51_11_), .A4(div_n227), .Y(div_n73) );
  AO222X1_LVT div_U109 ( .A1(div_n_T_51_20_), .A2(div_n223), .A3(div_n679), 
        .A4(div_n_T_87[12]), .A5(io_fpu_fromint_data[12]), .A6(div_n235), .Y(
        div_n72) );
  NAND3X0_LVT div_U108 ( .A1(div_n70), .A2(div_n633), .A3(div_n71), .Y(
        div_N380) );
  NAND2X0_LVT div_U107 ( .A1(div_n655), .A2(n_T_702[57]), .Y(div_n71) );
  NAND2X0_LVT div_U106 ( .A1(div_subtractor_57_), .A2(div_n754), .Y(div_n70)
         );
  AO22X1_LVT div_U105 ( .A1(div_n224), .A2(div_negated_remainder[48]), .A3(
        div_n225), .A4(div_n_T_442[48]), .Y(div_n69) );
  AO22X1_LVT div_U103 ( .A1(div_n_T_51_56_), .A2(div_n223), .A3(
        io_fpu_fromint_data[48]), .A4(div_n655), .Y(div_n66) );
  INVX0_LVT div_U102 ( .A(div_n658), .Y(div_n65) );
  AO22X1_LVT div_U101 ( .A1(div_n209), .A2(div_result_22_), .A3(div_result_54_), .A4(div_n146), .Y(div_io_resp_bits_data[22]) );
  NAND2X0_LVT div_U100 ( .A1(div_n343), .A2(div_n64), .Y(div_n207) );
  INVX0_LVT div_U99 ( .A(div_subtractor_64_), .Y(div_n64) );
  NAND3X0_LVT div_U98 ( .A1(div_n62), .A2(div_n633), .A3(div_n63), .Y(div_N372) );
  NAND2X0_LVT div_U97 ( .A1(div_n655), .A2(n_T_702[49]), .Y(div_n63) );
  NAND2X0_LVT div_U96 ( .A1(div_subtractor_49_), .A2(div_n754), .Y(div_n62) );
  NAND4X0_LVT div_U95 ( .A1(div_n790), .A2(div_n980), .A3(div_n60), .A4(
        div_n61), .Y(div_n338) );
  NAND2X0_LVT div_U94 ( .A1(div_n1000), .A2(div_n800), .Y(div_n61) );
  AND4X1_LVT div_U93 ( .A1(div_n51), .A2(div_n54), .A3(div_n56), .A4(div_n59), 
        .Y(div_n60) );
  NAND2X0_LVT div_U92 ( .A1(div_n210), .A2(div_n58), .Y(div_n59) );
  NAND3X0_LVT div_U90 ( .A1(div_n55), .A2(div_n148), .A3(div_n210), .Y(div_n56) );
  NAND2X0_LVT div_U89 ( .A1(div_n732), .A2(div_n779), .Y(div_n55) );
  AND4X1_LVT div_U88 ( .A1(div_n781), .A2(div_n189), .A3(div_n296), .A4(
        div_n53), .Y(div_n54) );
  NOR4X0_LVT div_U87 ( .A1(div_n302), .A2(div_n305), .A3(div_n304), .A4(
        div_n52), .Y(div_n53) );
  OA22X1_LVT div_U86 ( .A1(div_n148), .A2(div_n210), .A3(div_n973), .A4(
        div_n974), .Y(div_n52) );
  OA22X1_LVT div_U85 ( .A1(div_n773), .A2(div_n789), .A3(div_n775), .A4(
        div_n788), .Y(div_n51) );
  NAND3X0_LVT div_U84 ( .A1(div_n49), .A2(div_n633), .A3(div_n50), .Y(div_N381) );
  NAND2X0_LVT div_U83 ( .A1(div_n655), .A2(n_T_702[58]), .Y(div_n50) );
  NAND2X0_LVT div_U82 ( .A1(div_subtractor_58_), .A2(div_n754), .Y(div_n49) );
  AO22X1_LVT div_U81 ( .A1(div_n_T_51_55_), .A2(div_n227), .A3(div_n225), .A4(
        div_n_T_442[56]), .Y(div_n48) );
  AO22X1_LVT div_U79 ( .A1(div_n_T_65[0]), .A2(div_n223), .A3(
        io_fpu_fromint_data[56]), .A4(div_n655), .Y(div_n45) );
  INVX0_LVT div_U78 ( .A(div_n658), .Y(div_n44) );
  AND2X1_LVT div_U77 ( .A1(div_n246), .A2(div_n43), .Y(div_n756) );
  AOI222X1_LVT div_U76 ( .A1(div_n_T_51_39_), .A2(div_n741), .A3(
        div_n_T_51_35_), .A4(div_n742), .A5(div_n_T_51_43_), .A6(div_n771), 
        .Y(div_n43) );
  NAND3X0_LVT div_U74 ( .A1(div_n40), .A2(div_n633), .A3(div_n41), .Y(div_N378) );
  NAND2X0_LVT div_U73 ( .A1(div_n655), .A2(n_T_702[55]), .Y(div_n41) );
  NAND2X0_LVT div_U72 ( .A1(div_subtractor_55_), .A2(div_n754), .Y(div_n40) );
  NAND3X0_LVT div_U71 ( .A1(div_n38), .A2(div_n633), .A3(div_n39), .Y(div_N364) );
  NAND2X0_LVT div_U70 ( .A1(div_n655), .A2(n_T_702[41]), .Y(div_n39) );
  NAND2X0_LVT div_U69 ( .A1(div_subtractor_41_), .A2(div_n754), .Y(div_n38) );
  NAND3X0_LVT div_U68 ( .A1(div_n36), .A2(div_n633), .A3(div_n37), .Y(div_N376) );
  NAND2X0_LVT div_U67 ( .A1(div_n655), .A2(n_T_702[53]), .Y(div_n37) );
  NAND2X0_LVT div_U66 ( .A1(div_subtractor_53_), .A2(div_n754), .Y(div_n36) );
  NAND3X0_LVT div_U65 ( .A1(div_n774), .A2(div_n33), .A3(div_n35), .Y(
        div_n_T_429[2]) );
  AO21X1_LVT div_U64 ( .A1(div_n771), .A2(div_n34), .A3(div_n972), .Y(div_n35)
         );
  NAND2X0_LVT div_U63 ( .A1(div_n971), .A2(div_n772), .Y(div_n34) );
  OA22X1_LVT div_U62 ( .A1(div_n_T_430_5_), .A2(div_n31), .A3(div_n779), .A4(
        div_n32), .Y(div_n33) );
  INVX0_LVT div_U61 ( .A(div_n773), .Y(div_n32) );
  OA21X1_LVT div_U60 ( .A1(div_n1000), .A2(div_n781), .A3(div_n780), .Y(
        div_n30) );
  AND2X1_LVT div_U59 ( .A1(div_n309), .A2(alu_io_fn[2]), .Y(div_n29) );
  NAND3X0_LVT div_U58 ( .A1(div_n27), .A2(div_n633), .A3(div_n28), .Y(div_N377) );
  NAND2X0_LVT div_U57 ( .A1(div_n655), .A2(n_T_702[54]), .Y(div_n28) );
  NAND2X0_LVT div_U56 ( .A1(div_subtractor_54_), .A2(div_n754), .Y(div_n27) );
  AND2X1_LVT div_U55 ( .A1(div_n149), .A2(div_n26), .Y(div_n758) );
  AOI222X1_LVT div_U54 ( .A1(div_n_T_51_51_), .A2(div_n747), .A3(
        div_n_T_51_55_), .A4(div_n773), .A5(div_n_T_51_59_), .A6(div_n774), 
        .Y(div_n26) );
  NAND3X0_LVT div_U53 ( .A1(div_n24), .A2(div_n633), .A3(div_n25), .Y(div_N370) );
  NAND2X0_LVT div_U52 ( .A1(div_n655), .A2(n_T_702[47]), .Y(div_n25) );
  NAND2X0_LVT div_U51 ( .A1(div_subtractor_47_), .A2(div_n754), .Y(div_n24) );
  AO22X1_LVT div_U49 ( .A1(div_n1002), .A2(div_n18), .A3(div_n1001), .A4(
        div_n21), .Y(div_n22) );
  NAND4X0_LVT div_U48 ( .A1(div_n282), .A2(div_n757), .A3(div_n19), .A4(
        div_n20), .Y(div_n21) );
  OR2X1_LVT div_U47 ( .A1(div_n286), .A2(div_n743), .Y(div_n20) );
  AOI22X1_LVT div_U46 ( .A1(div_n304), .A2(div_n745), .A3(div_n_T_51_6_), .A4(
        div_n744), .Y(div_n19) );
  NAND4X0_LVT div_U45 ( .A1(div_n247), .A2(div_n756), .A3(div_n16), .A4(
        div_n17), .Y(div_n18) );
  OR2X1_LVT div_U44 ( .A1(div_n251), .A2(div_n740), .Y(div_n17) );
  AOI22X1_LVT div_U43 ( .A1(div_n_T_51_34_), .A2(div_n742), .A3(div_n_T_51_38_), .A4(div_n741), .Y(div_n16) );
  NAND4X0_LVT div_U42 ( .A1(div_n264), .A2(div_n755), .A3(div_n13), .A4(
        div_n14), .Y(div_n15) );
  OR2X1_LVT div_U41 ( .A1(div_n268), .A2(div_n748), .Y(div_n14) );
  AOI22X1_LVT div_U40 ( .A1(div_n775), .A2(div_n_T_51_22_), .A3(div_n_T_51_18_), .A4(div_n749), .Y(div_n13) );
  NAND4X0_LVT div_U39 ( .A1(div_n9), .A2(div_n758), .A3(div_n10), .A4(div_n11), 
        .Y(div_n12) );
  NAND2X0_LVT div_U38 ( .A1(div_n747), .A2(div_n_T_51_50_), .Y(div_n11) );
  NAND2X0_LVT div_U37 ( .A1(div_n773), .A2(div_n_T_51_54_), .Y(div_n10) );
  OA21X1_LVT div_U36 ( .A1(div_n232), .A2(div_n746), .A3(div_n228), .Y(div_n9)
         );
  NAND3X0_LVT div_U35 ( .A1(div_n7), .A2(div_n633), .A3(div_n8), .Y(div_N373)
         );
  NAND2X0_LVT div_U34 ( .A1(div_n655), .A2(n_T_702[50]), .Y(div_n8) );
  NAND2X0_LVT div_U33 ( .A1(div_subtractor_50_), .A2(div_n754), .Y(div_n7) );
  NAND3X0_LVT div_U32 ( .A1(div_n5), .A2(div_n633), .A3(div_n6), .Y(div_N363)
         );
  NAND2X0_LVT div_U31 ( .A1(div_n655), .A2(n_T_702[40]), .Y(div_n6) );
  NAND2X0_LVT div_U30 ( .A1(div_subtractor_40_), .A2(div_n754), .Y(div_n5) );
  NAND3X0_LVT div_U29 ( .A1(div_n3), .A2(div_n633), .A3(div_n4), .Y(div_N369)
         );
  NAND2X0_LVT div_U28 ( .A1(div_n655), .A2(n_T_702[46]), .Y(div_n4) );
  NAND2X0_LVT div_U27 ( .A1(div_subtractor_46_), .A2(div_n754), .Y(div_n3) );
  AND2X1_LVT div_U26 ( .A1(div_n263), .A2(div_n2), .Y(div_n755) );
  AOI222X1_LVT div_U25 ( .A1(div_n_T_51_23_), .A2(div_n775), .A3(div_n749), 
        .A4(div_n_T_51_19_), .A5(div_n_T_51_27_), .A6(div_n776), .Y(div_n2) );
  INVX1_LVT div_U24 ( .A(div_n209), .Y(div_n146) );
  OA221X1_LVT div_U23 ( .A1(div_n975), .A2(div_n30), .A3(div_n777), .A4(
        div_n997), .A5(div_n776), .Y(div_n31) );
  AO221X1_LVT div_U22 ( .A1(1'b1), .A2(div_n12), .A3(div_n1003), .A4(div_n15), 
        .A5(div_n22), .Y(div_n_T_429[1]) );
  AO222X1_LVT div_U21 ( .A1(div_n753), .A2(div_n224), .A3(div_n680), .A4(1'b1), 
        .A5(div_n29), .A6(div_n235), .Y(div_N283) );
  AO221X1_LVT div_U20 ( .A1(1'b1), .A2(div_n47), .A3(div_n224), .A4(
        div_negated_remainder[56]), .A5(div_n48), .Y(div_N450) );
  AO221X1_LVT div_U19 ( .A1(1'b1), .A2(div_n44), .A3(div_n_T_87[56]), .A4(
        div_n679), .A5(div_n45), .Y(div_n47) );
  AO221X1_LVT div_U18 ( .A1(1'b1), .A2(div_n971), .A3(div_n999), .A4(div_n795), 
        .A5(div_n970), .Y(div_n58) );
  AO221X1_LVT div_U17 ( .A1(1'b1), .A2(div_n68), .A3(div_n_T_51_47_), .A4(
        div_n227), .A5(div_n69), .Y(div_N442) );
  AO221X1_LVT div_U16 ( .A1(1'b1), .A2(div_n65), .A3(div_n_T_87[48]), .A4(
        div_n679), .A5(div_n66), .Y(div_n68) );
  AO221X1_LVT div_U15 ( .A1(1'b1), .A2(div_n72), .A3(div_n225), .A4(
        div_n_T_442[12]), .A5(div_n73), .Y(div_N406) );
  AO221X1_LVT div_U14 ( .A1(1'b1), .A2(div_n80), .A3(div_n_T_51_39_), .A4(
        div_n227), .A5(div_n81), .Y(div_N434) );
  AO221X1_LVT div_U13 ( .A1(1'b1), .A2(div_n77), .A3(div_n_T_87[40]), .A4(
        div_n679), .A5(div_n78), .Y(div_n80) );
  AO221X1_LVT div_U12 ( .A1(1'b1), .A2(div_n977), .A3(div_n_T_51_63_), .A4(
        div_n224), .A5(div_N293), .Y(div_N493) );
  AO221X1_LVT div_U11 ( .A1(1'b1), .A2(div_n87), .A3(div_n157), .A4(
        div_n_T_442[24]), .A5(div_n88), .Y(div_N418) );
  AO221X1_LVT div_U10 ( .A1(1'b1), .A2(div_n92), .A3(div_n225), .A4(
        div_n_T_442[2]), .A5(div_n93), .Y(div_N396) );
  AO221X1_LVT div_U9 ( .A1(1'b1), .A2(div_n97), .A3(div_n227), .A4(
        div_n_T_51_15_), .A5(div_n98), .Y(div_n100) );
  AO221X1_LVT div_U8 ( .A1(1'b1), .A2(div_n105), .A3(div_n225), .A4(
        div_n_T_442[4]), .A5(div_n106), .Y(div_N398) );
  AO221X1_LVT div_U7 ( .A1(1'b1), .A2(div_n117), .A3(div_n225), .A4(
        div_n_T_442[1]), .A5(div_n118), .Y(div_N395) );
  AO221X1_LVT div_U6 ( .A1(1'b1), .A2(div_n123), .A3(div_n_T_51_31_), .A4(
        div_n227), .A5(div_n124), .Y(div_N426) );
  AO221X1_LVT div_U5 ( .A1(1'b1), .A2(div_n120), .A3(div_n_T_87[32]), .A4(
        div_n679), .A5(div_n121), .Y(div_n123) );
  AO221X1_LVT div_U4 ( .A1(1'b1), .A2(div_n135), .A3(div_n_T_51_51_), .A4(
        div_n227), .A5(div_n136), .Y(div_N446) );
  AO221X1_LVT div_U3 ( .A1(1'b1), .A2(div_n132), .A3(div_n_T_87[52]), .A4(
        div_n679), .A5(div_n133), .Y(div_n135) );
  DFFX1_LVT div_isHi_reg ( .D(div_n145), .CLK(div_net34690), .Q(div_n189), 
        .QN(div_isHi) );
  OA21X1_LVT div_isHi_reg_U2 ( .A1(alu_io_fn[2]), .A2(div_n786), .A3(div_n785), 
        .Y(div_n145) );
  DFFX1_LVT div_count_reg_0_ ( .D(div_N294), .CLK(div_net34695), .Q(div_n300), 
        .QN(div_n204) );
  DFFX1_LVT div_resHi_reg ( .D(div_n794), .CLK(div_net34700), .Q(div_resHi) );
  DFFSSRX1_LVT div_remainder_reg_129_ ( .D(div_n230), .SETB(div_n_T_65[72]), 
        .RSTB(1'b1), .CLK(div_n245), .QN(div_n_T_51_128_) );
  DFFX1_LVT div_remainder_reg_128_ ( .D(div_N523), .CLK(div_n245), .Q(
        div_n_T_51_127_) );
  DFFX1_LVT div_remainder_reg_127_ ( .D(div_N522), .CLK(div_n245), .Q(
        div_n_T_51_126_) );
  DFFX1_LVT div_remainder_reg_126_ ( .D(div_N521), .CLK(div_n245), .Q(
        div_n_T_51_125_) );
  DFFX1_LVT div_remainder_reg_125_ ( .D(div_N520), .CLK(div_n245), .Q(
        div_n_T_51_124_) );
  DFFX1_LVT div_remainder_reg_124_ ( .D(div_N519), .CLK(div_n245), .Q(
        div_n_T_51_123_) );
  DFFX1_LVT div_remainder_reg_123_ ( .D(div_N518), .CLK(div_n245), .Q(
        div_n_T_51_122_) );
  DFFX1_LVT div_remainder_reg_122_ ( .D(div_N517), .CLK(div_n245), .Q(
        div_n_T_51_121_) );
  DFFX1_LVT div_remainder_reg_121_ ( .D(div_N516), .CLK(div_n245), .Q(
        div_n_T_51_120_) );
  DFFX1_LVT div_remainder_reg_120_ ( .D(div_N515), .CLK(div_n245), .Q(
        div_n_T_51_119_) );
  DFFX1_LVT div_remainder_reg_119_ ( .D(div_N514), .CLK(div_n245), .Q(
        div_n_T_51_118_) );
  DFFX1_LVT div_remainder_reg_118_ ( .D(div_N513), .CLK(div_n245), .Q(
        div_n_T_51_117_) );
  DFFX1_LVT div_remainder_reg_117_ ( .D(div_N512), .CLK(div_n253), .Q(
        div_n_T_51_116_) );
  DFFX1_LVT div_remainder_reg_116_ ( .D(div_N511), .CLK(div_n253), .Q(
        div_n_T_51_115_) );
  DFFX1_LVT div_remainder_reg_115_ ( .D(div_N510), .CLK(div_n253), .Q(
        div_n_T_51_114_) );
  DFFX1_LVT div_remainder_reg_114_ ( .D(div_N509), .CLK(div_n253), .Q(
        div_n_T_51_113_) );
  DFFX1_LVT div_remainder_reg_113_ ( .D(div_N508), .CLK(div_n253), .Q(
        div_n_T_51_112_) );
  DFFX1_LVT div_remainder_reg_112_ ( .D(div_N507), .CLK(div_n253), .Q(
        div_n_T_51_111_) );
  DFFX1_LVT div_remainder_reg_111_ ( .D(div_N506), .CLK(div_n253), .Q(
        div_n_T_51_110_) );
  DFFX1_LVT div_remainder_reg_110_ ( .D(div_N505), .CLK(div_n253), .Q(
        div_n_T_51_109_) );
  DFFX1_LVT div_remainder_reg_109_ ( .D(div_N504), .CLK(div_n253), .Q(
        div_n_T_51_108_) );
  DFFX1_LVT div_remainder_reg_108_ ( .D(div_N503), .CLK(div_n253), .Q(
        div_n_T_51_107_) );
  DFFX1_LVT div_remainder_reg_107_ ( .D(div_N502), .CLK(div_n253), .Q(
        div_n_T_51_106_) );
  DFFX1_LVT div_remainder_reg_106_ ( .D(div_N501), .CLK(div_n253), .Q(
        div_n_T_51_105_) );
  DFFX1_LVT div_remainder_reg_105_ ( .D(div_N500), .CLK(div_n262), .Q(
        div_n_T_51_104_) );
  DFFX1_LVT div_remainder_reg_104_ ( .D(div_N499), .CLK(div_n262), .Q(
        div_n_T_51_103_) );
  DFFX1_LVT div_remainder_reg_103_ ( .D(div_N498), .CLK(div_n262), .Q(
        div_n_T_51_102_) );
  DFFX1_LVT div_remainder_reg_102_ ( .D(div_N497), .CLK(div_n262), .Q(
        div_n_T_51_101_) );
  DFFX1_LVT div_remainder_reg_101_ ( .D(div_N496), .CLK(div_n262), .Q(
        div_n_T_51_100_) );
  DFFX1_LVT div_remainder_reg_100_ ( .D(div_N495), .CLK(div_n262), .Q(
        div_n_T_51_99_) );
  DFFX1_LVT div_remainder_reg_99_ ( .D(div_N494), .CLK(div_n262), .Q(
        div_n_T_51_98_) );
  DFFX1_LVT div_remainder_reg_98_ ( .D(div_N492), .CLK(div_n262), .Q(
        div_n_T_51_97_) );
  DFFX1_LVT div_remainder_reg_97_ ( .D(div_N491), .CLK(div_n262), .Q(
        div_n_T_51_96_) );
  DFFX1_LVT div_remainder_reg_96_ ( .D(div_N490), .CLK(div_n262), .Q(
        div_n_T_51_95_) );
  DFFX1_LVT div_remainder_reg_95_ ( .D(div_N489), .CLK(div_n262), .Q(
        div_n_T_51_94_) );
  DFFX1_LVT div_remainder_reg_94_ ( .D(div_N488), .CLK(div_n262), .Q(
        div_n_T_51_93_) );
  DFFX1_LVT div_remainder_reg_93_ ( .D(div_N487), .CLK(div_n265), .Q(
        div_n_T_51_92_) );
  DFFX1_LVT div_remainder_reg_92_ ( .D(div_N486), .CLK(div_n265), .Q(
        div_n_T_51_91_) );
  DFFX1_LVT div_remainder_reg_91_ ( .D(div_N485), .CLK(div_n265), .Q(
        div_n_T_51_90_) );
  DFFX1_LVT div_remainder_reg_90_ ( .D(div_N484), .CLK(div_n265), .Q(
        div_n_T_51_89_) );
  DFFX1_LVT div_remainder_reg_89_ ( .D(div_N483), .CLK(div_n265), .Q(
        div_n_T_51_88_) );
  DFFX1_LVT div_remainder_reg_88_ ( .D(div_N482), .CLK(div_n265), .Q(
        div_n_T_51_87_) );
  DFFX1_LVT div_remainder_reg_87_ ( .D(div_N481), .CLK(div_n265), .Q(
        div_n_T_51_86_) );
  DFFX1_LVT div_remainder_reg_86_ ( .D(div_N480), .CLK(div_n265), .Q(
        div_n_T_51_85_) );
  DFFX1_LVT div_remainder_reg_85_ ( .D(div_N479), .CLK(div_n265), .Q(
        div_n_T_51_84_) );
  DFFX1_LVT div_remainder_reg_84_ ( .D(div_N478), .CLK(div_n265), .Q(
        div_n_T_51_83_) );
  DFFX1_LVT div_remainder_reg_83_ ( .D(div_N477), .CLK(div_n265), .Q(
        div_n_T_51_82_) );
  DFFX1_LVT div_remainder_reg_82_ ( .D(div_N476), .CLK(div_n265), .Q(
        div_n_T_51_81_) );
  DFFX1_LVT div_remainder_reg_81_ ( .D(div_N475), .CLK(div_n271), .Q(
        div_n_T_51_80_) );
  DFFX1_LVT div_remainder_reg_80_ ( .D(div_N474), .CLK(div_n271), .Q(
        div_n_T_51_79_) );
  DFFX1_LVT div_remainder_reg_79_ ( .D(div_N473), .CLK(div_n271), .Q(
        div_n_T_51_78_) );
  DFFX1_LVT div_remainder_reg_78_ ( .D(div_N472), .CLK(div_n271), .Q(
        div_n_T_51_77_) );
  DFFX1_LVT div_remainder_reg_77_ ( .D(div_N471), .CLK(div_n271), .Q(
        div_n_T_51_76_) );
  DFFX1_LVT div_remainder_reg_76_ ( .D(div_N470), .CLK(div_n271), .Q(
        div_n_T_51_75_) );
  DFFX1_LVT div_remainder_reg_75_ ( .D(div_N469), .CLK(div_n271), .Q(
        div_n_T_51_74_) );
  DFFX1_LVT div_remainder_reg_74_ ( .D(div_N468), .CLK(div_n271), .Q(
        div_n_T_51_73_) );
  DFFX1_LVT div_remainder_reg_73_ ( .D(div_N467), .CLK(div_n271), .Q(
        div_n_T_51_72_) );
  DFFX1_LVT div_remainder_reg_72_ ( .D(div_N466), .CLK(div_n271), .Q(
        div_n_T_51_71_) );
  DFFX1_LVT div_remainder_reg_71_ ( .D(div_N465), .CLK(div_n271), .Q(
        div_n_T_51_70_) );
  DFFX1_LVT div_remainder_reg_70_ ( .D(div_N464), .CLK(div_n271), .Q(
        div_n_T_51_69_) );
  DFFX1_LVT div_remainder_reg_69_ ( .D(div_N463), .CLK(div_n276), .Q(
        div_n_T_51_68_) );
  DFFX1_LVT div_remainder_reg_68_ ( .D(div_N462), .CLK(div_n276), .Q(
        div_n_T_51_67_) );
  DFFX1_LVT div_remainder_reg_67_ ( .D(div_N461), .CLK(div_n276), .Q(
        div_n_T_51_66_) );
  DFFX1_LVT div_remainder_reg_66_ ( .D(div_N460), .CLK(div_n276), .Q(
        div_n_T_51_65_) );
  DFFX1_LVT div_remainder_reg_65_ ( .D(div_N459), .CLK(div_n276), .Q(
        div_n_T_51_64_) );
  DFFX1_LVT div_remainder_reg_64_ ( .D(div_N458), .CLK(div_n276), .Q(
        div_n_T_59_8_) );
  DFFX1_LVT div_remainder_reg_63_ ( .D(div_N457), .CLK(div_n276), .Q(
        div_n_T_51_63_), .QN(div_n149) );
  DFFX1_LVT div_remainder_reg_62_ ( .D(div_N456), .CLK(div_n276), .Q(
        div_n_T_51_62_), .QN(div_n228) );
  DFFX1_LVT div_remainder_reg_61_ ( .D(div_N455), .CLK(div_n276), .Q(
        div_n_T_51_61_), .QN(div_n229) );
  DFFX1_LVT div_remainder_reg_60_ ( .D(div_N454), .CLK(div_n276), .Q(
        div_n_T_51_60_), .QN(div_n187) );
  DFFX1_LVT div_remainder_reg_59_ ( .D(div_N453), .CLK(div_n276), .Q(
        div_n_T_51_59_), .QN(div_n231) );
  DFFX1_LVT div_remainder_reg_58_ ( .D(div_N452), .CLK(div_n276), .Q(
        div_n_T_51_58_), .QN(div_n232) );
  DFFX1_LVT div_remainder_reg_57_ ( .D(div_N451), .CLK(div_n279), .Q(
        div_n_T_51_57_), .QN(div_n233) );
  DFFX1_LVT div_remainder_reg_56_ ( .D(div_N450), .CLK(div_n279), .Q(
        div_n_T_51_56_), .QN(div_n234) );
  DFFX1_LVT div_remainder_reg_55_ ( .D(div_N449), .CLK(div_n279), .Q(
        div_n_T_51_55_), .QN(div_n236) );
  DFFX1_LVT div_remainder_reg_54_ ( .D(div_N448), .CLK(div_n279), .Q(
        div_n_T_51_54_), .QN(div_n237) );
  DFFX1_LVT div_remainder_reg_53_ ( .D(div_N447), .CLK(div_n279), .Q(
        div_n_T_51_53_), .QN(div_n238) );
  DFFX1_LVT div_remainder_reg_52_ ( .D(div_N446), .CLK(div_n279), .Q(
        div_n_T_51_52_), .QN(div_n239) );
  DFFX1_LVT div_remainder_reg_51_ ( .D(div_N445), .CLK(div_n279), .Q(
        div_n_T_51_51_), .QN(div_n240) );
  DFFX1_LVT div_remainder_reg_50_ ( .D(div_N444), .CLK(div_n279), .Q(
        div_n_T_51_50_), .QN(div_n241) );
  DFFX1_LVT div_remainder_reg_49_ ( .D(div_N443), .CLK(div_n279), .Q(
        div_n_T_51_49_), .QN(div_n182) );
  DFFX1_LVT div_remainder_reg_48_ ( .D(div_N442), .CLK(div_n279), .Q(
        div_n_T_51_48_), .QN(div_n243) );
  DFFX1_LVT div_remainder_reg_47_ ( .D(div_N441), .CLK(div_n279), .Q(
        div_n_T_51_47_), .QN(div_n246) );
  DFFX1_LVT div_remainder_reg_46_ ( .D(div_N440), .CLK(div_n279), .Q(
        div_n_T_51_46_), .QN(div_n247) );
  DFFX1_LVT div_remainder_reg_45_ ( .D(div_N439), .CLK(div_n280), .Q(
        div_n_T_51_45_), .QN(div_n248) );
  DFFX1_LVT div_remainder_reg_44_ ( .D(div_N438), .CLK(div_n280), .Q(
        div_n_T_51_44_), .QN(div_n249) );
  DFFX1_LVT div_remainder_reg_43_ ( .D(div_N437), .CLK(div_n280), .Q(
        div_n_T_51_43_), .QN(div_n250) );
  DFFX1_LVT div_remainder_reg_42_ ( .D(div_N436), .CLK(div_n280), .Q(
        div_n_T_51_42_), .QN(div_n251) );
  DFFX1_LVT div_remainder_reg_41_ ( .D(div_N435), .CLK(div_n280), .Q(
        div_n_T_51_41_), .QN(div_n252) );
  DFFX1_LVT div_remainder_reg_40_ ( .D(div_N434), .CLK(div_n280), .Q(
        div_n_T_51_40_), .QN(div_n188) );
  DFFX1_LVT div_remainder_reg_39_ ( .D(div_N433), .CLK(div_n280), .Q(
        div_n_T_51_39_), .QN(div_n254) );
  DFFX1_LVT div_remainder_reg_38_ ( .D(div_N432), .CLK(div_n280), .Q(
        div_n_T_51_38_), .QN(div_n255) );
  DFFX1_LVT div_remainder_reg_37_ ( .D(div_N431), .CLK(div_n280), .Q(
        div_n_T_51_37_), .QN(div_n256) );
  DFFX1_LVT div_remainder_reg_36_ ( .D(div_N430), .CLK(div_n280), .Q(
        div_n_T_51_36_), .QN(div_n257) );
  DFFX1_LVT div_remainder_reg_35_ ( .D(div_N429), .CLK(div_n280), .Q(
        div_n_T_51_35_), .QN(div_n258) );
  DFFX1_LVT div_remainder_reg_34_ ( .D(div_N428), .CLK(div_n280), .Q(
        div_n_T_51_34_), .QN(div_n259) );
  DFFX1_LVT div_remainder_reg_33_ ( .D(div_N427), .CLK(div_n285), .Q(
        div_n_T_51_33_), .QN(div_n260) );
  DFFX1_LVT div_remainder_reg_32_ ( .D(div_N426), .CLK(div_n285), .Q(
        div_n_T_51_32_), .QN(div_n261) );
  DFFX1_LVT div_divisor_reg_0_ ( .D(div_N323), .CLK(div_n289), .Q(
        div_divisor_0_) );
  DFFX1_LVT div_divisor_reg_1_ ( .D(div_N324), .CLK(div_n289), .Q(
        div_divisor_1_) );
  DFFX1_LVT div_divisor_reg_2_ ( .D(div_N325), .CLK(div_n289), .Q(
        div_divisor_2_), .QN(div_n205) );
  DFFX1_LVT div_divisor_reg_3_ ( .D(div_N326), .CLK(div_n289), .Q(
        div_divisor_3_) );
  DFFX1_LVT div_divisor_reg_4_ ( .D(div_N327), .CLK(div_n289), .Q(
        div_divisor_4_) );
  DFFX1_LVT div_divisor_reg_5_ ( .D(div_N328), .CLK(div_n289), .Q(
        div_divisor_5_) );
  DFFX1_LVT div_divisor_reg_6_ ( .D(div_N329), .CLK(div_n289), .Q(
        div_divisor_6_), .QN(div_n191) );
  DFFX1_LVT div_divisor_reg_7_ ( .D(div_N330), .CLK(div_n289), .Q(
        div_divisor_7_) );
  DFFX1_LVT div_divisor_reg_8_ ( .D(div_N331), .CLK(div_n289), .Q(
        div_divisor_8_), .QN(div_n165) );
  DFFX1_LVT div_divisor_reg_9_ ( .D(div_N332), .CLK(div_n289), .Q(
        div_divisor_9_) );
  DFFX1_LVT div_divisor_reg_10_ ( .D(div_N333), .CLK(div_n289), .Q(
        div_divisor_10_), .QN(div_n202) );
  DFFX1_LVT div_divisor_reg_11_ ( .D(div_N334), .CLK(div_n289), .Q(
        div_divisor_11_) );
  DFFX1_LVT div_divisor_reg_12_ ( .D(div_N335), .CLK(div_n294), .Q(
        div_divisor_12_) );
  DFFX1_LVT div_divisor_reg_13_ ( .D(div_N336), .CLK(div_n294), .Q(
        div_divisor_13_), .QN(div_n172) );
  DFFX1_LVT div_divisor_reg_14_ ( .D(div_N337), .CLK(div_n294), .Q(
        div_divisor_14_), .QN(div_n193) );
  DFFX1_LVT div_divisor_reg_15_ ( .D(div_N338), .CLK(div_n294), .Q(
        div_divisor_15_), .QN(div_n162) );
  DFFX1_LVT div_divisor_reg_16_ ( .D(div_N339), .CLK(div_n294), .Q(
        div_divisor_16_) );
  DFFX1_LVT div_divisor_reg_17_ ( .D(div_N340), .CLK(div_n294), .Q(
        div_divisor_17_) );
  DFFX1_LVT div_divisor_reg_18_ ( .D(div_N341), .CLK(div_n294), .Q(
        div_divisor_18_), .QN(div_n161) );
  DFFX1_LVT div_divisor_reg_19_ ( .D(div_N342), .CLK(div_n294), .Q(
        div_divisor_19_) );
  DFFX1_LVT div_divisor_reg_20_ ( .D(div_N343), .CLK(div_n294), .Q(
        div_divisor_20_) );
  DFFX1_LVT div_divisor_reg_21_ ( .D(div_N344), .CLK(div_n294), .Q(
        div_divisor_21_) );
  DFFX1_LVT div_divisor_reg_22_ ( .D(div_N345), .CLK(div_n294), .Q(
        div_divisor_22_), .QN(div_n190) );
  DFFX1_LVT div_divisor_reg_23_ ( .D(div_N346), .CLK(div_n294), .Q(
        div_divisor_23_) );
  DFFX1_LVT div_divisor_reg_24_ ( .D(div_N347), .CLK(div_n295), .Q(
        div_divisor_24_), .QN(div_n164) );
  DFFX1_LVT div_divisor_reg_25_ ( .D(div_N348), .CLK(div_n295), .Q(
        div_divisor_25_) );
  DFFX1_LVT div_divisor_reg_26_ ( .D(div_N349), .CLK(div_n295), .Q(
        div_divisor_26_), .QN(div_n196) );
  DFFX1_LVT div_divisor_reg_27_ ( .D(div_N350), .CLK(div_n295), .Q(
        div_divisor_27_) );
  DFFX1_LVT div_divisor_reg_28_ ( .D(div_N351), .CLK(div_n295), .Q(
        div_divisor_28_) );
  DFFX1_LVT div_divisor_reg_29_ ( .D(div_N352), .CLK(div_n295), .Q(
        div_divisor_29_) );
  DFFX1_LVT div_divisor_reg_30_ ( .D(div_N353), .CLK(div_n295), .Q(
        div_divisor_30_), .QN(div_n174) );
  DFFX1_LVT div_divisor_reg_31_ ( .D(div_N354), .CLK(div_n295), .Q(
        div_divisor_31_), .QN(div_n176) );
  DFFX1_LVT div_divisor_reg_32_ ( .D(div_N355), .CLK(div_n295), .Q(
        div_divisor_32_) );
  DFFX1_LVT div_divisor_reg_33_ ( .D(div_N356), .CLK(div_n295), .Q(
        div_divisor_33_) );
  DFFX1_LVT div_divisor_reg_34_ ( .D(div_N357), .CLK(div_n295), .Q(
        div_divisor_34_), .QN(div_n160) );
  DFFX1_LVT div_divisor_reg_35_ ( .D(div_N358), .CLK(div_n295), .Q(
        div_divisor_35_) );
  DFFX1_LVT div_divisor_reg_36_ ( .D(div_N359), .CLK(div_n297), .Q(
        div_divisor_36_) );
  DFFX1_LVT div_divisor_reg_37_ ( .D(div_N360), .CLK(div_n297), .Q(
        div_divisor_37_) );
  DFFX1_LVT div_divisor_reg_38_ ( .D(div_N361), .CLK(div_n297), .Q(
        div_divisor_38_), .QN(div_n192) );
  DFFX1_LVT div_divisor_reg_39_ ( .D(div_N362), .CLK(div_n297), .Q(
        div_divisor_39_) );
  DFFX1_LVT div_divisor_reg_40_ ( .D(div_N363), .CLK(div_n297), .Q(
        div_divisor_40_), .QN(div_n163) );
  DFFX1_LVT div_divisor_reg_41_ ( .D(div_N364), .CLK(div_n297), .Q(
        div_divisor_41_) );
  DFFX1_LVT div_divisor_reg_42_ ( .D(div_N365), .CLK(div_n297), .Q(
        div_divisor_42_), .QN(div_n185) );
  DFFX1_LVT div_divisor_reg_43_ ( .D(div_N366), .CLK(div_n297), .Q(
        div_divisor_43_) );
  DFFX1_LVT div_divisor_reg_44_ ( .D(div_N367), .CLK(div_n297), .Q(
        div_divisor_44_) );
  DFFX1_LVT div_divisor_reg_45_ ( .D(div_N368), .CLK(div_n297), .Q(
        div_divisor_45_), .QN(div_n173) );
  DFFX1_LVT div_divisor_reg_46_ ( .D(div_N369), .CLK(div_n297), .Q(
        div_divisor_46_), .QN(div_n194) );
  DFFX1_LVT div_divisor_reg_47_ ( .D(div_N370), .CLK(div_n297), .Q(
        div_divisor_47_), .QN(div_n178) );
  DFFX1_LVT div_divisor_reg_48_ ( .D(div_N371), .CLK(div_n298), .Q(
        div_divisor_48_) );
  DFFX1_LVT div_divisor_reg_49_ ( .D(div_N372), .CLK(div_n298), .Q(
        div_divisor_49_) );
  DFFX1_LVT div_divisor_reg_50_ ( .D(div_N373), .CLK(div_n298), .Q(
        div_divisor_50_), .QN(div_n159) );
  DFFX1_LVT div_divisor_reg_51_ ( .D(div_N374), .CLK(div_n298), .Q(
        div_divisor_51_) );
  DFFX1_LVT div_divisor_reg_52_ ( .D(div_N375), .CLK(div_n298), .Q(
        div_divisor_52_) );
  DFFX1_LVT div_divisor_reg_53_ ( .D(div_N376), .CLK(div_n298), .Q(
        div_divisor_53_) );
  DFFX1_LVT div_divisor_reg_54_ ( .D(div_N377), .CLK(div_n298), .Q(
        div_divisor_54_), .QN(div_n195) );
  DFFX1_LVT div_divisor_reg_55_ ( .D(div_N378), .CLK(div_n298), .Q(
        div_divisor_55_) );
  DFFX1_LVT div_divisor_reg_56_ ( .D(div_N379), .CLK(div_n298), .Q(
        div_divisor_56_) );
  DFFX1_LVT div_divisor_reg_57_ ( .D(div_N380), .CLK(div_n298), .Q(
        div_divisor_57_) );
  DFFX1_LVT div_divisor_reg_58_ ( .D(div_N381), .CLK(div_n298), .Q(
        div_divisor_58_), .QN(div_n179) );
  DFFX1_LVT div_divisor_reg_59_ ( .D(div_N382), .CLK(div_n298), .Q(
        div_divisor_59_), .QN(div_n180) );
  DFFX1_LVT div_divisor_reg_60_ ( .D(div_N383), .CLK(div_n299), .Q(
        div_divisor_60_) );
  DFFX1_LVT div_divisor_reg_61_ ( .D(div_N384), .CLK(div_n299), .Q(
        div_divisor_61_) );
  DFFX1_LVT div_divisor_reg_62_ ( .D(div_N385), .CLK(div_n299), .Q(
        div_divisor_62_), .QN(div_n177) );
  DFFX1_LVT div_divisor_reg_63_ ( .D(div_N386), .CLK(div_n299), .Q(
        div_divisor_63_), .QN(div_n175) );
  DFFX1_LVT div_divisor_reg_64_ ( .D(div_N387), .CLK(div_n299), .Q(
        div_divisor_64_) );
  DFFX1_LVT div_neg_out_reg ( .D(div_n793), .CLK(div_net34695), .Q(div_neg_out), .QN(div_n212) );
  DFFX1_LVT div_count_reg_1_ ( .D(div_N295), .CLK(div_net34695), .Q(
        div_n_T_69_4_), .QN(div_n148) );
  DFFX1_LVT div_count_reg_2_ ( .D(div_N296), .CLK(div_net34695), .Q(
        div_n_T_71_39_), .QN(div_n210) );
  DFFX1_LVT div_count_reg_3_ ( .D(div_N297), .CLK(div_net34695), .Q(
        div_n_T_69_6_), .QN(div_n198) );
  DFFX1_LVT div_count_reg_4_ ( .D(div_N298), .CLK(div_net34695), .Q(
        div_n_T_69_7_) );
  DFFX1_LVT div_count_reg_5_ ( .D(div_N299), .CLK(div_net34695), .Q(
        div_n_T_69_8_), .QN(div_n197) );
  DFFSSRX1_LVT div_count_reg_6_ ( .D(div_n783), .SETB(div_n200), .RSTB(
        div_n_T_97_6_), .CLK(div_net34695), .Q(div_n_T_69_9_), .QN(div_n155)
         );
  DFFX1_LVT div_req_tag_reg_0_ ( .D(io_dmem_req_bits_tag[1]), .CLK(
        div_net34690), .Q(div_io_resp_bits_tag[0]) );
  DFFX1_LVT div_req_tag_reg_1_ ( .D(io_dmem_req_bits_tag[2]), .CLK(
        div_net34690), .QN(div_io_resp_bits_tag[1]) );
  DFFX1_LVT div_req_tag_reg_2_ ( .D(io_dmem_req_bits_tag[3]), .CLK(
        div_net34690), .Q(div_io_resp_bits_tag[2]) );
  DFFX1_LVT div_req_tag_reg_3_ ( .D(io_dmem_req_bits_tag[4]), .CLK(
        div_net34690), .QN(div_io_resp_bits_tag[3]) );
  DFFX1_LVT div_req_tag_reg_4_ ( .D(io_dmem_req_bits_tag[5]), .CLK(
        div_net34690), .QN(div_io_resp_bits_tag[4]) );
  DFFX1_LVT div_req_dw_reg ( .D(alu_io_dw), .CLK(div_net34690), .Q(div_n206), 
        .QN(div_n156) );
  DFFX1_LVT div_state_reg_2_ ( .D(div_N285), .CLK(div_net34700), .Q(div_n154), 
        .QN(div_n217) );
  DFFX1_LVT div_state_reg_1_ ( .D(div_N284), .CLK(div_net34700), .Q(div_n184), 
        .QN(div_n219) );
  DFFX1_LVT div_state_reg_0_ ( .D(div_N283), .CLK(div_net34700), .Q(div_n150), 
        .QN(div_n220) );
  DFFX1_LVT div_remainder_reg_31_ ( .D(div_N425), .CLK(div_n285), .Q(
        div_n_T_51_31_), .QN(div_n263) );
  DFFX1_LVT div_remainder_reg_30_ ( .D(div_N424), .CLK(div_n285), .Q(
        div_n_T_51_30_), .QN(div_n264) );
  DFFX1_LVT div_remainder_reg_29_ ( .D(div_N423), .CLK(div_n285), .Q(
        div_n_T_51_29_), .QN(div_n181) );
  DFFX1_LVT div_remainder_reg_28_ ( .D(div_N422), .CLK(div_n285), .Q(
        div_n_T_51_28_), .QN(div_n266) );
  DFFX1_LVT div_remainder_reg_27_ ( .D(div_N421), .CLK(div_n285), .Q(
        div_n_T_51_27_), .QN(div_n267) );
  DFFX1_LVT div_remainder_reg_26_ ( .D(div_N420), .CLK(div_n285), .Q(
        div_n_T_51_26_), .QN(div_n268) );
  DFFX1_LVT div_remainder_reg_25_ ( .D(div_N419), .CLK(div_n285), .Q(
        div_n_T_51_25_), .QN(div_n269) );
  DFFX1_LVT div_remainder_reg_24_ ( .D(div_N418), .CLK(div_n285), .Q(
        div_n_T_51_24_), .QN(div_n270) );
  DFFX1_LVT div_remainder_reg_23_ ( .D(div_N417), .CLK(div_n285), .Q(
        div_n_T_51_23_), .QN(div_n272) );
  DFFX1_LVT div_remainder_reg_22_ ( .D(div_N416), .CLK(div_n285), .Q(
        div_n_T_51_22_), .QN(div_n273) );
  DFFX1_LVT div_remainder_reg_21_ ( .D(div_N415), .CLK(div_n287), .Q(
        div_n_T_51_21_), .QN(div_n274) );
  DFFX1_LVT div_remainder_reg_20_ ( .D(div_N414), .CLK(div_n287), .Q(
        div_n_T_51_20_), .QN(div_n275) );
  DFFX1_LVT div_remainder_reg_19_ ( .D(div_N413), .CLK(div_n287), .Q(
        div_n_T_51_19_), .QN(div_n152) );
  DFFX1_LVT div_remainder_reg_18_ ( .D(div_N412), .CLK(div_n287), .Q(
        div_n_T_51_18_), .QN(div_n277) );
  DFFX1_LVT div_remainder_reg_17_ ( .D(div_N411), .CLK(div_n287), .Q(
        div_n_T_51_17_), .QN(div_n278) );
  DFFX1_LVT div_remainder_reg_16_ ( .D(div_N410), .CLK(div_n287), .Q(
        div_n_T_51_16_), .QN(div_n183) );
  DFFX1_LVT div_remainder_reg_15_ ( .D(div_N409), .CLK(div_n287), .Q(
        div_n_T_51_15_), .QN(div_n281) );
  DFFX1_LVT div_remainder_reg_14_ ( .D(div_N408), .CLK(div_n287), .Q(
        div_n_T_51_14_), .QN(div_n282) );
  DFFX1_LVT div_remainder_reg_13_ ( .D(div_N407), .CLK(div_n287), .Q(
        div_n_T_51_13_), .QN(div_n283) );
  DFFX1_LVT div_remainder_reg_12_ ( .D(div_N406), .CLK(div_n287), .Q(
        div_n_T_51_12_), .QN(div_n284) );
  DFFX1_LVT div_remainder_reg_11_ ( .D(div_N405), .CLK(div_n287), .Q(
        div_n_T_51_11_), .QN(div_n153) );
  DFFX1_LVT div_remainder_reg_10_ ( .D(div_N404), .CLK(div_n287), .Q(
        div_n_T_51_10_), .QN(div_n286) );
  DFFX1_LVT div_remainder_reg_9_ ( .D(div_N403), .CLK(div_n288), .Q(
        div_n_T_51_9_), .QN(div_n147) );
  DFFX1_LVT div_remainder_reg_8_ ( .D(div_N402), .CLK(div_n288), .Q(
        div_n_T_51_8_), .QN(div_n186) );
  DFFX1_LVT div_remainder_reg_7_ ( .D(div_N401), .CLK(div_n288), .Q(
        div_n_T_51_7_), .QN(div_n290) );
  DFFX1_LVT div_remainder_reg_6_ ( .D(div_N400), .CLK(div_n288), .Q(
        div_n_T_51_6_), .QN(div_n291) );
  DFFX1_LVT div_remainder_reg_5_ ( .D(div_N399), .CLK(div_n288), .Q(
        div_n_T_51_5_), .QN(div_n292) );
  DFFX1_LVT div_remainder_reg_4_ ( .D(div_N398), .CLK(div_n288), .Q(
        div_n_T_51_4_), .QN(div_n293) );
  DFFX1_LVT div_remainder_reg_3_ ( .D(div_N397), .CLK(div_n288), .Q(
        div_n_T_51_3_) );
  DFFX1_LVT div_remainder_reg_2_ ( .D(div_N396), .CLK(div_n288), .QN(div_n208)
         );
  DFFX1_LVT div_remainder_reg_1_ ( .D(div_N395), .CLK(div_n288), .Q(
        div_n_T_51_1_), .QN(div_n296) );
  DFFX1_LVT div_remainder_reg_0_ ( .D(div_N394), .CLK(div_n288), .Q(
        div_n_T_51_0_) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_1 div_clk_gate_remainder_reg ( .CLK(n3785), .EN(
        div_N493), .ENCLK(div_net34705), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_2 div_clk_gate_state_reg ( .CLK(n3785), .EN(
        div_N282), .ENCLK(div_net34700), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_3 div_clk_gate_count_reg ( .CLK(n3785), .EN(
        div_N293), .ENCLK(div_net34695), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_4 div_clk_gate_req_dw_reg ( .CLK(n3785), .EN(
        div_n235), .ENCLK(div_net34690), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_0 div_clk_gate_divisor_reg ( .CLK(n3785), .EN(
        div_N322), .ENCLK(div_net34684), .TE(1'b0) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2790 ( .A1(div_n301), .A2(
        div_divisor_0_), .Y(div_DP_OP_279J39_124_314_n2787) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2789 ( .A1(
        div_DP_OP_279J39_124_314_n2787), .A2(div_DP_OP_279J39_124_314_n2588), 
        .Y(div_DP_OP_279J39_124_314_n1593) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U2788 ( .A0(div_n_T_51_72_), .B0(
        div_DP_OP_279J39_124_314_n2787), .SO(div_DP_OP_279J39_124_314_n1594)
         );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2787 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2583), .Y(div_DP_OP_279J39_124_314_n1653) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2786 ( .A1(div_n301), .A2(
        div_divisor_62_), .Y(div_DP_OP_279J39_124_314_n1654) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2785 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2582), .Y(div_DP_OP_279J39_124_314_n1655) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2784 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2581), .Y(div_DP_OP_279J39_124_314_n1656) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2783 ( .A1(div_n301), .A2(
        div_divisor_59_), .Y(div_DP_OP_279J39_124_314_n1657) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2782 ( .A1(div_n301), .A2(
        div_divisor_58_), .Y(div_DP_OP_279J39_124_314_n1658) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2781 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2580), .Y(div_DP_OP_279J39_124_314_n1659) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2780 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2579), .Y(div_DP_OP_279J39_124_314_n1660) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2779 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2578), .Y(div_DP_OP_279J39_124_314_n1661) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2778 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2577), .Y(div_DP_OP_279J39_124_314_n1662) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2777 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2576), .Y(div_DP_OP_279J39_124_314_n1663) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2776 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2575), .Y(div_DP_OP_279J39_124_314_n1664) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2775 ( .A1(div_n301), .A2(
        div_divisor_51_), .Y(div_DP_OP_279J39_124_314_n1665) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2774 ( .A1(div_n301), .A2(
        div_divisor_50_), .Y(div_DP_OP_279J39_124_314_n1666) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2773 ( .A1(div_n301), .A2(
        div_divisor_49_), .Y(div_DP_OP_279J39_124_314_n1667) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2772 ( .A1(div_n301), .A2(
        div_divisor_48_), .Y(div_DP_OP_279J39_124_314_n1668) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2771 ( .A1(div_n301), .A2(
        div_divisor_47_), .Y(div_DP_OP_279J39_124_314_n1669) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2770 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2574), .Y(div_DP_OP_279J39_124_314_n1670) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2769 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2573), .Y(div_DP_OP_279J39_124_314_n1671) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2768 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2572), .Y(div_DP_OP_279J39_124_314_n1672) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2767 ( .A1(div_n301), .A2(
        div_divisor_43_), .Y(div_DP_OP_279J39_124_314_n1673) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2766 ( .A1(div_n301), .A2(
        div_divisor_42_), .Y(div_DP_OP_279J39_124_314_n1674) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2765 ( .A1(div_n301), .A2(
        div_divisor_41_), .Y(div_DP_OP_279J39_124_314_n1675) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2764 ( .A1(div_n301), .A2(
        div_divisor_40_), .Y(div_DP_OP_279J39_124_314_n1676) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2763 ( .A1(div_n301), .A2(
        div_divisor_39_), .Y(div_DP_OP_279J39_124_314_n1677) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2762 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2571), .Y(div_DP_OP_279J39_124_314_n1678) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2761 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2570), .Y(div_DP_OP_279J39_124_314_n1679) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2760 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2569), .Y(div_DP_OP_279J39_124_314_n1680) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2759 ( .A1(div_n301), .A2(
        div_divisor_35_), .Y(div_DP_OP_279J39_124_314_n1681) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2758 ( .A1(div_n301), .A2(
        div_divisor_34_), .Y(div_DP_OP_279J39_124_314_n1682) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2757 ( .A1(div_n301), .A2(
        div_divisor_33_), .Y(div_DP_OP_279J39_124_314_n1683) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2756 ( .A1(div_n301), .A2(
        div_divisor_32_), .Y(div_DP_OP_279J39_124_314_n1684) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2755 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2568), .Y(div_DP_OP_279J39_124_314_n1685) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2754 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2567), .Y(div_DP_OP_279J39_124_314_n1686) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2753 ( .A1(div_n301), .A2(
        div_divisor_29_), .Y(div_DP_OP_279J39_124_314_n1687) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2752 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2566), .Y(div_DP_OP_279J39_124_314_n1688) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2751 ( .A1(div_n301), .A2(
        div_divisor_27_), .Y(div_DP_OP_279J39_124_314_n1689) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2750 ( .A1(div_n301), .A2(
        div_divisor_26_), .Y(div_DP_OP_279J39_124_314_n1690) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2749 ( .A1(div_n301), .A2(
        div_divisor_25_), .Y(div_DP_OP_279J39_124_314_n1691) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2748 ( .A1(div_n301), .A2(
        div_divisor_24_), .Y(div_DP_OP_279J39_124_314_n1692) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2747 ( .A1(div_n301), .A2(
        div_divisor_23_), .Y(div_DP_OP_279J39_124_314_n1693) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2746 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2565), .Y(div_DP_OP_279J39_124_314_n1694) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2745 ( .A1(div_n301), .A2(
        div_divisor_21_), .Y(div_DP_OP_279J39_124_314_n1695) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2744 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2564), .Y(div_DP_OP_279J39_124_314_n1696) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2743 ( .A1(div_n301), .A2(
        div_divisor_19_), .Y(div_DP_OP_279J39_124_314_n1697) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2742 ( .A1(div_n301), .A2(
        div_divisor_18_), .Y(div_DP_OP_279J39_124_314_n1698) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2741 ( .A1(div_n301), .A2(
        div_divisor_17_), .Y(div_DP_OP_279J39_124_314_n1699) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2740 ( .A1(div_n301), .A2(
        div_divisor_16_), .Y(div_DP_OP_279J39_124_314_n1700) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2739 ( .A1(div_n301), .A2(
        div_divisor_15_), .Y(div_DP_OP_279J39_124_314_n1701) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2738 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2563), .Y(div_DP_OP_279J39_124_314_n1702) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2737 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2562), .Y(div_DP_OP_279J39_124_314_n1703) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2736 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2561), .Y(div_DP_OP_279J39_124_314_n1704) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2735 ( .A1(div_n301), .A2(
        div_divisor_11_), .Y(div_DP_OP_279J39_124_314_n1705) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2734 ( .A1(div_n301), .A2(
        div_divisor_10_), .Y(div_DP_OP_279J39_124_314_n1706) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2733 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2560), .Y(div_DP_OP_279J39_124_314_n1707) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2732 ( .A1(div_n301), .A2(
        div_divisor_8_), .Y(div_DP_OP_279J39_124_314_n1708) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2731 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2559), .Y(div_DP_OP_279J39_124_314_n1709) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2730 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2558), .Y(div_DP_OP_279J39_124_314_n1710) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2729 ( .A1(div_n301), .A2(
        div_divisor_5_), .Y(div_DP_OP_279J39_124_314_n1711) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2728 ( .A1(div_n301), .A2(
        div_DP_OP_279J39_124_314_n2557), .Y(div_DP_OP_279J39_124_314_n1712) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2727 ( .A1(div_n301), .A2(
        div_divisor_3_), .Y(div_DP_OP_279J39_124_314_n1713) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2726 ( .A1(div_n301), .A2(
        div_divisor_2_), .Y(div_DP_OP_279J39_124_314_n1714) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2725 ( .A1(div_n301), .A2(
        div_divisor_1_), .Y(div_DP_OP_279J39_124_314_n1715) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2724 ( .A1(div_divisor_64_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1717) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2723 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1718) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2722 ( .A1(div_divisor_62_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1719) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2721 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1720) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2720 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1721) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2719 ( .A1(div_divisor_59_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1722) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2718 ( .A1(div_divisor_58_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1723) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2717 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1724) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2716 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1725) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2715 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1726) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2714 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1727) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2713 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1728) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2712 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1729) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2711 ( .A1(div_divisor_51_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1730) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2710 ( .A1(div_divisor_50_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1731) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2709 ( .A1(div_divisor_49_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1732) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2708 ( .A1(div_divisor_48_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1733) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2707 ( .A1(div_divisor_47_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1734) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2706 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1735) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2705 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1736) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2704 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1737) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2703 ( .A1(div_divisor_43_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1738) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2702 ( .A1(div_divisor_42_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1739) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2701 ( .A1(div_divisor_41_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1740) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2700 ( .A1(div_divisor_40_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1741) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2699 ( .A1(div_divisor_39_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1742) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2698 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1743) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2697 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1744) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2696 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1745) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2695 ( .A1(div_divisor_35_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1746) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2694 ( .A1(div_divisor_34_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1747) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2693 ( .A1(div_divisor_33_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1748) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2692 ( .A1(div_divisor_32_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1749) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2691 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1750) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2690 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1751) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2689 ( .A1(div_divisor_29_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1752) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2688 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1753) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2687 ( .A1(div_divisor_27_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1754) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2686 ( .A1(div_divisor_26_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1755) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2685 ( .A1(div_divisor_25_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1756) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2684 ( .A1(div_divisor_24_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1757) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2683 ( .A1(div_divisor_23_), .A2(
        div_n_T_51_7_), .Y(div_DP_OP_279J39_124_314_n1758) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2682 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n_T_51_7_), .Y(
        div_DP_OP_279J39_124_314_n1759) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2681 ( .A1(div_divisor_21_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1760) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2680 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_n_T_51_7_), .Y(
        div_DP_OP_279J39_124_314_n1761) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2679 ( .A1(div_divisor_19_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1762) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2678 ( .A1(div_divisor_18_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1763) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2677 ( .A1(div_divisor_17_), .A2(
        div_n_T_51_7_), .Y(div_DP_OP_279J39_124_314_n1764) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2676 ( .A1(div_divisor_16_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1765) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2675 ( .A1(div_divisor_15_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1766) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2674 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1767) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2673 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1768) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2672 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n_T_51_7_), .Y(
        div_DP_OP_279J39_124_314_n1769) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2671 ( .A1(div_divisor_11_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1770) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2670 ( .A1(div_divisor_10_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1771) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2669 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1772) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2668 ( .A1(div_divisor_8_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1773) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2667 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1774) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2666 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1775) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2665 ( .A1(div_divisor_5_), .A2(
        div_DP_OP_279J39_124_314_n2585), .Y(div_DP_OP_279J39_124_314_n1776) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2664 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_DP_OP_279J39_124_314_n2585), 
        .Y(div_DP_OP_279J39_124_314_n1777) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2663 ( .A1(div_divisor_3_), .A2(
        div_n_T_51_7_), .Y(div_DP_OP_279J39_124_314_n1778) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2662 ( .A1(div_divisor_2_), .A2(
        div_n_T_51_7_), .Y(div_DP_OP_279J39_124_314_n1779) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2661 ( .A1(div_divisor_1_), .A2(
        div_n_T_51_7_), .Y(div_DP_OP_279J39_124_314_n1780) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2660 ( .A1(div_divisor_0_), .A2(
        div_n_T_51_7_), .Y(div_DP_OP_279J39_124_314_n1781) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2659 ( .A1(div_divisor_64_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1782) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2658 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1783) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2657 ( .A1(div_divisor_62_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1784) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2656 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1785) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2655 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1786) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2654 ( .A1(div_divisor_59_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1787) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2653 ( .A1(div_divisor_58_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1788) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2652 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1789) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2651 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1790) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2650 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1791) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2649 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1792) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2648 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1793) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2647 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1794) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2646 ( .A1(div_divisor_51_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1795) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2645 ( .A1(div_divisor_50_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1796) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2644 ( .A1(div_divisor_49_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1797) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2643 ( .A1(div_divisor_48_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1798) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2642 ( .A1(div_divisor_47_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1799) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2641 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1800) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2640 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1801) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2639 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1802) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2638 ( .A1(div_divisor_43_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1803) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2637 ( .A1(div_divisor_42_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1804) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2636 ( .A1(div_divisor_41_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1805) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2635 ( .A1(div_divisor_40_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1806) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2634 ( .A1(div_divisor_39_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1807) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2633 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1808) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2632 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1809) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2631 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1810) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2630 ( .A1(div_divisor_35_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1811) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2629 ( .A1(div_divisor_34_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1812) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2628 ( .A1(div_divisor_33_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1813) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2627 ( .A1(div_divisor_32_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1814) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2626 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1815) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2625 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1816) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2624 ( .A1(div_divisor_29_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1817) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2623 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1818) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2622 ( .A1(div_divisor_27_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1819) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2621 ( .A1(div_divisor_26_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1820) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2620 ( .A1(div_divisor_25_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1821) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2619 ( .A1(div_divisor_24_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1822) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2618 ( .A1(div_divisor_23_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1823) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2617 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1824) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2616 ( .A1(div_divisor_21_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1825) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2615 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1826) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2614 ( .A1(div_divisor_19_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1827) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2613 ( .A1(div_divisor_18_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1828) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2612 ( .A1(div_divisor_17_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1829) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2611 ( .A1(div_divisor_16_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1830) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2610 ( .A1(div_divisor_15_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1831) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2609 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1832) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2608 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1833) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2607 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1834) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2606 ( .A1(div_divisor_11_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1835) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2605 ( .A1(div_divisor_10_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1836) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2604 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1837) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2603 ( .A1(div_divisor_8_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1838) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2602 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1839) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2601 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1840) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2600 ( .A1(div_divisor_5_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1841) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2599 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_n307), .Y(
        div_DP_OP_279J39_124_314_n1842) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2598 ( .A1(div_divisor_3_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1843) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2597 ( .A1(div_divisor_2_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1844) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2596 ( .A1(div_divisor_1_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1845) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2595 ( .A1(div_divisor_0_), .A2(
        div_n307), .Y(div_DP_OP_279J39_124_314_n1846) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2594 ( .A1(div_divisor_64_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1847) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2593 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1848) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2592 ( .A1(div_divisor_62_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1849) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2591 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1850) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2590 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1851) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2589 ( .A1(div_divisor_59_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1852) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2588 ( .A1(div_divisor_58_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1853) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2587 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1854) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2586 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1855) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2585 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1856) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2584 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1857) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2583 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1858) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2582 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1859) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2581 ( .A1(div_divisor_51_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1860) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2580 ( .A1(div_divisor_50_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1861) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2579 ( .A1(div_divisor_49_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1862) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2578 ( .A1(div_divisor_48_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1863) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2577 ( .A1(div_divisor_47_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1864) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2576 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1865) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2575 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1866) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2574 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1867) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2573 ( .A1(div_divisor_43_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1868) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2572 ( .A1(div_divisor_42_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1869) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2571 ( .A1(div_divisor_41_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1870) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2570 ( .A1(div_divisor_40_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1871) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2569 ( .A1(div_divisor_39_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1872) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2568 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1873) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2567 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1874) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2566 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1875) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2565 ( .A1(div_divisor_35_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1876) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2564 ( .A1(div_divisor_34_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1877) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2563 ( .A1(div_divisor_33_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1878) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2562 ( .A1(div_divisor_32_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1879) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2561 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1880) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2560 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1881) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2559 ( .A1(div_divisor_29_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1882) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2558 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1883) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2557 ( .A1(div_divisor_27_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1884) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2556 ( .A1(div_divisor_26_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1885) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2555 ( .A1(div_divisor_25_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1886) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2554 ( .A1(div_divisor_24_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1887) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2553 ( .A1(div_divisor_23_), .A2(
        div_n_T_51_5_), .Y(div_DP_OP_279J39_124_314_n1888) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2552 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n_T_51_5_), .Y(
        div_DP_OP_279J39_124_314_n1889) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2551 ( .A1(div_divisor_21_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1890) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2550 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1891) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2549 ( .A1(div_divisor_19_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1892) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2548 ( .A1(div_divisor_18_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1893) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2547 ( .A1(div_divisor_17_), .A2(
        div_n_T_51_5_), .Y(div_DP_OP_279J39_124_314_n1894) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2546 ( .A1(div_divisor_16_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1895) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2545 ( .A1(div_divisor_15_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1896) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2544 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1897) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2543 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1898) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2542 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n_T_51_5_), .Y(
        div_DP_OP_279J39_124_314_n1899) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2541 ( .A1(div_divisor_11_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1900) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2540 ( .A1(div_divisor_10_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1901) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2539 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1902) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2538 ( .A1(div_divisor_8_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1903) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2537 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1904) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2536 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1905) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2535 ( .A1(div_divisor_5_), .A2(
        div_DP_OP_279J39_124_314_n2584), .Y(div_DP_OP_279J39_124_314_n1906) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2534 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_DP_OP_279J39_124_314_n2584), 
        .Y(div_DP_OP_279J39_124_314_n1907) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2533 ( .A1(div_divisor_3_), .A2(
        div_n_T_51_5_), .Y(div_DP_OP_279J39_124_314_n1908) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2532 ( .A1(div_divisor_2_), .A2(
        div_n_T_51_5_), .Y(div_DP_OP_279J39_124_314_n1909) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2531 ( .A1(div_divisor_1_), .A2(
        div_n_T_51_5_), .Y(div_DP_OP_279J39_124_314_n1910) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2530 ( .A1(div_divisor_0_), .A2(
        div_n_T_51_5_), .Y(div_DP_OP_279J39_124_314_n1911) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2529 ( .A1(div_divisor_64_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1912) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2528 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1913) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2527 ( .A1(div_divisor_62_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1914) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2526 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1915) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2525 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1916) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2524 ( .A1(div_divisor_59_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1917) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2523 ( .A1(div_divisor_58_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1918) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2522 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1919) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2521 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1920) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2520 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1921) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2519 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1922) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2518 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1923) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2517 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1924) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2516 ( .A1(div_divisor_51_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1925) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2515 ( .A1(div_divisor_50_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1926) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2514 ( .A1(div_divisor_49_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1927) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2513 ( .A1(div_divisor_48_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1928) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2512 ( .A1(div_divisor_47_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1929) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2511 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1930) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2510 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1931) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2509 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1932) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2508 ( .A1(div_divisor_43_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1933) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2507 ( .A1(div_divisor_42_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1934) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2506 ( .A1(div_divisor_41_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1935) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2505 ( .A1(div_divisor_40_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1936) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2504 ( .A1(div_divisor_39_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1937) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2503 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1938) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2502 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1939) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2501 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1940) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2500 ( .A1(div_divisor_35_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1941) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2499 ( .A1(div_divisor_34_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1942) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2498 ( .A1(div_divisor_33_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1943) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2497 ( .A1(div_divisor_32_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1944) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2496 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1945) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2495 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1946) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2494 ( .A1(div_divisor_29_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1947) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2493 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1948) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2492 ( .A1(div_divisor_27_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1949) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2491 ( .A1(div_divisor_26_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1950) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2490 ( .A1(div_divisor_25_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1951) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2489 ( .A1(div_divisor_24_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1952) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2488 ( .A1(div_divisor_23_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1953) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2487 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1954) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2486 ( .A1(div_divisor_21_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1955) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2485 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1956) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2484 ( .A1(div_divisor_19_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1957) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2483 ( .A1(div_divisor_18_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1958) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2482 ( .A1(div_divisor_17_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1959) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2481 ( .A1(div_divisor_16_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1960) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2480 ( .A1(div_divisor_15_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1961) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2479 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1962) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2478 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1963) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2477 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1964) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2476 ( .A1(div_divisor_11_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1965) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2475 ( .A1(div_divisor_10_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1966) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2474 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1967) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2473 ( .A1(div_divisor_8_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1968) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2472 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1969) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2471 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1970) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2470 ( .A1(div_divisor_5_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1971) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2469 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_n306), .Y(
        div_DP_OP_279J39_124_314_n1972) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2468 ( .A1(div_divisor_3_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1973) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2467 ( .A1(div_divisor_2_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1974) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2466 ( .A1(div_divisor_1_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1975) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2465 ( .A1(div_divisor_0_), .A2(
        div_n306), .Y(div_DP_OP_279J39_124_314_n1976) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2464 ( .A1(div_divisor_64_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1977) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2463 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1978) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2462 ( .A1(div_divisor_62_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1979) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2461 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1980) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2460 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1981) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2459 ( .A1(div_divisor_59_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1982) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2458 ( .A1(div_divisor_58_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1983) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2457 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1984) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2456 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1985) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2455 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1986) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2454 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1987) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2453 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1988) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2452 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1989) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2451 ( .A1(div_divisor_51_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1990) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2450 ( .A1(div_divisor_50_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1991) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2449 ( .A1(div_divisor_49_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1992) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2448 ( .A1(div_divisor_48_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1993) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2447 ( .A1(div_divisor_47_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1994) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2446 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1995) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2445 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1996) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2444 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n1997) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2443 ( .A1(div_divisor_43_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1998) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2442 ( .A1(div_divisor_42_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n1999) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2441 ( .A1(div_divisor_41_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2000) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2440 ( .A1(div_divisor_40_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2001) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2439 ( .A1(div_divisor_39_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2002) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2438 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2003) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2437 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2004) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2436 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2005) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2435 ( .A1(div_divisor_35_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2006) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2434 ( .A1(div_divisor_34_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2007) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2433 ( .A1(div_divisor_33_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2008) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2432 ( .A1(div_divisor_32_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2009) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2431 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2010) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2430 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2011) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2429 ( .A1(div_divisor_29_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2012) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2428 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2013) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2427 ( .A1(div_divisor_27_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2014) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2426 ( .A1(div_divisor_26_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2015) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2425 ( .A1(div_divisor_25_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2016) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2424 ( .A1(div_divisor_24_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2017) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2423 ( .A1(div_divisor_23_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2018) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2422 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2019) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2421 ( .A1(div_divisor_21_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2020) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2420 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2021) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2419 ( .A1(div_divisor_19_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2022) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2418 ( .A1(div_divisor_18_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2023) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2417 ( .A1(div_divisor_17_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2024) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2416 ( .A1(div_divisor_16_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2025) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2415 ( .A1(div_divisor_15_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2026) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2414 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2027) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2413 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2028) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2412 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2029) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2411 ( .A1(div_divisor_11_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2030) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2410 ( .A1(div_divisor_10_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2031) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2409 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2032) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2408 ( .A1(div_divisor_8_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2033) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2407 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2034) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2406 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2035) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2405 ( .A1(div_divisor_5_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2036) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2404 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_n305), .Y(
        div_DP_OP_279J39_124_314_n2037) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2403 ( .A1(div_divisor_3_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2038) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2402 ( .A1(div_divisor_2_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2039) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2401 ( .A1(div_divisor_1_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2040) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2400 ( .A1(div_divisor_0_), .A2(
        div_n305), .Y(div_DP_OP_279J39_124_314_n2041) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2399 ( .A1(div_divisor_64_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2042) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2398 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2043) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2397 ( .A1(div_divisor_62_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2044) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2396 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2045) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2395 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2046) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2394 ( .A1(div_divisor_59_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2047) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2393 ( .A1(div_divisor_58_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2048) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2392 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2049) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2391 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2050) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2390 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2051) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2389 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2052) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2388 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2053) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2387 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2054) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2386 ( .A1(div_divisor_51_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2055) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2385 ( .A1(div_divisor_50_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2056) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2384 ( .A1(div_divisor_49_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2057) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2383 ( .A1(div_divisor_48_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2058) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2382 ( .A1(div_divisor_47_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2059) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2381 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2060) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2380 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2061) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2379 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2062) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2378 ( .A1(div_divisor_43_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2063) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2377 ( .A1(div_divisor_42_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2064) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2376 ( .A1(div_divisor_41_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2065) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2375 ( .A1(div_divisor_40_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2066) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2374 ( .A1(div_divisor_39_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2067) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2373 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2068) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2372 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2069) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2371 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2070) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2370 ( .A1(div_divisor_35_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2071) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2369 ( .A1(div_divisor_34_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2072) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2368 ( .A1(div_divisor_33_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2073) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2367 ( .A1(div_divisor_32_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2074) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2366 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2075) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2365 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2076) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2364 ( .A1(div_divisor_29_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2077) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2363 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2078) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2362 ( .A1(div_divisor_27_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2079) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2361 ( .A1(div_divisor_26_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2080) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2360 ( .A1(div_divisor_25_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2081) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2359 ( .A1(div_divisor_24_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2082) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2358 ( .A1(div_divisor_23_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2083) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2357 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2084) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2356 ( .A1(div_divisor_21_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2085) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2355 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2086) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2354 ( .A1(div_divisor_19_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2087) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2353 ( .A1(div_divisor_18_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2088) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2352 ( .A1(div_divisor_17_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2089) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2351 ( .A1(div_divisor_16_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2090) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2350 ( .A1(div_divisor_15_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2091) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2349 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2092) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2348 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2093) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2347 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2094) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2346 ( .A1(div_divisor_11_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2095) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2345 ( .A1(div_divisor_10_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2096) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2344 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2097) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2343 ( .A1(div_divisor_8_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2098) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2342 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2099) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2341 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2100) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2340 ( .A1(div_divisor_5_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2101) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2339 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_n304), .Y(
        div_DP_OP_279J39_124_314_n2102) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2338 ( .A1(div_divisor_3_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2103) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2337 ( .A1(div_divisor_2_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2104) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2336 ( .A1(div_divisor_1_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2105) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2335 ( .A1(div_divisor_0_), .A2(
        div_n304), .Y(div_DP_OP_279J39_124_314_n2106) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2334 ( .A1(div_divisor_64_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2107) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2333 ( .A1(
        div_DP_OP_279J39_124_314_n2583), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2108) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2332 ( .A1(div_divisor_62_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2109) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2331 ( .A1(
        div_DP_OP_279J39_124_314_n2582), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2110) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2330 ( .A1(
        div_DP_OP_279J39_124_314_n2581), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2111) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2329 ( .A1(div_divisor_59_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2112) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2328 ( .A1(div_divisor_58_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2113) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2327 ( .A1(
        div_DP_OP_279J39_124_314_n2580), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2114) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2326 ( .A1(
        div_DP_OP_279J39_124_314_n2579), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2115) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2325 ( .A1(
        div_DP_OP_279J39_124_314_n2578), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2116) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2324 ( .A1(
        div_DP_OP_279J39_124_314_n2577), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2117) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2323 ( .A1(
        div_DP_OP_279J39_124_314_n2576), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2118) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2322 ( .A1(
        div_DP_OP_279J39_124_314_n2575), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2119) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2321 ( .A1(div_divisor_51_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2120) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2320 ( .A1(div_divisor_50_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2121) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2319 ( .A1(div_divisor_49_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2122) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2318 ( .A1(div_divisor_48_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2123) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2317 ( .A1(div_divisor_47_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2124) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2316 ( .A1(
        div_DP_OP_279J39_124_314_n2574), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2125) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2315 ( .A1(
        div_DP_OP_279J39_124_314_n2573), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2126) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2314 ( .A1(
        div_DP_OP_279J39_124_314_n2572), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2127) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2313 ( .A1(div_divisor_43_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2128) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2312 ( .A1(div_divisor_42_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2129) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2311 ( .A1(div_divisor_41_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2130) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2310 ( .A1(div_divisor_40_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2131) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2309 ( .A1(div_divisor_39_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2132) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2308 ( .A1(
        div_DP_OP_279J39_124_314_n2571), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2133) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2307 ( .A1(
        div_DP_OP_279J39_124_314_n2570), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2134) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2306 ( .A1(
        div_DP_OP_279J39_124_314_n2569), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2135) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2305 ( .A1(div_divisor_35_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2136) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2304 ( .A1(div_divisor_34_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2137) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2303 ( .A1(div_divisor_33_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2138) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2302 ( .A1(div_divisor_32_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2139) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2301 ( .A1(
        div_DP_OP_279J39_124_314_n2568), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2140) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2300 ( .A1(
        div_DP_OP_279J39_124_314_n2567), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2141) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2299 ( .A1(div_divisor_29_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2142) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2298 ( .A1(
        div_DP_OP_279J39_124_314_n2566), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2143) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2297 ( .A1(div_divisor_27_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2144) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2296 ( .A1(div_divisor_26_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2145) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2295 ( .A1(div_divisor_25_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2146) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2294 ( .A1(div_divisor_24_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2147) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2293 ( .A1(div_divisor_23_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2148) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2292 ( .A1(
        div_DP_OP_279J39_124_314_n2565), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2149) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2291 ( .A1(div_divisor_21_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2150) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2290 ( .A1(
        div_DP_OP_279J39_124_314_n2564), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2151) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2289 ( .A1(div_divisor_19_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2152) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2288 ( .A1(div_divisor_18_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2153) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2287 ( .A1(div_divisor_17_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2154) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2286 ( .A1(div_divisor_16_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2155) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2285 ( .A1(div_divisor_15_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2156) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2284 ( .A1(
        div_DP_OP_279J39_124_314_n2563), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2157) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2283 ( .A1(
        div_DP_OP_279J39_124_314_n2562), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2158) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2282 ( .A1(
        div_DP_OP_279J39_124_314_n2561), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2159) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2281 ( .A1(div_divisor_11_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2160) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2280 ( .A1(div_divisor_10_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2161) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2279 ( .A1(
        div_DP_OP_279J39_124_314_n2560), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2162) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2278 ( .A1(div_divisor_8_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2163) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2277 ( .A1(
        div_DP_OP_279J39_124_314_n2559), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2164) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2276 ( .A1(
        div_DP_OP_279J39_124_314_n2558), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2165) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2275 ( .A1(div_divisor_5_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2166) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2274 ( .A1(
        div_DP_OP_279J39_124_314_n2557), .A2(div_n303), .Y(
        div_DP_OP_279J39_124_314_n2167) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2273 ( .A1(div_divisor_3_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2168) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2272 ( .A1(div_divisor_2_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2169) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2271 ( .A1(div_divisor_1_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2170) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2270 ( .A1(div_divisor_0_), .A2(
        div_n303), .Y(div_DP_OP_279J39_124_314_n2171) );
  NAND2X0_LVT div_DP_OP_279J39_124_314_U2269 ( .A1(div_divisor_64_), .A2(
        div_n302), .Y(div_DP_OP_279J39_124_314_n2172) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2268 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2583), .Y(div_DP_OP_279J39_124_314_n2173) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2267 ( .A1(div_n302), .A2(
        div_divisor_62_), .Y(div_DP_OP_279J39_124_314_n2174) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2266 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2582), .Y(div_DP_OP_279J39_124_314_n2175) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2265 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2581), .Y(div_DP_OP_279J39_124_314_n2176) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2264 ( .A1(div_n302), .A2(
        div_divisor_59_), .Y(div_DP_OP_279J39_124_314_n2177) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2263 ( .A1(div_n302), .A2(
        div_divisor_58_), .Y(div_DP_OP_279J39_124_314_n2178) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2262 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2580), .Y(div_DP_OP_279J39_124_314_n2179) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2261 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2579), .Y(div_DP_OP_279J39_124_314_n2180) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2260 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2578), .Y(div_DP_OP_279J39_124_314_n2181) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2259 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2577), .Y(div_DP_OP_279J39_124_314_n2182) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2258 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2576), .Y(div_DP_OP_279J39_124_314_n2183) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2257 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2575), .Y(div_DP_OP_279J39_124_314_n2184) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2256 ( .A1(div_n302), .A2(
        div_divisor_51_), .Y(div_DP_OP_279J39_124_314_n2185) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2255 ( .A1(div_n302), .A2(
        div_divisor_50_), .Y(div_DP_OP_279J39_124_314_n2186) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2254 ( .A1(div_n302), .A2(
        div_divisor_49_), .Y(div_DP_OP_279J39_124_314_n2187) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2253 ( .A1(div_n302), .A2(
        div_divisor_48_), .Y(div_DP_OP_279J39_124_314_n2188) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2252 ( .A1(div_n302), .A2(
        div_divisor_47_), .Y(div_DP_OP_279J39_124_314_n2189) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2251 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2574), .Y(div_DP_OP_279J39_124_314_n2190) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2250 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2573), .Y(div_DP_OP_279J39_124_314_n2191) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2249 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2572), .Y(div_DP_OP_279J39_124_314_n2192) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2248 ( .A1(div_n302), .A2(
        div_divisor_43_), .Y(div_DP_OP_279J39_124_314_n2193) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2247 ( .A1(div_n302), .A2(
        div_divisor_42_), .Y(div_DP_OP_279J39_124_314_n2194) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2246 ( .A1(div_n302), .A2(
        div_divisor_41_), .Y(div_DP_OP_279J39_124_314_n2195) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2245 ( .A1(div_n302), .A2(
        div_divisor_40_), .Y(div_DP_OP_279J39_124_314_n2196) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2244 ( .A1(div_n302), .A2(
        div_divisor_39_), .Y(div_DP_OP_279J39_124_314_n2197) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2243 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2571), .Y(div_DP_OP_279J39_124_314_n2198) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2242 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2570), .Y(div_DP_OP_279J39_124_314_n2199) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2241 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2569), .Y(div_DP_OP_279J39_124_314_n2200) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2240 ( .A1(div_n302), .A2(
        div_divisor_35_), .Y(div_DP_OP_279J39_124_314_n2201) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2239 ( .A1(div_n302), .A2(
        div_divisor_34_), .Y(div_DP_OP_279J39_124_314_n2202) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2238 ( .A1(div_n302), .A2(
        div_divisor_33_), .Y(div_DP_OP_279J39_124_314_n2203) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2237 ( .A1(div_n302), .A2(
        div_divisor_32_), .Y(div_DP_OP_279J39_124_314_n2204) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2236 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2568), .Y(div_DP_OP_279J39_124_314_n2205) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2235 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2567), .Y(div_DP_OP_279J39_124_314_n2206) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2234 ( .A1(div_n302), .A2(
        div_divisor_29_), .Y(div_DP_OP_279J39_124_314_n2207) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2233 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2566), .Y(div_DP_OP_279J39_124_314_n2208) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2232 ( .A1(div_n302), .A2(
        div_divisor_27_), .Y(div_DP_OP_279J39_124_314_n2209) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2231 ( .A1(div_n302), .A2(
        div_divisor_26_), .Y(div_DP_OP_279J39_124_314_n2210) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2230 ( .A1(div_n302), .A2(
        div_divisor_25_), .Y(div_DP_OP_279J39_124_314_n2211) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2229 ( .A1(div_n302), .A2(
        div_divisor_24_), .Y(div_DP_OP_279J39_124_314_n2212) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2228 ( .A1(div_n302), .A2(
        div_divisor_23_), .Y(div_DP_OP_279J39_124_314_n2213) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2227 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2565), .Y(div_DP_OP_279J39_124_314_n2214) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2226 ( .A1(div_n302), .A2(
        div_divisor_21_), .Y(div_DP_OP_279J39_124_314_n2215) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2225 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2564), .Y(div_DP_OP_279J39_124_314_n2216) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2224 ( .A1(div_n302), .A2(
        div_divisor_19_), .Y(div_DP_OP_279J39_124_314_n2217) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2223 ( .A1(div_n302), .A2(
        div_divisor_18_), .Y(div_DP_OP_279J39_124_314_n2218) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2222 ( .A1(div_n302), .A2(
        div_divisor_17_), .Y(div_DP_OP_279J39_124_314_n2219) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2221 ( .A1(div_n302), .A2(
        div_divisor_16_), .Y(div_DP_OP_279J39_124_314_n2220) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2220 ( .A1(div_n302), .A2(
        div_divisor_15_), .Y(div_DP_OP_279J39_124_314_n2221) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2219 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2563), .Y(div_DP_OP_279J39_124_314_n2222) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2218 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2562), .Y(div_DP_OP_279J39_124_314_n2223) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2217 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2561), .Y(div_DP_OP_279J39_124_314_n2224) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2216 ( .A1(div_n302), .A2(
        div_divisor_11_), .Y(div_DP_OP_279J39_124_314_n2225) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2215 ( .A1(div_n302), .A2(
        div_divisor_10_), .Y(div_DP_OP_279J39_124_314_n2226) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2214 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2560), .Y(div_DP_OP_279J39_124_314_n2227) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2213 ( .A1(div_n302), .A2(
        div_divisor_8_), .Y(div_DP_OP_279J39_124_314_n2228) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2212 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2559), .Y(div_DP_OP_279J39_124_314_n2229) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2211 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2558), .Y(div_DP_OP_279J39_124_314_n2230) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2210 ( .A1(div_n302), .A2(
        div_divisor_5_), .Y(div_DP_OP_279J39_124_314_n2231) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2209 ( .A1(div_n302), .A2(
        div_DP_OP_279J39_124_314_n2557), .Y(div_DP_OP_279J39_124_314_n2232) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2208 ( .A1(div_n302), .A2(
        div_divisor_3_), .Y(div_DP_OP_279J39_124_314_n2233) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2207 ( .A1(div_n302), .A2(
        div_divisor_2_), .Y(div_DP_OP_279J39_124_314_n2234) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2206 ( .A1(div_n302), .A2(
        div_divisor_1_), .Y(div_DP_OP_279J39_124_314_n2235) );
  NAND3X0_LVT div_DP_OP_279J39_124_314_U2205 ( .A1(div_divisor_0_), .A2(
        div_n302), .A3(div_n_T_51_64_), .Y(div_DP_OP_279J39_124_314_n2589) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2204 ( .A(div_DP_OP_279J39_124_314_n551), .B(div_DP_OP_279J39_124_314_n1646), .CI(div_DP_OP_279J39_124_314_n1648), .S(
        div_n_T_65[2]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2203 ( .A1(
        div_DP_OP_279J39_124_314_n1646), .A2(div_DP_OP_279J39_124_314_n1648), 
        .Y(div_DP_OP_279J39_124_314_n2784) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2202 ( .A1(
        div_DP_OP_279J39_124_314_n1646), .A2(div_DP_OP_279J39_124_314_n1648), 
        .Y(div_DP_OP_279J39_124_314_n2785) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2201 ( .A1(
        div_DP_OP_279J39_124_314_n551), .A2(div_DP_OP_279J39_124_314_n2784), 
        .A3(div_DP_OP_279J39_124_314_n2785), .Y(div_DP_OP_279J39_124_314_n2786) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2200 ( .A(
        div_DP_OP_279J39_124_314_n1645), .B(div_DP_OP_279J39_124_314_n1640), 
        .CI(div_DP_OP_279J39_124_314_n2786), .S(div_n_T_65[3]) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2199 ( .A(
        div_DP_OP_279J39_124_314_n2778), .B(div_DP_OP_279J39_124_314_n1639), 
        .CI(div_DP_OP_279J39_124_314_n1632), .S(div_n_T_65[4]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2198 ( .A1(
        div_DP_OP_279J39_124_314_n1639), .A2(div_DP_OP_279J39_124_314_n1632), 
        .Y(div_DP_OP_279J39_124_314_n2782) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2197 ( .A1(
        div_DP_OP_279J39_124_314_n2778), .A2(div_DP_OP_279J39_124_314_n2782), 
        .A3(div_DP_OP_279J39_124_314_n1639), .A4(
        div_DP_OP_279J39_124_314_n1632), .Y(div_DP_OP_279J39_124_314_n2783) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2196 ( .A(
        div_DP_OP_279J39_124_314_n1631), .B(div_DP_OP_279J39_124_314_n1622), 
        .CI(div_DP_OP_279J39_124_314_n2783), .S(div_n_T_65[5]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2195 ( .A1(
        div_DP_OP_279J39_124_314_n1639), .A2(div_DP_OP_279J39_124_314_n1632), 
        .A3(div_DP_OP_279J39_124_314_n1631), .A4(
        div_DP_OP_279J39_124_314_n1622), .Y(div_DP_OP_279J39_124_314_n2779) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2194 ( .A1(
        div_DP_OP_279J39_124_314_n2779), .A2(div_DP_OP_279J39_124_314_n2778), 
        .A3(div_DP_OP_279J39_124_314_n2776), .Y(div_DP_OP_279J39_124_314_n2781) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2193 ( .A(
        div_DP_OP_279J39_124_314_n1621), .B(div_DP_OP_279J39_124_314_n1610), 
        .CI(div_DP_OP_279J39_124_314_n2781), .S(div_n_T_65[6]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2192 ( .A1(
        div_DP_OP_279J39_124_314_n1621), .A2(div_DP_OP_279J39_124_314_n1610), 
        .Y(div_DP_OP_279J39_124_314_n2777) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2191 ( .A1(
        div_DP_OP_279J39_124_314_n2781), .A2(div_DP_OP_279J39_124_314_n1621), 
        .A3(div_DP_OP_279J39_124_314_n2781), .A4(
        div_DP_OP_279J39_124_314_n1610), .A5(div_DP_OP_279J39_124_314_n2777), 
        .Y(div_DP_OP_279J39_124_314_n2780) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2190 ( .A(
        div_DP_OP_279J39_124_314_n1609), .B(div_DP_OP_279J39_124_314_n1596), 
        .CI(div_DP_OP_279J39_124_314_n2780), .S(div_n_T_65[7]) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2189 ( .A(
        div_DP_OP_279J39_124_314_n1580), .B(div_DP_OP_279J39_124_314_n1595), 
        .CI(div_DP_OP_279J39_124_314_n2757), .S(div_n_T_65[8]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2188 ( .A1(
        div_DP_OP_279J39_124_314_n1580), .A2(div_DP_OP_279J39_124_314_n1595), 
        .Y(div_DP_OP_279J39_124_314_n2774) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2187 ( .A1(
        div_DP_OP_279J39_124_314_n2757), .A2(div_DP_OP_279J39_124_314_n1580), 
        .A3(div_DP_OP_279J39_124_314_n2757), .A4(
        div_DP_OP_279J39_124_314_n1595), .A5(div_DP_OP_279J39_124_314_n2774), 
        .Y(div_DP_OP_279J39_124_314_n2775) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2186 ( .A(
        div_DP_OP_279J39_124_314_n1579), .B(div_DP_OP_279J39_124_314_n1564), 
        .CI(div_DP_OP_279J39_124_314_n2775), .S(div_n_T_65[9]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2185 ( .A1(
        div_DP_OP_279J39_124_314_n1579), .A2(div_DP_OP_279J39_124_314_n1564), 
        .A3(div_DP_OP_279J39_124_314_n1580), .A4(
        div_DP_OP_279J39_124_314_n1595), .Y(div_DP_OP_279J39_124_314_n2771) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2184 ( .A1(
        div_DP_OP_279J39_124_314_n2771), .A2(div_DP_OP_279J39_124_314_n2757), 
        .A3(div_DP_OP_279J39_124_314_n2770), .Y(div_DP_OP_279J39_124_314_n2773) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2183 ( .A(
        div_DP_OP_279J39_124_314_n1548), .B(div_DP_OP_279J39_124_314_n1563), 
        .CI(div_DP_OP_279J39_124_314_n2773), .S(div_n_T_65[10]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2182 ( .A1(
        div_DP_OP_279J39_124_314_n1548), .A2(div_DP_OP_279J39_124_314_n1563), 
        .Y(div_DP_OP_279J39_124_314_n2767) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2181 ( .A1(
        div_DP_OP_279J39_124_314_n2767), .A2(div_DP_OP_279J39_124_314_n2773), 
        .A3(div_DP_OP_279J39_124_314_n1548), .A4(
        div_DP_OP_279J39_124_314_n1563), .Y(div_DP_OP_279J39_124_314_n2772) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2180 ( .A(
        div_DP_OP_279J39_124_314_n1547), .B(div_DP_OP_279J39_124_314_n1532), 
        .CI(div_DP_OP_279J39_124_314_n2772), .S(div_n_T_65[11]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2179 ( .A1(
        div_DP_OP_279J39_124_314_n1547), .A2(div_DP_OP_279J39_124_314_n1532), 
        .A3(div_DP_OP_279J39_124_314_n1548), .A4(
        div_DP_OP_279J39_124_314_n1563), .Y(div_DP_OP_279J39_124_314_n2769) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2178 ( .A1(
        div_DP_OP_279J39_124_314_n2769), .A2(div_DP_OP_279J39_124_314_n2771), 
        .Y(div_DP_OP_279J39_124_314_n2756) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2177 ( .A1(
        div_DP_OP_279J39_124_314_n1532), .A2(div_DP_OP_279J39_124_314_n1547), 
        .Y(div_DP_OP_279J39_124_314_n2768) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2176 ( .A1(
        div_DP_OP_279J39_124_314_n1547), .A2(div_DP_OP_279J39_124_314_n1532), 
        .A3(div_DP_OP_279J39_124_314_n2767), .A4(
        div_DP_OP_279J39_124_314_n2768), .A5(div_DP_OP_279J39_124_314_n2769), 
        .A6(div_DP_OP_279J39_124_314_n2770), .Y(div_DP_OP_279J39_124_314_n2759) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2175 ( .A1(
        div_DP_OP_279J39_124_314_n2756), .A2(div_DP_OP_279J39_124_314_n2757), 
        .A3(div_DP_OP_279J39_124_314_n2759), .Y(div_DP_OP_279J39_124_314_n2764) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2174 ( .A(
        div_DP_OP_279J39_124_314_n1531), .B(div_DP_OP_279J39_124_314_n1516), 
        .CI(div_DP_OP_279J39_124_314_n2764), .S(div_n_T_65[12]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2173 ( .A1(
        div_DP_OP_279J39_124_314_n1531), .A2(div_DP_OP_279J39_124_314_n1516), 
        .Y(div_DP_OP_279J39_124_314_n2765) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2172 ( .A1(
        div_DP_OP_279J39_124_314_n2765), .A2(div_DP_OP_279J39_124_314_n2764), 
        .A3(div_DP_OP_279J39_124_314_n1531), .A4(
        div_DP_OP_279J39_124_314_n1516), .Y(div_DP_OP_279J39_124_314_n2766) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2171 ( .A(
        div_DP_OP_279J39_124_314_n1515), .B(div_DP_OP_279J39_124_314_n1500), 
        .CI(div_DP_OP_279J39_124_314_n2766), .S(div_n_T_65[13]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2170 ( .A1(
        div_DP_OP_279J39_124_314_n1515), .A2(div_DP_OP_279J39_124_314_n1500), 
        .A3(div_DP_OP_279J39_124_314_n1531), .A4(
        div_DP_OP_279J39_124_314_n1516), .Y(div_DP_OP_279J39_124_314_n2761) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2169 ( .A1(
        div_DP_OP_279J39_124_314_n2761), .A2(div_DP_OP_279J39_124_314_n2764), 
        .A3(div_DP_OP_279J39_124_314_n2758), .Y(div_DP_OP_279J39_124_314_n2763) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2168 ( .A(
        div_DP_OP_279J39_124_314_n1499), .B(div_DP_OP_279J39_124_314_n1484), 
        .CI(div_DP_OP_279J39_124_314_n2763), .S(div_n_T_65[14]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2167 ( .A1(
        div_DP_OP_279J39_124_314_n1499), .A2(div_DP_OP_279J39_124_314_n1484), 
        .Y(div_DP_OP_279J39_124_314_n2760) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2166 ( .A1(
        div_DP_OP_279J39_124_314_n2760), .A2(div_DP_OP_279J39_124_314_n2763), 
        .A3(div_DP_OP_279J39_124_314_n1499), .A4(
        div_DP_OP_279J39_124_314_n1484), .Y(div_DP_OP_279J39_124_314_n2762) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2165 ( .A(
        div_DP_OP_279J39_124_314_n1483), .B(div_DP_OP_279J39_124_314_n1468), 
        .CI(div_DP_OP_279J39_124_314_n2762), .S(div_n_T_65[15]) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2164 ( .A(
        div_DP_OP_279J39_124_314_n2716), .B(div_DP_OP_279J39_124_314_n1467), 
        .CI(div_DP_OP_279J39_124_314_n1452), .S(div_n_T_65[16]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2163 ( .A1(
        div_DP_OP_279J39_124_314_n1467), .A2(div_DP_OP_279J39_124_314_n1452), 
        .Y(div_DP_OP_279J39_124_314_n2754) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2162 ( .A1(
        div_DP_OP_279J39_124_314_n2716), .A2(div_DP_OP_279J39_124_314_n2754), 
        .A3(div_DP_OP_279J39_124_314_n1467), .A4(
        div_DP_OP_279J39_124_314_n1452), .Y(div_DP_OP_279J39_124_314_n2755) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2161 ( .A(
        div_DP_OP_279J39_124_314_n1451), .B(div_DP_OP_279J39_124_314_n1436), 
        .CI(div_DP_OP_279J39_124_314_n2755), .S(div_n_T_65[17]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2160 ( .A1(
        div_DP_OP_279J39_124_314_n1451), .A2(div_DP_OP_279J39_124_314_n1436), 
        .A3(div_DP_OP_279J39_124_314_n1467), .A4(
        div_DP_OP_279J39_124_314_n1452), .Y(div_DP_OP_279J39_124_314_n2751) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2159 ( .A1(
        div_DP_OP_279J39_124_314_n2751), .A2(div_DP_OP_279J39_124_314_n2716), 
        .A3(div_DP_OP_279J39_124_314_n2750), .Y(div_DP_OP_279J39_124_314_n2753) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2158 ( .A(
        div_DP_OP_279J39_124_314_n1435), .B(div_DP_OP_279J39_124_314_n1420), 
        .CI(div_DP_OP_279J39_124_314_n2753), .S(div_n_T_65[18]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2157 ( .A1(
        div_DP_OP_279J39_124_314_n1435), .A2(div_DP_OP_279J39_124_314_n1420), 
        .Y(div_DP_OP_279J39_124_314_n2747) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2156 ( .A1(
        div_DP_OP_279J39_124_314_n2753), .A2(div_DP_OP_279J39_124_314_n1435), 
        .A3(div_DP_OP_279J39_124_314_n2753), .A4(
        div_DP_OP_279J39_124_314_n1420), .A5(div_DP_OP_279J39_124_314_n2747), 
        .Y(div_DP_OP_279J39_124_314_n2752) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2155 ( .A(
        div_DP_OP_279J39_124_314_n1419), .B(div_DP_OP_279J39_124_314_n1404), 
        .CI(div_DP_OP_279J39_124_314_n2752), .S(div_n_T_65[19]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2154 ( .A1(
        div_DP_OP_279J39_124_314_n1419), .A2(div_DP_OP_279J39_124_314_n1404), 
        .A3(div_DP_OP_279J39_124_314_n1435), .A4(
        div_DP_OP_279J39_124_314_n1420), .Y(div_DP_OP_279J39_124_314_n2749) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2153 ( .A1(
        div_DP_OP_279J39_124_314_n2749), .A2(div_DP_OP_279J39_124_314_n2751), 
        .Y(div_DP_OP_279J39_124_314_n2740) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2152 ( .A1(
        div_DP_OP_279J39_124_314_n1404), .A2(div_DP_OP_279J39_124_314_n1419), 
        .Y(div_DP_OP_279J39_124_314_n2748) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2151 ( .A1(
        div_DP_OP_279J39_124_314_n1419), .A2(div_DP_OP_279J39_124_314_n1404), 
        .A3(div_DP_OP_279J39_124_314_n2747), .A4(
        div_DP_OP_279J39_124_314_n2748), .A5(div_DP_OP_279J39_124_314_n2749), 
        .A6(div_DP_OP_279J39_124_314_n2750), .Y(div_DP_OP_279J39_124_314_n2737) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2150 ( .A1(
        div_DP_OP_279J39_124_314_n2716), .A2(div_DP_OP_279J39_124_314_n2740), 
        .A3(div_DP_OP_279J39_124_314_n2737), .Y(div_DP_OP_279J39_124_314_n2744) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2149 ( .A(
        div_DP_OP_279J39_124_314_n1403), .B(div_DP_OP_279J39_124_314_n1388), 
        .CI(div_DP_OP_279J39_124_314_n2744), .S(div_n_T_65[20]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2148 ( .A1(
        div_DP_OP_279J39_124_314_n1403), .A2(div_DP_OP_279J39_124_314_n1388), 
        .Y(div_DP_OP_279J39_124_314_n2745) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2147 ( .A1(
        div_DP_OP_279J39_124_314_n2744), .A2(div_DP_OP_279J39_124_314_n1403), 
        .A3(div_DP_OP_279J39_124_314_n2744), .A4(
        div_DP_OP_279J39_124_314_n1388), .A5(div_DP_OP_279J39_124_314_n2745), 
        .Y(div_DP_OP_279J39_124_314_n2746) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2146 ( .A(
        div_DP_OP_279J39_124_314_n1387), .B(div_DP_OP_279J39_124_314_n1372), 
        .CI(div_DP_OP_279J39_124_314_n2746), .S(div_n_T_65[21]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2145 ( .A1(
        div_DP_OP_279J39_124_314_n1387), .A2(div_DP_OP_279J39_124_314_n1372), 
        .A3(div_DP_OP_279J39_124_314_n1403), .A4(
        div_DP_OP_279J39_124_314_n1388), .Y(div_DP_OP_279J39_124_314_n2741) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2144 ( .A1(
        div_DP_OP_279J39_124_314_n2741), .A2(div_DP_OP_279J39_124_314_n2744), 
        .A3(div_DP_OP_279J39_124_314_n2736), .Y(div_DP_OP_279J39_124_314_n2743) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2143 ( .A(
        div_DP_OP_279J39_124_314_n1371), .B(div_DP_OP_279J39_124_314_n1356), 
        .CI(div_DP_OP_279J39_124_314_n2743), .S(div_n_T_65[22]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2142 ( .A1(
        div_DP_OP_279J39_124_314_n1371), .A2(div_DP_OP_279J39_124_314_n1356), 
        .Y(div_DP_OP_279J39_124_314_n2739) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2141 ( .A1(
        div_DP_OP_279J39_124_314_n2743), .A2(div_DP_OP_279J39_124_314_n1371), 
        .A3(div_DP_OP_279J39_124_314_n2743), .A4(
        div_DP_OP_279J39_124_314_n1356), .A5(div_DP_OP_279J39_124_314_n2739), 
        .Y(div_DP_OP_279J39_124_314_n2742) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2140 ( .A(
        div_DP_OP_279J39_124_314_n1355), .B(div_DP_OP_279J39_124_314_n1340), 
        .CI(div_DP_OP_279J39_124_314_n2742), .S(div_n_T_65[23]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2139 ( .A1(
        div_DP_OP_279J39_124_314_n1355), .A2(div_DP_OP_279J39_124_314_n1340), 
        .A3(div_DP_OP_279J39_124_314_n1371), .A4(
        div_DP_OP_279J39_124_314_n1356), .Y(div_DP_OP_279J39_124_314_n2735) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2138 ( .A1(
        div_DP_OP_279J39_124_314_n2735), .A2(div_DP_OP_279J39_124_314_n2741), 
        .Y(div_DP_OP_279J39_124_314_n2738) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2137 ( .A1(
        div_DP_OP_279J39_124_314_n2740), .A2(div_DP_OP_279J39_124_314_n2738), 
        .Y(div_DP_OP_279J39_124_314_n2717) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2136 ( .A1(
        div_DP_OP_279J39_124_314_n2717), .A2(div_DP_OP_279J39_124_314_n2716), 
        .A3(div_DP_OP_279J39_124_314_n2712), .Y(div_DP_OP_279J39_124_314_n2725) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2135 ( .A(
        div_DP_OP_279J39_124_314_n1339), .B(div_DP_OP_279J39_124_314_n1324), 
        .CI(div_DP_OP_279J39_124_314_n2725), .S(div_n_T_65[24]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2134 ( .A1(
        div_DP_OP_279J39_124_314_n1339), .A2(div_DP_OP_279J39_124_314_n1324), 
        .Y(div_DP_OP_279J39_124_314_n2733) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2133 ( .A1(
        div_DP_OP_279J39_124_314_n2725), .A2(div_DP_OP_279J39_124_314_n1339), 
        .A3(div_DP_OP_279J39_124_314_n2725), .A4(
        div_DP_OP_279J39_124_314_n1324), .A5(div_DP_OP_279J39_124_314_n2733), 
        .Y(div_DP_OP_279J39_124_314_n2734) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2132 ( .A(
        div_DP_OP_279J39_124_314_n1323), .B(div_DP_OP_279J39_124_314_n1308), 
        .CI(div_DP_OP_279J39_124_314_n2734), .S(div_n_T_65[25]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2131 ( .A1(
        div_DP_OP_279J39_124_314_n1323), .A2(div_DP_OP_279J39_124_314_n1308), 
        .A3(div_DP_OP_279J39_124_314_n1339), .A4(
        div_DP_OP_279J39_124_314_n1324), .Y(div_DP_OP_279J39_124_314_n2730) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2130 ( .A1(
        div_DP_OP_279J39_124_314_n2730), .A2(div_DP_OP_279J39_124_314_n2725), 
        .A3(div_DP_OP_279J39_124_314_n2729), .Y(div_DP_OP_279J39_124_314_n2732) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2129 ( .A(
        div_DP_OP_279J39_124_314_n1307), .B(div_DP_OP_279J39_124_314_n1292), 
        .CI(div_DP_OP_279J39_124_314_n2732), .S(div_n_T_65[26]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2128 ( .A1(
        div_DP_OP_279J39_124_314_n1307), .A2(div_DP_OP_279J39_124_314_n1292), 
        .Y(div_DP_OP_279J39_124_314_n2726) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2127 ( .A1(
        div_DP_OP_279J39_124_314_n2732), .A2(div_DP_OP_279J39_124_314_n1307), 
        .A3(div_DP_OP_279J39_124_314_n2732), .A4(
        div_DP_OP_279J39_124_314_n1292), .A5(div_DP_OP_279J39_124_314_n2726), 
        .Y(div_DP_OP_279J39_124_314_n2731) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2126 ( .A(
        div_DP_OP_279J39_124_314_n1291), .B(div_DP_OP_279J39_124_314_n1276), 
        .CI(div_DP_OP_279J39_124_314_n2731), .S(div_n_T_65[27]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2125 ( .A1(
        div_DP_OP_279J39_124_314_n1291), .A2(div_DP_OP_279J39_124_314_n1276), 
        .A3(div_DP_OP_279J39_124_314_n1307), .A4(
        div_DP_OP_279J39_124_314_n1292), .Y(div_DP_OP_279J39_124_314_n2728) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2124 ( .A1(
        div_DP_OP_279J39_124_314_n2728), .A2(div_DP_OP_279J39_124_314_n2730), 
        .Y(div_DP_OP_279J39_124_314_n2718) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2123 ( .A1(
        div_DP_OP_279J39_124_314_n1276), .A2(div_DP_OP_279J39_124_314_n1291), 
        .Y(div_DP_OP_279J39_124_314_n2727) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2122 ( .A1(
        div_DP_OP_279J39_124_314_n1291), .A2(div_DP_OP_279J39_124_314_n1276), 
        .A3(div_DP_OP_279J39_124_314_n2726), .A4(
        div_DP_OP_279J39_124_314_n2727), .A5(div_DP_OP_279J39_124_314_n2728), 
        .A6(div_DP_OP_279J39_124_314_n2729), .Y(div_DP_OP_279J39_124_314_n2714) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2121 ( .A1(
        div_DP_OP_279J39_124_314_n2718), .A2(div_DP_OP_279J39_124_314_n2725), 
        .A3(div_DP_OP_279J39_124_314_n2714), .Y(div_DP_OP_279J39_124_314_n2722) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2120 ( .A(
        div_DP_OP_279J39_124_314_n1275), .B(div_DP_OP_279J39_124_314_n1260), 
        .CI(div_DP_OP_279J39_124_314_n2722), .S(div_n_T_65[28]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2119 ( .A1(
        div_DP_OP_279J39_124_314_n1275), .A2(div_DP_OP_279J39_124_314_n1260), 
        .Y(div_DP_OP_279J39_124_314_n2723) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2118 ( .A1(
        div_DP_OP_279J39_124_314_n2722), .A2(div_DP_OP_279J39_124_314_n1275), 
        .A3(div_DP_OP_279J39_124_314_n2722), .A4(
        div_DP_OP_279J39_124_314_n1260), .A5(div_DP_OP_279J39_124_314_n2723), 
        .Y(div_DP_OP_279J39_124_314_n2724) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2117 ( .A(
        div_DP_OP_279J39_124_314_n1259), .B(div_DP_OP_279J39_124_314_n1244), 
        .CI(div_DP_OP_279J39_124_314_n2724), .S(div_n_T_65[29]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2116 ( .A1(
        div_DP_OP_279J39_124_314_n1259), .A2(div_DP_OP_279J39_124_314_n1244), 
        .A3(div_DP_OP_279J39_124_314_n1275), .A4(
        div_DP_OP_279J39_124_314_n1260), .Y(div_DP_OP_279J39_124_314_n2719) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2115 ( .A1(
        div_DP_OP_279J39_124_314_n2719), .A2(div_DP_OP_279J39_124_314_n2722), 
        .A3(div_DP_OP_279J39_124_314_n2713), .Y(div_DP_OP_279J39_124_314_n2721) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2114 ( .A(
        div_DP_OP_279J39_124_314_n1243), .B(div_DP_OP_279J39_124_314_n1228), 
        .CI(div_DP_OP_279J39_124_314_n2721), .S(div_n_T_65[30]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2113 ( .A1(
        div_DP_OP_279J39_124_314_n1243), .A2(div_DP_OP_279J39_124_314_n1228), 
        .Y(div_DP_OP_279J39_124_314_n2715) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2112 ( .A1(
        div_DP_OP_279J39_124_314_n2721), .A2(div_DP_OP_279J39_124_314_n1243), 
        .A3(div_DP_OP_279J39_124_314_n2721), .A4(
        div_DP_OP_279J39_124_314_n1228), .A5(div_DP_OP_279J39_124_314_n2715), 
        .Y(div_DP_OP_279J39_124_314_n2720) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2111 ( .A(
        div_DP_OP_279J39_124_314_n1227), .B(div_DP_OP_279J39_124_314_n1212), 
        .CI(div_DP_OP_279J39_124_314_n2720), .S(div_n_T_65[31]) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2110 ( .A(
        div_DP_OP_279J39_124_314_n1211), .B(div_DP_OP_279J39_124_314_n1196), 
        .CI(div_DP_OP_279J39_124_314_n2618), .S(div_n_T_65[32]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2109 ( .A1(
        div_DP_OP_279J39_124_314_n1211), .A2(div_DP_OP_279J39_124_314_n1196), 
        .Y(div_DP_OP_279J39_124_314_n2710) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2108 ( .A1(
        div_DP_OP_279J39_124_314_n2618), .A2(div_DP_OP_279J39_124_314_n1211), 
        .A3(div_DP_OP_279J39_124_314_n2618), .A4(
        div_DP_OP_279J39_124_314_n1196), .A5(div_DP_OP_279J39_124_314_n2710), 
        .Y(div_DP_OP_279J39_124_314_n2711) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2107 ( .A(
        div_DP_OP_279J39_124_314_n1195), .B(div_DP_OP_279J39_124_314_n1180), 
        .CI(div_DP_OP_279J39_124_314_n2711), .S(div_n_T_65[33]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2106 ( .A1(
        div_DP_OP_279J39_124_314_n1195), .A2(div_DP_OP_279J39_124_314_n1180), 
        .A3(div_DP_OP_279J39_124_314_n1211), .A4(
        div_DP_OP_279J39_124_314_n1196), .Y(div_DP_OP_279J39_124_314_n2707) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2105 ( .A1(
        div_DP_OP_279J39_124_314_n2707), .A2(div_DP_OP_279J39_124_314_n2618), 
        .A3(div_DP_OP_279J39_124_314_n2706), .Y(div_DP_OP_279J39_124_314_n2709) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2104 ( .A(
        div_DP_OP_279J39_124_314_n1179), .B(div_DP_OP_279J39_124_314_n1164), 
        .CI(div_DP_OP_279J39_124_314_n2709), .S(div_n_T_65[34]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2103 ( .A1(
        div_DP_OP_279J39_124_314_n1179), .A2(div_DP_OP_279J39_124_314_n1164), 
        .Y(div_DP_OP_279J39_124_314_n2703) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2102 ( .A1(
        div_DP_OP_279J39_124_314_n2703), .A2(div_DP_OP_279J39_124_314_n2709), 
        .A3(div_DP_OP_279J39_124_314_n1179), .A4(
        div_DP_OP_279J39_124_314_n1164), .Y(div_DP_OP_279J39_124_314_n2708) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2101 ( .A(
        div_DP_OP_279J39_124_314_n1163), .B(div_DP_OP_279J39_124_314_n1148), 
        .CI(div_DP_OP_279J39_124_314_n2708), .S(div_n_T_65[35]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2100 ( .A1(
        div_DP_OP_279J39_124_314_n1163), .A2(div_DP_OP_279J39_124_314_n1148), 
        .A3(div_DP_OP_279J39_124_314_n1179), .A4(
        div_DP_OP_279J39_124_314_n1164), .Y(div_DP_OP_279J39_124_314_n2705) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2099 ( .A1(
        div_DP_OP_279J39_124_314_n2705), .A2(div_DP_OP_279J39_124_314_n2707), 
        .Y(div_DP_OP_279J39_124_314_n2696) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2098 ( .A1(
        div_DP_OP_279J39_124_314_n1148), .A2(div_DP_OP_279J39_124_314_n1163), 
        .Y(div_DP_OP_279J39_124_314_n2704) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2097 ( .A1(
        div_DP_OP_279J39_124_314_n1163), .A2(div_DP_OP_279J39_124_314_n1148), 
        .A3(div_DP_OP_279J39_124_314_n2703), .A4(
        div_DP_OP_279J39_124_314_n2704), .A5(div_DP_OP_279J39_124_314_n2705), 
        .A6(div_DP_OP_279J39_124_314_n2706), .Y(div_DP_OP_279J39_124_314_n2693) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2096 ( .A1(
        div_DP_OP_279J39_124_314_n2696), .A2(div_DP_OP_279J39_124_314_n2618), 
        .A3(div_DP_OP_279J39_124_314_n2693), .Y(div_DP_OP_279J39_124_314_n2700) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2095 ( .A(
        div_DP_OP_279J39_124_314_n1147), .B(div_DP_OP_279J39_124_314_n1132), 
        .CI(div_DP_OP_279J39_124_314_n2700), .S(div_n_T_65[36]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2094 ( .A1(
        div_DP_OP_279J39_124_314_n1147), .A2(div_DP_OP_279J39_124_314_n1132), 
        .Y(div_DP_OP_279J39_124_314_n2701) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2093 ( .A1(
        div_DP_OP_279J39_124_314_n2701), .A2(div_DP_OP_279J39_124_314_n2700), 
        .A3(div_DP_OP_279J39_124_314_n1147), .A4(
        div_DP_OP_279J39_124_314_n1132), .Y(div_DP_OP_279J39_124_314_n2702) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2092 ( .A(
        div_DP_OP_279J39_124_314_n1131), .B(div_DP_OP_279J39_124_314_n1116), 
        .CI(div_DP_OP_279J39_124_314_n2702), .S(div_n_T_65[37]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2091 ( .A1(
        div_DP_OP_279J39_124_314_n1131), .A2(div_DP_OP_279J39_124_314_n1116), 
        .A3(div_DP_OP_279J39_124_314_n1147), .A4(
        div_DP_OP_279J39_124_314_n1132), .Y(div_DP_OP_279J39_124_314_n2697) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2090 ( .A1(
        div_DP_OP_279J39_124_314_n2697), .A2(div_DP_OP_279J39_124_314_n2700), 
        .A3(div_DP_OP_279J39_124_314_n2692), .Y(div_DP_OP_279J39_124_314_n2699) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2089 ( .A(
        div_DP_OP_279J39_124_314_n1115), .B(div_DP_OP_279J39_124_314_n1100), 
        .CI(div_DP_OP_279J39_124_314_n2699), .S(div_n_T_65[38]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2088 ( .A1(
        div_DP_OP_279J39_124_314_n1115), .A2(div_DP_OP_279J39_124_314_n1100), 
        .Y(div_DP_OP_279J39_124_314_n2695) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2087 ( .A1(
        div_DP_OP_279J39_124_314_n2695), .A2(div_DP_OP_279J39_124_314_n2699), 
        .A3(div_DP_OP_279J39_124_314_n1115), .A4(
        div_DP_OP_279J39_124_314_n1100), .Y(div_DP_OP_279J39_124_314_n2698) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2086 ( .A(
        div_DP_OP_279J39_124_314_n1099), .B(div_DP_OP_279J39_124_314_n1084), 
        .CI(div_DP_OP_279J39_124_314_n2698), .S(div_n_T_65[39]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2085 ( .A1(
        div_DP_OP_279J39_124_314_n1099), .A2(div_DP_OP_279J39_124_314_n1084), 
        .A3(div_DP_OP_279J39_124_314_n1115), .A4(
        div_DP_OP_279J39_124_314_n1100), .Y(div_DP_OP_279J39_124_314_n2691) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2084 ( .A1(
        div_DP_OP_279J39_124_314_n2691), .A2(div_DP_OP_279J39_124_314_n2697), 
        .Y(div_DP_OP_279J39_124_314_n2694) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2083 ( .A1(
        div_DP_OP_279J39_124_314_n2694), .A2(div_DP_OP_279J39_124_314_n2696), 
        .Y(div_DP_OP_279J39_124_314_n2673) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2082 ( .A1(
        div_DP_OP_279J39_124_314_n2673), .A2(div_DP_OP_279J39_124_314_n2618), 
        .A3(div_DP_OP_279J39_124_314_n2667), .Y(div_DP_OP_279J39_124_314_n2681) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2081 ( .A(
        div_DP_OP_279J39_124_314_n1083), .B(div_DP_OP_279J39_124_314_n1068), 
        .CI(div_DP_OP_279J39_124_314_n2681), .S(div_n_T_65[40]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2080 ( .A1(
        div_DP_OP_279J39_124_314_n1083), .A2(div_DP_OP_279J39_124_314_n1068), 
        .Y(div_DP_OP_279J39_124_314_n2689) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2079 ( .A1(
        div_DP_OP_279J39_124_314_n2689), .A2(div_DP_OP_279J39_124_314_n2681), 
        .A3(div_DP_OP_279J39_124_314_n1083), .A4(
        div_DP_OP_279J39_124_314_n1068), .Y(div_DP_OP_279J39_124_314_n2690) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2078 ( .A(
        div_DP_OP_279J39_124_314_n1067), .B(div_DP_OP_279J39_124_314_n1052), 
        .CI(div_DP_OP_279J39_124_314_n2690), .S(div_n_T_65[41]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2077 ( .A1(
        div_DP_OP_279J39_124_314_n1067), .A2(div_DP_OP_279J39_124_314_n1052), 
        .A3(div_DP_OP_279J39_124_314_n1083), .A4(
        div_DP_OP_279J39_124_314_n1068), .Y(div_DP_OP_279J39_124_314_n2686) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2076 ( .A1(
        div_DP_OP_279J39_124_314_n2686), .A2(div_DP_OP_279J39_124_314_n2681), 
        .A3(div_DP_OP_279J39_124_314_n2685), .Y(div_DP_OP_279J39_124_314_n2688) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2075 ( .A(
        div_DP_OP_279J39_124_314_n1051), .B(div_DP_OP_279J39_124_314_n1036), 
        .CI(div_DP_OP_279J39_124_314_n2688), .S(div_n_T_65[42]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2074 ( .A1(
        div_DP_OP_279J39_124_314_n1051), .A2(div_DP_OP_279J39_124_314_n1036), 
        .Y(div_DP_OP_279J39_124_314_n2682) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2073 ( .A1(
        div_DP_OP_279J39_124_314_n2682), .A2(div_DP_OP_279J39_124_314_n2688), 
        .A3(div_DP_OP_279J39_124_314_n1051), .A4(
        div_DP_OP_279J39_124_314_n1036), .Y(div_DP_OP_279J39_124_314_n2687) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2072 ( .A(
        div_DP_OP_279J39_124_314_n1035), .B(div_DP_OP_279J39_124_314_n1020), 
        .CI(div_DP_OP_279J39_124_314_n2687), .S(div_n_T_65[43]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2071 ( .A1(
        div_DP_OP_279J39_124_314_n1035), .A2(div_DP_OP_279J39_124_314_n1020), 
        .A3(div_DP_OP_279J39_124_314_n1051), .A4(
        div_DP_OP_279J39_124_314_n1036), .Y(div_DP_OP_279J39_124_314_n2684) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2070 ( .A1(
        div_DP_OP_279J39_124_314_n2684), .A2(div_DP_OP_279J39_124_314_n2686), 
        .Y(div_DP_OP_279J39_124_314_n2674) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2069 ( .A1(
        div_DP_OP_279J39_124_314_n1020), .A2(div_DP_OP_279J39_124_314_n1035), 
        .Y(div_DP_OP_279J39_124_314_n2683) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2068 ( .A1(
        div_DP_OP_279J39_124_314_n1035), .A2(div_DP_OP_279J39_124_314_n1020), 
        .A3(div_DP_OP_279J39_124_314_n2682), .A4(
        div_DP_OP_279J39_124_314_n2683), .A5(div_DP_OP_279J39_124_314_n2684), 
        .A6(div_DP_OP_279J39_124_314_n2685), .Y(div_DP_OP_279J39_124_314_n2664) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2067 ( .A1(
        div_DP_OP_279J39_124_314_n2674), .A2(div_DP_OP_279J39_124_314_n2681), 
        .A3(div_DP_OP_279J39_124_314_n2664), .Y(div_DP_OP_279J39_124_314_n2678) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2066 ( .A(
        div_DP_OP_279J39_124_314_n1019), .B(div_DP_OP_279J39_124_314_n1004), 
        .CI(div_DP_OP_279J39_124_314_n2678), .S(div_n_T_65[44]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2065 ( .A1(
        div_DP_OP_279J39_124_314_n1019), .A2(div_DP_OP_279J39_124_314_n1004), 
        .Y(div_DP_OP_279J39_124_314_n2679) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2064 ( .A1(
        div_DP_OP_279J39_124_314_n2679), .A2(div_DP_OP_279J39_124_314_n2678), 
        .A3(div_DP_OP_279J39_124_314_n1019), .A4(
        div_DP_OP_279J39_124_314_n1004), .Y(div_DP_OP_279J39_124_314_n2680) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2063 ( .A(
        div_DP_OP_279J39_124_314_n1003), .B(div_DP_OP_279J39_124_314_n988), 
        .CI(div_DP_OP_279J39_124_314_n2680), .S(div_n_T_65[45]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2062 ( .A1(
        div_DP_OP_279J39_124_314_n1003), .A2(div_DP_OP_279J39_124_314_n988), 
        .A3(div_DP_OP_279J39_124_314_n1019), .A4(
        div_DP_OP_279J39_124_314_n1004), .Y(div_DP_OP_279J39_124_314_n2675) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2061 ( .A1(
        div_DP_OP_279J39_124_314_n2675), .A2(div_DP_OP_279J39_124_314_n2678), 
        .A3(div_DP_OP_279J39_124_314_n2672), .Y(div_DP_OP_279J39_124_314_n2677) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2060 ( .A(div_DP_OP_279J39_124_314_n987), .B(div_DP_OP_279J39_124_314_n972), .CI(div_DP_OP_279J39_124_314_n2677), .S(
        div_n_T_65[46]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2059 ( .A1(
        div_DP_OP_279J39_124_314_n987), .A2(div_DP_OP_279J39_124_314_n972), 
        .Y(div_DP_OP_279J39_124_314_n2669) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2058 ( .A1(
        div_DP_OP_279J39_124_314_n2669), .A2(div_DP_OP_279J39_124_314_n2677), 
        .A3(div_DP_OP_279J39_124_314_n987), .A4(div_DP_OP_279J39_124_314_n972), 
        .Y(div_DP_OP_279J39_124_314_n2676) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2057 ( .A(div_DP_OP_279J39_124_314_n971), .B(div_DP_OP_279J39_124_314_n956), .CI(div_DP_OP_279J39_124_314_n2676), .S(
        div_n_T_65[47]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2056 ( .A1(
        div_DP_OP_279J39_124_314_n971), .A2(div_DP_OP_279J39_124_314_n956), 
        .A3(div_DP_OP_279J39_124_314_n987), .A4(div_DP_OP_279J39_124_314_n972), 
        .Y(div_DP_OP_279J39_124_314_n2671) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2055 ( .A1(
        div_DP_OP_279J39_124_314_n2671), .A2(div_DP_OP_279J39_124_314_n2675), 
        .Y(div_DP_OP_279J39_124_314_n2665) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2054 ( .A1(
        div_DP_OP_279J39_124_314_n2674), .A2(div_DP_OP_279J39_124_314_n2665), 
        .Y(div_DP_OP_279J39_124_314_n2666) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2053 ( .A1(
        div_DP_OP_279J39_124_314_n2666), .A2(div_DP_OP_279J39_124_314_n2673), 
        .Y(div_DP_OP_279J39_124_314_n2617) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2052 ( .A1(div_DP_OP_279J39_124_314_n956), .A2(div_DP_OP_279J39_124_314_n971), .Y(div_DP_OP_279J39_124_314_n2670) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2051 ( .A1(
        div_DP_OP_279J39_124_314_n971), .A2(div_DP_OP_279J39_124_314_n956), 
        .A3(div_DP_OP_279J39_124_314_n2669), .A4(
        div_DP_OP_279J39_124_314_n2670), .A5(div_DP_OP_279J39_124_314_n2671), 
        .A6(div_DP_OP_279J39_124_314_n2672), .Y(div_DP_OP_279J39_124_314_n2668) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2050 ( .A1(
        div_DP_OP_279J39_124_314_n2664), .A2(div_DP_OP_279J39_124_314_n2665), 
        .A3(div_DP_OP_279J39_124_314_n2666), .A4(
        div_DP_OP_279J39_124_314_n2667), .A5(div_DP_OP_279J39_124_314_n2668), 
        .Y(div_DP_OP_279J39_124_314_n2619) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2049 ( .A1(
        div_DP_OP_279J39_124_314_n2617), .A2(div_DP_OP_279J39_124_314_n2618), 
        .A3(div_DP_OP_279J39_124_314_n2619), .Y(div_DP_OP_279J39_124_314_n2642) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2048 ( .A(div_DP_OP_279J39_124_314_n955), .B(div_DP_OP_279J39_124_314_n940), .CI(div_DP_OP_279J39_124_314_n2642), .S(
        div_n_T_65[48]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2047 ( .A1(
        div_DP_OP_279J39_124_314_n955), .A2(div_DP_OP_279J39_124_314_n940), 
        .Y(div_DP_OP_279J39_124_314_n2662) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2046 ( .A1(
        div_DP_OP_279J39_124_314_n2662), .A2(div_DP_OP_279J39_124_314_n2642), 
        .A3(div_DP_OP_279J39_124_314_n955), .A4(div_DP_OP_279J39_124_314_n940), 
        .Y(div_DP_OP_279J39_124_314_n2663) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2045 ( .A(div_DP_OP_279J39_124_314_n939), .B(div_DP_OP_279J39_124_314_n924), .CI(div_DP_OP_279J39_124_314_n2663), .S(
        div_n_T_65[49]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2044 ( .A1(
        div_DP_OP_279J39_124_314_n939), .A2(div_DP_OP_279J39_124_314_n924), 
        .A3(div_DP_OP_279J39_124_314_n955), .A4(div_DP_OP_279J39_124_314_n940), 
        .Y(div_DP_OP_279J39_124_314_n2659) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2043 ( .A1(
        div_DP_OP_279J39_124_314_n2659), .A2(div_DP_OP_279J39_124_314_n2642), 
        .A3(div_DP_OP_279J39_124_314_n2658), .Y(div_DP_OP_279J39_124_314_n2661) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2042 ( .A(div_DP_OP_279J39_124_314_n923), .B(div_DP_OP_279J39_124_314_n908), .CI(div_DP_OP_279J39_124_314_n2661), .S(
        div_n_T_65[50]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2041 ( .A1(
        div_DP_OP_279J39_124_314_n923), .A2(div_DP_OP_279J39_124_314_n908), 
        .Y(div_DP_OP_279J39_124_314_n2655) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2040 ( .A1(
        div_DP_OP_279J39_124_314_n2655), .A2(div_DP_OP_279J39_124_314_n2661), 
        .A3(div_DP_OP_279J39_124_314_n923), .A4(div_DP_OP_279J39_124_314_n908), 
        .Y(div_DP_OP_279J39_124_314_n2660) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2039 ( .A(div_DP_OP_279J39_124_314_n907), .B(div_DP_OP_279J39_124_314_n892), .CI(div_DP_OP_279J39_124_314_n2660), .S(
        div_n_T_65[51]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2038 ( .A1(
        div_DP_OP_279J39_124_314_n907), .A2(div_DP_OP_279J39_124_314_n892), 
        .A3(div_DP_OP_279J39_124_314_n923), .A4(div_DP_OP_279J39_124_314_n908), 
        .Y(div_DP_OP_279J39_124_314_n2657) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2037 ( .A1(
        div_DP_OP_279J39_124_314_n2657), .A2(div_DP_OP_279J39_124_314_n2659), 
        .Y(div_DP_OP_279J39_124_314_n2648) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2036 ( .A1(div_DP_OP_279J39_124_314_n892), .A2(div_DP_OP_279J39_124_314_n907), .Y(div_DP_OP_279J39_124_314_n2656) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2035 ( .A1(
        div_DP_OP_279J39_124_314_n907), .A2(div_DP_OP_279J39_124_314_n892), 
        .A3(div_DP_OP_279J39_124_314_n2655), .A4(
        div_DP_OP_279J39_124_314_n2656), .A5(div_DP_OP_279J39_124_314_n2657), 
        .A6(div_DP_OP_279J39_124_314_n2658), .Y(div_DP_OP_279J39_124_314_n2645) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2034 ( .A1(
        div_DP_OP_279J39_124_314_n2648), .A2(div_DP_OP_279J39_124_314_n2642), 
        .A3(div_DP_OP_279J39_124_314_n2645), .Y(div_DP_OP_279J39_124_314_n2652) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2033 ( .A(div_DP_OP_279J39_124_314_n891), .B(div_DP_OP_279J39_124_314_n876), .CI(div_DP_OP_279J39_124_314_n2652), .S(
        div_n_T_65[52]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2032 ( .A1(
        div_DP_OP_279J39_124_314_n891), .A2(div_DP_OP_279J39_124_314_n876), 
        .Y(div_DP_OP_279J39_124_314_n2653) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2031 ( .A1(
        div_DP_OP_279J39_124_314_n2653), .A2(div_DP_OP_279J39_124_314_n2652), 
        .A3(div_DP_OP_279J39_124_314_n891), .A4(div_DP_OP_279J39_124_314_n876), 
        .Y(div_DP_OP_279J39_124_314_n2654) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2030 ( .A(div_DP_OP_279J39_124_314_n875), .B(div_DP_OP_279J39_124_314_n860), .CI(div_DP_OP_279J39_124_314_n2654), .S(
        div_n_T_65[53]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2029 ( .A1(
        div_DP_OP_279J39_124_314_n875), .A2(div_DP_OP_279J39_124_314_n860), 
        .A3(div_DP_OP_279J39_124_314_n891), .A4(div_DP_OP_279J39_124_314_n876), 
        .Y(div_DP_OP_279J39_124_314_n2649) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2028 ( .A1(
        div_DP_OP_279J39_124_314_n2649), .A2(div_DP_OP_279J39_124_314_n2652), 
        .A3(div_DP_OP_279J39_124_314_n2644), .Y(div_DP_OP_279J39_124_314_n2651) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2027 ( .A(div_DP_OP_279J39_124_314_n859), .B(div_DP_OP_279J39_124_314_n844), .CI(div_DP_OP_279J39_124_314_n2651), .S(
        div_n_T_65[54]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2026 ( .A1(
        div_DP_OP_279J39_124_314_n859), .A2(div_DP_OP_279J39_124_314_n844), 
        .Y(div_DP_OP_279J39_124_314_n2647) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2025 ( .A1(
        div_DP_OP_279J39_124_314_n2647), .A2(div_DP_OP_279J39_124_314_n2651), 
        .A3(div_DP_OP_279J39_124_314_n859), .A4(div_DP_OP_279J39_124_314_n844), 
        .Y(div_DP_OP_279J39_124_314_n2650) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2024 ( .A(div_DP_OP_279J39_124_314_n843), .B(div_DP_OP_279J39_124_314_n828), .CI(div_DP_OP_279J39_124_314_n2650), .S(
        div_n_T_65[55]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2023 ( .A1(
        div_DP_OP_279J39_124_314_n843), .A2(div_DP_OP_279J39_124_314_n828), 
        .A3(div_DP_OP_279J39_124_314_n859), .A4(div_DP_OP_279J39_124_314_n844), 
        .Y(div_DP_OP_279J39_124_314_n2643) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2022 ( .A1(
        div_DP_OP_279J39_124_314_n2643), .A2(div_DP_OP_279J39_124_314_n2649), 
        .Y(div_DP_OP_279J39_124_314_n2646) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2021 ( .A1(
        div_DP_OP_279J39_124_314_n2646), .A2(div_DP_OP_279J39_124_314_n2648), 
        .Y(div_DP_OP_279J39_124_314_n2625) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2020 ( .A1(
        div_DP_OP_279J39_124_314_n2625), .A2(div_DP_OP_279J39_124_314_n2642), 
        .A3(div_DP_OP_279J39_124_314_n2620), .Y(div_DP_OP_279J39_124_314_n2632) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2019 ( .A(div_DP_OP_279J39_124_314_n827), .B(div_DP_OP_279J39_124_314_n812), .CI(div_DP_OP_279J39_124_314_n2632), .S(
        div_n_T_65[56]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2018 ( .A1(
        div_DP_OP_279J39_124_314_n827), .A2(div_DP_OP_279J39_124_314_n812), 
        .Y(div_DP_OP_279J39_124_314_n2640) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2017 ( .A1(
        div_DP_OP_279J39_124_314_n2640), .A2(div_DP_OP_279J39_124_314_n2632), 
        .A3(div_DP_OP_279J39_124_314_n827), .A4(div_DP_OP_279J39_124_314_n812), 
        .Y(div_DP_OP_279J39_124_314_n2641) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2016 ( .A(div_DP_OP_279J39_124_314_n811), .B(div_DP_OP_279J39_124_314_n796), .CI(div_DP_OP_279J39_124_314_n2641), .S(
        div_n_T_65[57]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2015 ( .A1(
        div_DP_OP_279J39_124_314_n811), .A2(div_DP_OP_279J39_124_314_n796), 
        .A3(div_DP_OP_279J39_124_314_n827), .A4(div_DP_OP_279J39_124_314_n812), 
        .Y(div_DP_OP_279J39_124_314_n2637) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2014 ( .A1(
        div_DP_OP_279J39_124_314_n2637), .A2(div_DP_OP_279J39_124_314_n2632), 
        .A3(div_DP_OP_279J39_124_314_n2636), .Y(div_DP_OP_279J39_124_314_n2639) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2013 ( .A(div_DP_OP_279J39_124_314_n795), .B(div_DP_OP_279J39_124_314_n780), .CI(div_DP_OP_279J39_124_314_n2639), .S(
        div_n_T_65[58]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2012 ( .A1(
        div_DP_OP_279J39_124_314_n795), .A2(div_DP_OP_279J39_124_314_n780), 
        .Y(div_DP_OP_279J39_124_314_n2633) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2011 ( .A1(
        div_DP_OP_279J39_124_314_n2633), .A2(div_DP_OP_279J39_124_314_n2639), 
        .A3(div_DP_OP_279J39_124_314_n795), .A4(div_DP_OP_279J39_124_314_n780), 
        .Y(div_DP_OP_279J39_124_314_n2638) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2010 ( .A(div_DP_OP_279J39_124_314_n779), .B(div_DP_OP_279J39_124_314_n764), .CI(div_DP_OP_279J39_124_314_n2638), .S(
        div_n_T_65[59]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2009 ( .A1(
        div_DP_OP_279J39_124_314_n779), .A2(div_DP_OP_279J39_124_314_n764), 
        .A3(div_DP_OP_279J39_124_314_n795), .A4(div_DP_OP_279J39_124_314_n780), 
        .Y(div_DP_OP_279J39_124_314_n2635) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2008 ( .A1(
        div_DP_OP_279J39_124_314_n2635), .A2(div_DP_OP_279J39_124_314_n2637), 
        .Y(div_DP_OP_279J39_124_314_n2626) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U2007 ( .A1(div_DP_OP_279J39_124_314_n764), .A2(div_DP_OP_279J39_124_314_n779), .Y(div_DP_OP_279J39_124_314_n2634) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U2006 ( .A1(
        div_DP_OP_279J39_124_314_n779), .A2(div_DP_OP_279J39_124_314_n764), 
        .A3(div_DP_OP_279J39_124_314_n2633), .A4(
        div_DP_OP_279J39_124_314_n2634), .A5(div_DP_OP_279J39_124_314_n2635), 
        .A6(div_DP_OP_279J39_124_314_n2636), .Y(div_DP_OP_279J39_124_314_n2624) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U2005 ( .A1(
        div_DP_OP_279J39_124_314_n2626), .A2(div_DP_OP_279J39_124_314_n2632), 
        .A3(div_DP_OP_279J39_124_314_n2624), .Y(div_DP_OP_279J39_124_314_n2629) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2004 ( .A(div_DP_OP_279J39_124_314_n763), .B(div_DP_OP_279J39_124_314_n748), .CI(div_DP_OP_279J39_124_314_n2629), .S(
        div_n_T_65[60]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U2003 ( .A1(
        div_DP_OP_279J39_124_314_n763), .A2(div_DP_OP_279J39_124_314_n748), 
        .Y(div_DP_OP_279J39_124_314_n2630) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U2002 ( .A1(
        div_DP_OP_279J39_124_314_n2629), .A2(div_DP_OP_279J39_124_314_n763), 
        .A3(div_DP_OP_279J39_124_314_n2629), .A4(div_DP_OP_279J39_124_314_n748), .A5(div_DP_OP_279J39_124_314_n2630), .Y(div_DP_OP_279J39_124_314_n2631) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U2001 ( .A(div_DP_OP_279J39_124_314_n747), .B(div_DP_OP_279J39_124_314_n732), .CI(div_DP_OP_279J39_124_314_n2631), .S(
        div_n_T_65[61]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U2000 ( .A1(
        div_DP_OP_279J39_124_314_n747), .A2(div_DP_OP_279J39_124_314_n732), 
        .A3(div_DP_OP_279J39_124_314_n763), .A4(div_DP_OP_279J39_124_314_n748), 
        .Y(div_DP_OP_279J39_124_314_n2623) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1999 ( .A1(
        div_DP_OP_279J39_124_314_n2623), .A2(div_DP_OP_279J39_124_314_n2629), 
        .A3(div_DP_OP_279J39_124_314_n2622), .Y(div_DP_OP_279J39_124_314_n2628) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1998 ( .A(div_DP_OP_279J39_124_314_n731), .B(div_DP_OP_279J39_124_314_n716), .CI(div_DP_OP_279J39_124_314_n2628), .S(
        div_n_T_65[62]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1997 ( .A1(div_DP_OP_279J39_124_314_n731), .A2(div_DP_OP_279J39_124_314_n716), .Y(div_DP_OP_279J39_124_314_n2621) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1996 ( .A1(
        div_DP_OP_279J39_124_314_n731), .A2(div_DP_OP_279J39_124_314_n716), 
        .A3(div_DP_OP_279J39_124_314_n2628), .A4(
        div_DP_OP_279J39_124_314_n2621), .Y(div_DP_OP_279J39_124_314_n2627) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1995 ( .A(div_DP_OP_279J39_124_314_n715), .B(div_DP_OP_279J39_124_314_n700), .CI(div_DP_OP_279J39_124_314_n2627), .S(
        div_n_T_65[63]) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1994 ( .A(div_DP_OP_279J39_124_314_n699), .B(div_DP_OP_279J39_124_314_n684), .CI(div_DP_OP_279J39_124_314_n2594), .S(
        div_n_T_65[64]) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U1993 ( .A1(
        div_DP_OP_279J39_124_314_n699), .A2(div_DP_OP_279J39_124_314_n684), 
        .Y(div_DP_OP_279J39_124_314_n2615) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U1992 ( .A1(
        div_DP_OP_279J39_124_314_n699), .A2(div_DP_OP_279J39_124_314_n684), 
        .A3(div_DP_OP_279J39_124_314_n2615), .A4(
        div_DP_OP_279J39_124_314_n2594), .Y(div_DP_OP_279J39_124_314_n2616) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1991 ( .A(div_DP_OP_279J39_124_314_n683), .B(div_DP_OP_279J39_124_314_n670), .CI(div_DP_OP_279J39_124_314_n2616), .S(
        div_n_T_65[65]) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U1990 ( .A1(
        div_DP_OP_279J39_124_314_n683), .A2(div_DP_OP_279J39_124_314_n670), 
        .A3(div_DP_OP_279J39_124_314_n699), .A4(div_DP_OP_279J39_124_314_n684), 
        .Y(div_DP_OP_279J39_124_314_n2612) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1989 ( .A1(
        div_DP_OP_279J39_124_314_n2612), .A2(div_DP_OP_279J39_124_314_n2594), 
        .A3(div_DP_OP_279J39_124_314_n2608), .Y(div_DP_OP_279J39_124_314_n2614) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1988 ( .A(div_DP_OP_279J39_124_314_n669), .B(div_DP_OP_279J39_124_314_n658), .CI(div_DP_OP_279J39_124_314_n2614), .S(
        div_n_T_65[66]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1987 ( .A1(div_DP_OP_279J39_124_314_n669), .A2(div_DP_OP_279J39_124_314_n658), .Y(div_DP_OP_279J39_124_314_n2611) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1986 ( .A1(
        div_DP_OP_279J39_124_314_n669), .A2(div_DP_OP_279J39_124_314_n658), 
        .A3(div_DP_OP_279J39_124_314_n2614), .A4(
        div_DP_OP_279J39_124_314_n2611), .Y(div_DP_OP_279J39_124_314_n2613) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1985 ( .A(div_DP_OP_279J39_124_314_n657), .B(div_DP_OP_279J39_124_314_n648), .CI(div_DP_OP_279J39_124_314_n2613), .S(
        div_n_T_65[67]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1984 ( .A1(div_DP_OP_279J39_124_314_n657), .A2(div_DP_OP_279J39_124_314_n648), .Y(div_DP_OP_279J39_124_314_n2610) );
  AND3X1_LVT div_DP_OP_279J39_124_314_U1983 ( .A1(
        div_DP_OP_279J39_124_314_n2612), .A2(div_DP_OP_279J39_124_314_n2611), 
        .A3(div_DP_OP_279J39_124_314_n2610), .Y(div_DP_OP_279J39_124_314_n2604) );
  OA21X1_LVT div_DP_OP_279J39_124_314_U1982 ( .A1(
        div_DP_OP_279J39_124_314_n648), .A2(div_DP_OP_279J39_124_314_n657), 
        .A3(div_DP_OP_279J39_124_314_n2611), .Y(div_DP_OP_279J39_124_314_n2607) );
  AND3X1_LVT div_DP_OP_279J39_124_314_U1981 ( .A1(
        div_DP_OP_279J39_124_314_n669), .A2(div_DP_OP_279J39_124_314_n658), 
        .A3(div_DP_OP_279J39_124_314_n2610), .Y(div_DP_OP_279J39_124_314_n2609) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U1980 ( .A1(
        div_DP_OP_279J39_124_314_n657), .A2(div_DP_OP_279J39_124_314_n648), 
        .A3(div_DP_OP_279J39_124_314_n2607), .A4(
        div_DP_OP_279J39_124_314_n2608), .A5(div_DP_OP_279J39_124_314_n2609), 
        .Y(div_DP_OP_279J39_124_314_n2601) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1979 ( .A1(
        div_DP_OP_279J39_124_314_n2594), .A2(div_DP_OP_279J39_124_314_n2604), 
        .A3(div_DP_OP_279J39_124_314_n2601), .Y(div_DP_OP_279J39_124_314_n2606) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1978 ( .A(div_DP_OP_279J39_124_314_n647), .B(div_DP_OP_279J39_124_314_n640), .CI(div_DP_OP_279J39_124_314_n2606), .S(
        div_n_T_65[68]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1977 ( .A1(div_DP_OP_279J39_124_314_n647), .A2(div_DP_OP_279J39_124_314_n640), .Y(div_DP_OP_279J39_124_314_n2602) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1976 ( .A1(
        div_DP_OP_279J39_124_314_n647), .A2(div_DP_OP_279J39_124_314_n640), 
        .A3(div_DP_OP_279J39_124_314_n2606), .A4(
        div_DP_OP_279J39_124_314_n2602), .Y(div_DP_OP_279J39_124_314_n2605) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1975 ( .A(div_DP_OP_279J39_124_314_n639), .B(div_DP_OP_279J39_124_314_n634), .CI(div_DP_OP_279J39_124_314_n2605), .S(
        div_n_T_65[69]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1974 ( .A1(div_DP_OP_279J39_124_314_n639), .A2(div_DP_OP_279J39_124_314_n634), .Y(div_DP_OP_279J39_124_314_n2603) );
  AND3X1_LVT div_DP_OP_279J39_124_314_U1973 ( .A1(
        div_DP_OP_279J39_124_314_n2604), .A2(div_DP_OP_279J39_124_314_n2602), 
        .A3(div_DP_OP_279J39_124_314_n2603), .Y(div_DP_OP_279J39_124_314_n2599) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1972 ( .A1(
        div_DP_OP_279J39_124_314_n2599), .A2(div_DP_OP_279J39_124_314_n2594), 
        .A3(div_DP_OP_279J39_124_314_n2598), .Y(div_DP_OP_279J39_124_314_n2600) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1971 ( .A(
        div_DP_OP_279J39_124_314_n2600), .B(div_DP_OP_279J39_124_314_n630), 
        .CI(div_DP_OP_279J39_124_314_n633), .S(div_n_T_65[70]) );
  OA21X1_LVT div_DP_OP_279J39_124_314_U1970 ( .A1(
        div_DP_OP_279J39_124_314_n630), .A2(div_DP_OP_279J39_124_314_n633), 
        .A3(div_DP_OP_279J39_124_314_n2599), .Y(div_DP_OP_279J39_124_314_n2593) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1969 ( .A1(
        div_DP_OP_279J39_124_314_n630), .A2(div_DP_OP_279J39_124_314_n633), 
        .A3(div_DP_OP_279J39_124_314_n630), .A4(div_DP_OP_279J39_124_314_n2598), .A5(div_DP_OP_279J39_124_314_n633), .A6(div_DP_OP_279J39_124_314_n2598), .Y(
        div_DP_OP_279J39_124_314_n2596) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1968 ( .A1(
        div_DP_OP_279J39_124_314_n2594), .A2(div_DP_OP_279J39_124_314_n2593), 
        .A3(div_DP_OP_279J39_124_314_n2596), .Y(div_DP_OP_279J39_124_314_n2597) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1967 ( .A(
        div_DP_OP_279J39_124_314_n2597), .B(div_DP_OP_279J39_124_314_n628), 
        .CI(div_DP_OP_279J39_124_314_n629), .S(div_n_T_65[71]) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1966 ( .A1(div_DP_OP_279J39_124_314_n628), .A2(div_DP_OP_279J39_124_314_n629), .Y(div_DP_OP_279J39_124_314_n2595) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1965 ( .A1(
        div_DP_OP_279J39_124_314_n2596), .A2(div_DP_OP_279J39_124_314_n2595), 
        .A3(div_DP_OP_279J39_124_314_n628), .A4(div_DP_OP_279J39_124_314_n629), 
        .Y(div_DP_OP_279J39_124_314_n2592) );
  OA222X1_LVT div_DP_OP_279J39_124_314_U1964 ( .A1(
        div_DP_OP_279J39_124_314_n2592), .A2(div_DP_OP_279J39_124_314_n2593), 
        .A3(div_DP_OP_279J39_124_314_n2592), .A4(
        div_DP_OP_279J39_124_314_n2594), .A5(div_DP_OP_279J39_124_314_n2592), 
        .A6(div_DP_OP_279J39_124_314_n2595), .Y(div_DP_OP_279J39_124_314_n2590) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U1963 ( .A1(div_n301), .A2(
        div_divisor_64_), .Y(div_DP_OP_279J39_124_314_n2591) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1962 ( .A(
        div_DP_OP_279J39_124_314_n2590), .B(div_DP_OP_279J39_124_314_n627), 
        .CI(div_DP_OP_279J39_124_314_n2591), .S(div_n_T_65[72]) );
  INVX1_LVT div_DP_OP_279J39_124_314_U1961 ( .A(div_n_T_51_72_), .Y(
        div_DP_OP_279J39_124_314_n2588) );
  INVX1_LVT div_DP_OP_279J39_124_314_U1960 ( .A(div_n_T_51_128_), .Y(
        div_DP_OP_279J39_124_314_n2587) );
  INVX1_LVT div_DP_OP_279J39_124_314_U1959 ( .A(div_DP_OP_279J39_124_314_n2589), .Y(div_DP_OP_279J39_124_314_n2586) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1958 ( .A(div_n_T_51_7_), .Y(
        div_DP_OP_279J39_124_314_n2585) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1957 ( .A(div_n_T_51_5_), .Y(
        div_DP_OP_279J39_124_314_n2584) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1956 ( .A(div_divisor_4_), .Y(
        div_DP_OP_279J39_124_314_n2557) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1955 ( .A(div_divisor_7_), .Y(
        div_DP_OP_279J39_124_314_n2559) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1954 ( .A(div_divisor_36_), .Y(
        div_DP_OP_279J39_124_314_n2569) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1953 ( .A(div_divisor_30_), .Y(
        div_DP_OP_279J39_124_314_n2567) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1952 ( .A(div_divisor_31_), .Y(
        div_DP_OP_279J39_124_314_n2568) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1951 ( .A(div_divisor_28_), .Y(
        div_DP_OP_279J39_124_314_n2566) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1950 ( .A(div_divisor_37_), .Y(
        div_DP_OP_279J39_124_314_n2570) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1949 ( .A(div_divisor_20_), .Y(
        div_DP_OP_279J39_124_314_n2564) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1948 ( .A(div_divisor_13_), .Y(
        div_DP_OP_279J39_124_314_n2562) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1947 ( .A(div_divisor_12_), .Y(
        div_DP_OP_279J39_124_314_n2561) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1946 ( .A(div_divisor_9_), .Y(
        div_DP_OP_279J39_124_314_n2560) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1945 ( .A(div_divisor_45_), .Y(
        div_DP_OP_279J39_124_314_n2573) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1944 ( .A(div_divisor_44_), .Y(
        div_DP_OP_279J39_124_314_n2572) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1943 ( .A(div_divisor_53_), .Y(
        div_DP_OP_279J39_124_314_n2576) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1942 ( .A(div_divisor_52_), .Y(
        div_DP_OP_279J39_124_314_n2575) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1941 ( .A(div_divisor_55_), .Y(
        div_DP_OP_279J39_124_314_n2578) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1940 ( .A(div_divisor_56_), .Y(
        div_DP_OP_279J39_124_314_n2579) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1939 ( .A(div_divisor_57_), .Y(
        div_DP_OP_279J39_124_314_n2580) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1938 ( .A(div_divisor_60_), .Y(
        div_DP_OP_279J39_124_314_n2581) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1937 ( .A(div_divisor_63_), .Y(
        div_DP_OP_279J39_124_314_n2583) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1936 ( .A(div_divisor_22_), .Y(
        div_DP_OP_279J39_124_314_n2565) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1935 ( .A(div_divisor_54_), .Y(
        div_DP_OP_279J39_124_314_n2577) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1934 ( .A(div_divisor_38_), .Y(
        div_DP_OP_279J39_124_314_n2571) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1933 ( .A(div_divisor_46_), .Y(
        div_DP_OP_279J39_124_314_n2574) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1932 ( .A(div_divisor_61_), .Y(
        div_DP_OP_279J39_124_314_n2582) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1931 ( .A(div_divisor_6_), .Y(
        div_DP_OP_279J39_124_314_n2558) );
  NBUFFX2_LVT div_DP_OP_279J39_124_314_U1930 ( .A(div_divisor_14_), .Y(
        div_DP_OP_279J39_124_314_n2563) );
  AND2X1_LVT div_DP_OP_279J39_124_314_U1929 ( .A1(
        div_DP_OP_279J39_124_314_n2603), .A2(div_DP_OP_279J39_124_314_n2556), 
        .Y(div_DP_OP_279J39_124_314_n2598) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1928 ( .A1(
        div_DP_OP_279J39_124_314_n639), .A2(div_DP_OP_279J39_124_314_n634), 
        .A3(div_DP_OP_279J39_124_314_n647), .A4(div_DP_OP_279J39_124_314_n640), 
        .A5(div_DP_OP_279J39_124_314_n2602), .A6(
        div_DP_OP_279J39_124_314_n2601), .Y(div_DP_OP_279J39_124_314_n2556) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1927 ( .A1(
        div_DP_OP_279J39_124_314_n1387), .A2(div_DP_OP_279J39_124_314_n1372), 
        .A3(div_DP_OP_279J39_124_314_n1387), .A4(
        div_DP_OP_279J39_124_314_n2745), .A5(div_DP_OP_279J39_124_314_n1372), 
        .A6(div_DP_OP_279J39_124_314_n2745), .Y(div_DP_OP_279J39_124_314_n2736) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1926 ( .A1(
        div_DP_OP_279J39_124_314_n1323), .A2(div_DP_OP_279J39_124_314_n1308), 
        .A3(div_DP_OP_279J39_124_314_n1323), .A4(
        div_DP_OP_279J39_124_314_n2733), .A5(div_DP_OP_279J39_124_314_n1308), 
        .A6(div_DP_OP_279J39_124_314_n2733), .Y(div_DP_OP_279J39_124_314_n2729) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1925 ( .A1(
        div_DP_OP_279J39_124_314_n1195), .A2(div_DP_OP_279J39_124_314_n1180), 
        .A3(div_DP_OP_279J39_124_314_n1195), .A4(
        div_DP_OP_279J39_124_314_n2710), .A5(div_DP_OP_279J39_124_314_n1180), 
        .A6(div_DP_OP_279J39_124_314_n2710), .Y(div_DP_OP_279J39_124_314_n2706) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1924 ( .A1(
        div_DP_OP_279J39_124_314_n1131), .A2(div_DP_OP_279J39_124_314_n1116), 
        .A3(div_DP_OP_279J39_124_314_n1131), .A4(
        div_DP_OP_279J39_124_314_n2701), .A5(div_DP_OP_279J39_124_314_n1116), 
        .A6(div_DP_OP_279J39_124_314_n2701), .Y(div_DP_OP_279J39_124_314_n2692) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1923 ( .A1(
        div_DP_OP_279J39_124_314_n1067), .A2(div_DP_OP_279J39_124_314_n1052), 
        .A3(div_DP_OP_279J39_124_314_n1067), .A4(
        div_DP_OP_279J39_124_314_n2689), .A5(div_DP_OP_279J39_124_314_n1052), 
        .A6(div_DP_OP_279J39_124_314_n2689), .Y(div_DP_OP_279J39_124_314_n2685) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1922 ( .A1(
        div_DP_OP_279J39_124_314_n1003), .A2(div_DP_OP_279J39_124_314_n988), 
        .A3(div_DP_OP_279J39_124_314_n1003), .A4(
        div_DP_OP_279J39_124_314_n2679), .A5(div_DP_OP_279J39_124_314_n988), 
        .A6(div_DP_OP_279J39_124_314_n2679), .Y(div_DP_OP_279J39_124_314_n2672) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1921 ( .A1(
        div_DP_OP_279J39_124_314_n939), .A2(div_DP_OP_279J39_124_314_n924), 
        .A3(div_DP_OP_279J39_124_314_n939), .A4(div_DP_OP_279J39_124_314_n2662), .A5(div_DP_OP_279J39_124_314_n924), .A6(div_DP_OP_279J39_124_314_n2662), .Y(
        div_DP_OP_279J39_124_314_n2658) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1920 ( .A1(
        div_DP_OP_279J39_124_314_n875), .A2(div_DP_OP_279J39_124_314_n860), 
        .A3(div_DP_OP_279J39_124_314_n875), .A4(div_DP_OP_279J39_124_314_n2653), .A5(div_DP_OP_279J39_124_314_n860), .A6(div_DP_OP_279J39_124_314_n2653), .Y(
        div_DP_OP_279J39_124_314_n2644) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1919 ( .A1(
        div_DP_OP_279J39_124_314_n811), .A2(div_DP_OP_279J39_124_314_n796), 
        .A3(div_DP_OP_279J39_124_314_n811), .A4(div_DP_OP_279J39_124_314_n2640), .A5(div_DP_OP_279J39_124_314_n796), .A6(div_DP_OP_279J39_124_314_n2640), .Y(
        div_DP_OP_279J39_124_314_n2636) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1918 ( .A1(
        div_DP_OP_279J39_124_314_n747), .A2(div_DP_OP_279J39_124_314_n732), 
        .A3(div_DP_OP_279J39_124_314_n747), .A4(div_DP_OP_279J39_124_314_n2630), .A5(div_DP_OP_279J39_124_314_n732), .A6(div_DP_OP_279J39_124_314_n2630), .Y(
        div_DP_OP_279J39_124_314_n2622) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1917 ( .A1(
        div_DP_OP_279J39_124_314_n1579), .A2(div_DP_OP_279J39_124_314_n1564), 
        .A3(div_DP_OP_279J39_124_314_n1579), .A4(
        div_DP_OP_279J39_124_314_n2774), .A5(div_DP_OP_279J39_124_314_n1564), 
        .A6(div_DP_OP_279J39_124_314_n2774), .Y(div_DP_OP_279J39_124_314_n2770) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1916 ( .A1(
        div_DP_OP_279J39_124_314_n1515), .A2(div_DP_OP_279J39_124_314_n1500), 
        .A3(div_DP_OP_279J39_124_314_n1515), .A4(
        div_DP_OP_279J39_124_314_n2765), .A5(div_DP_OP_279J39_124_314_n1500), 
        .A6(div_DP_OP_279J39_124_314_n2765), .Y(div_DP_OP_279J39_124_314_n2758) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1915 ( .A1(
        div_DP_OP_279J39_124_314_n1451), .A2(div_DP_OP_279J39_124_314_n1436), 
        .A3(div_DP_OP_279J39_124_314_n1451), .A4(
        div_DP_OP_279J39_124_314_n2754), .A5(div_DP_OP_279J39_124_314_n1436), 
        .A6(div_DP_OP_279J39_124_314_n2754), .Y(div_DP_OP_279J39_124_314_n2750) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1914 ( .A1(
        div_DP_OP_279J39_124_314_n1259), .A2(div_DP_OP_279J39_124_314_n1244), 
        .A3(div_DP_OP_279J39_124_314_n1259), .A4(
        div_DP_OP_279J39_124_314_n2723), .A5(div_DP_OP_279J39_124_314_n1244), 
        .A6(div_DP_OP_279J39_124_314_n2723), .Y(div_DP_OP_279J39_124_314_n2713) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U1913 ( .A1(
        div_DP_OP_279J39_124_314_n2555), .A2(div_DP_OP_279J39_124_314_n1099), 
        .A3(div_DP_OP_279J39_124_314_n2695), .A4(
        div_DP_OP_279J39_124_314_n1084), .A5(div_DP_OP_279J39_124_314_n2554), 
        .Y(div_DP_OP_279J39_124_314_n2667) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1912 ( .A1(
        div_DP_OP_279J39_124_314_n1084), .A2(div_DP_OP_279J39_124_314_n2695), 
        .Y(div_DP_OP_279J39_124_314_n2555) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1911 ( .A1(
        div_DP_OP_279J39_124_314_n2691), .A2(div_DP_OP_279J39_124_314_n2692), 
        .A3(div_DP_OP_279J39_124_314_n2694), .A4(
        div_DP_OP_279J39_124_314_n2693), .Y(div_DP_OP_279J39_124_314_n2554) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U1910 ( .A1(
        div_DP_OP_279J39_124_314_n2552), .A2(div_DP_OP_279J39_124_314_n843), 
        .A3(div_DP_OP_279J39_124_314_n2647), .A4(div_DP_OP_279J39_124_314_n828), .A5(div_DP_OP_279J39_124_314_n2553), .Y(div_DP_OP_279J39_124_314_n2620) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1909 ( .A1(
        div_DP_OP_279J39_124_314_n2643), .A2(div_DP_OP_279J39_124_314_n2644), 
        .A3(div_DP_OP_279J39_124_314_n2646), .A4(
        div_DP_OP_279J39_124_314_n2645), .Y(div_DP_OP_279J39_124_314_n2553) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1908 ( .A1(div_DP_OP_279J39_124_314_n828), .A2(div_DP_OP_279J39_124_314_n2647), .Y(div_DP_OP_279J39_124_314_n2552) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1907 ( .A1(
        div_DP_OP_279J39_124_314_n683), .A2(div_DP_OP_279J39_124_314_n670), 
        .A3(div_DP_OP_279J39_124_314_n683), .A4(div_DP_OP_279J39_124_314_n2615), .A5(div_DP_OP_279J39_124_314_n670), .A6(div_DP_OP_279J39_124_314_n2615), .Y(
        div_DP_OP_279J39_124_314_n2608) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1906 ( .A1(
        div_DP_OP_279J39_124_314_n2549), .A2(div_DP_OP_279J39_124_314_n2550), 
        .A3(div_DP_OP_279J39_124_314_n2551), .A4(
        div_DP_OP_279J39_124_314_n2760), .A5(div_DP_OP_279J39_124_314_n1468), 
        .A6(div_DP_OP_279J39_124_314_n1483), .Y(div_DP_OP_279J39_124_314_n2716) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1905 ( .A1(
        div_DP_OP_279J39_124_314_n1483), .A2(div_DP_OP_279J39_124_314_n1468), 
        .Y(div_DP_OP_279J39_124_314_n2551) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U1904 ( .A1(
        div_DP_OP_279J39_124_314_n1499), .A2(div_DP_OP_279J39_124_314_n1484), 
        .A3(div_DP_OP_279J39_124_314_n1483), .A4(
        div_DP_OP_279J39_124_314_n1468), .Y(div_DP_OP_279J39_124_314_n2550) );
  AND3X1_LVT div_DP_OP_279J39_124_314_U1902 ( .A1(
        div_DP_OP_279J39_124_314_n2757), .A2(div_DP_OP_279J39_124_314_n2761), 
        .A3(div_DP_OP_279J39_124_314_n2756), .Y(div_DP_OP_279J39_124_314_n2547) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1901 ( .A1(
        div_DP_OP_279J39_124_314_n1645), .A2(div_DP_OP_279J39_124_314_n1640), 
        .A3(div_DP_OP_279J39_124_314_n1645), .A4(
        div_DP_OP_279J39_124_314_n2546), .A5(div_DP_OP_279J39_124_314_n1640), 
        .A6(div_DP_OP_279J39_124_314_n2546), .Y(div_DP_OP_279J39_124_314_n2778) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1900 ( .A1(
        div_DP_OP_279J39_124_314_n2784), .A2(div_DP_OP_279J39_124_314_n551), 
        .A3(div_DP_OP_279J39_124_314_n2785), .Y(div_DP_OP_279J39_124_314_n2546) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U1899 ( .A1(
        div_DP_OP_279J39_124_314_n2544), .A2(div_DP_OP_279J39_124_314_n1355), 
        .A3(div_DP_OP_279J39_124_314_n2739), .A4(
        div_DP_OP_279J39_124_314_n1340), .A5(div_DP_OP_279J39_124_314_n2545), 
        .Y(div_DP_OP_279J39_124_314_n2712) );
  AO22X1_LVT div_DP_OP_279J39_124_314_U1898 ( .A1(
        div_DP_OP_279J39_124_314_n2735), .A2(div_DP_OP_279J39_124_314_n2736), 
        .A3(div_DP_OP_279J39_124_314_n2738), .A4(
        div_DP_OP_279J39_124_314_n2737), .Y(div_DP_OP_279J39_124_314_n2545) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1897 ( .A1(
        div_DP_OP_279J39_124_314_n1340), .A2(div_DP_OP_279J39_124_314_n2739), 
        .Y(div_DP_OP_279J39_124_314_n2544) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1896 ( .A1(
        div_DP_OP_279J39_124_314_n2541), .A2(div_DP_OP_279J39_124_314_n2542), 
        .A3(div_DP_OP_279J39_124_314_n2543), .A4(
        div_DP_OP_279J39_124_314_n2777), .A5(div_DP_OP_279J39_124_314_n1596), 
        .A6(div_DP_OP_279J39_124_314_n1609), .Y(div_DP_OP_279J39_124_314_n2757) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1895 ( .A1(
        div_DP_OP_279J39_124_314_n1609), .A2(div_DP_OP_279J39_124_314_n1596), 
        .Y(div_DP_OP_279J39_124_314_n2543) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U1894 ( .A1(
        div_DP_OP_279J39_124_314_n1621), .A2(div_DP_OP_279J39_124_314_n1610), 
        .A3(div_DP_OP_279J39_124_314_n1609), .A4(
        div_DP_OP_279J39_124_314_n1596), .Y(div_DP_OP_279J39_124_314_n2542) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1893 ( .A1(
        div_DP_OP_279J39_124_314_n2778), .A2(div_DP_OP_279J39_124_314_n2779), 
        .A3(div_DP_OP_279J39_124_314_n2776), .Y(div_DP_OP_279J39_124_314_n2541) );
  AO222X1_LVT div_DP_OP_279J39_124_314_U1891 ( .A1(
        div_DP_OP_279J39_124_314_n1631), .A2(div_DP_OP_279J39_124_314_n1622), 
        .A3(div_DP_OP_279J39_124_314_n1631), .A4(
        div_DP_OP_279J39_124_314_n2782), .A5(div_DP_OP_279J39_124_314_n1622), 
        .A6(div_DP_OP_279J39_124_314_n2782), .Y(div_DP_OP_279J39_124_314_n2776) );
  OA221X1_LVT div_DP_OP_279J39_124_314_U1890 ( .A1(div_n_T_51_64_), .A2(
        div_divisor_0_), .A3(div_n_T_51_64_), .A4(div_n302), .A5(
        div_DP_OP_279J39_124_314_n2589), .Y(div_n_T_65[0]) );
  AO21X1_LVT div_DP_OP_279J39_124_314_U1889 ( .A1(
        div_DP_OP_279J39_124_314_n1212), .A2(div_DP_OP_279J39_124_314_n1227), 
        .A3(div_DP_OP_279J39_124_314_n2539), .Y(div_DP_OP_279J39_124_314_n2618) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U1888 ( .A1(
        div_DP_OP_279J39_124_314_n2538), .A2(div_DP_OP_279J39_124_314_n2715), 
        .A3(div_DP_OP_279J39_124_314_n1227), .A4(
        div_DP_OP_279J39_124_314_n1212), .Y(div_DP_OP_279J39_124_314_n2539) );
  OA22X1_LVT div_DP_OP_279J39_124_314_U1887 ( .A1(
        div_DP_OP_279J39_124_314_n1243), .A2(div_DP_OP_279J39_124_314_n1228), 
        .A3(div_DP_OP_279J39_124_314_n2537), .A4(
        div_DP_OP_279J39_124_314_n2713), .Y(div_DP_OP_279J39_124_314_n2538) );
  OA221X1_LVT div_DP_OP_279J39_124_314_U1886 ( .A1(
        div_DP_OP_279J39_124_314_n2712), .A2(div_DP_OP_279J39_124_314_n2716), 
        .A3(div_DP_OP_279J39_124_314_n2712), .A4(
        div_DP_OP_279J39_124_314_n2717), .A5(div_DP_OP_279J39_124_314_n2718), 
        .Y(div_DP_OP_279J39_124_314_n2536) );
  NAND4X0_LVT div_DP_OP_279J39_124_314_U1885 ( .A1(
        div_DP_OP_279J39_124_314_n2529), .A2(div_DP_OP_279J39_124_314_n2533), 
        .A3(div_DP_OP_279J39_124_314_n2534), .A4(
        div_DP_OP_279J39_124_314_n2535), .Y(div_DP_OP_279J39_124_314_n2594) );
  NAND3X0_LVT div_DP_OP_279J39_124_314_U1884 ( .A1(
        div_DP_OP_279J39_124_314_n716), .A2(div_DP_OP_279J39_124_314_n731), 
        .A3(div_DP_OP_279J39_124_314_n2527), .Y(div_DP_OP_279J39_124_314_n2535) );
  NAND3X0_LVT div_DP_OP_279J39_124_314_U1883 ( .A1(
        div_DP_OP_279J39_124_314_n2621), .A2(div_DP_OP_279J39_124_314_n2622), 
        .A3(div_DP_OP_279J39_124_314_n2527), .Y(div_DP_OP_279J39_124_314_n2534) );
  NAND3X0_LVT div_DP_OP_279J39_124_314_U1882 ( .A1(
        div_DP_OP_279J39_124_314_n2626), .A2(div_DP_OP_279J39_124_314_n2528), 
        .A3(div_DP_OP_279J39_124_314_n2532), .Y(div_DP_OP_279J39_124_314_n2533) );
  AND3X1_LVT div_DP_OP_279J39_124_314_U1880 ( .A1(
        div_DP_OP_279J39_124_314_n2618), .A2(div_DP_OP_279J39_124_314_n2625), 
        .A3(div_DP_OP_279J39_124_314_n2617), .Y(div_DP_OP_279J39_124_314_n2530) );
  AOI22X1_LVT div_DP_OP_279J39_124_314_U1879 ( .A1(
        div_DP_OP_279J39_124_314_n715), .A2(div_DP_OP_279J39_124_314_n700), 
        .A3(div_DP_OP_279J39_124_314_n2528), .A4(
        div_DP_OP_279J39_124_314_n2624), .Y(div_DP_OP_279J39_124_314_n2529) );
  AND3X1_LVT div_DP_OP_279J39_124_314_U1878 ( .A1(
        div_DP_OP_279J39_124_314_n2621), .A2(div_DP_OP_279J39_124_314_n2623), 
        .A3(div_DP_OP_279J39_124_314_n2527), .Y(div_DP_OP_279J39_124_314_n2528) );
  OR2X1_LVT div_DP_OP_279J39_124_314_U1877 ( .A1(div_DP_OP_279J39_124_314_n715), .A2(div_DP_OP_279J39_124_314_n700), .Y(div_DP_OP_279J39_124_314_n2527) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U1876 ( .A1(1'b1), .A2(
        div_DP_OP_279J39_124_314_n2530), .A3(div_DP_OP_279J39_124_314_n2625), 
        .A4(div_DP_OP_279J39_124_314_n2619), .A5(
        div_DP_OP_279J39_124_314_n2620), .Y(div_DP_OP_279J39_124_314_n2532) );
  OA221X1_LVT div_DP_OP_279J39_124_314_U1875 ( .A1(
        div_DP_OP_279J39_124_314_n2714), .A2(1'b1), .A3(
        div_DP_OP_279J39_124_314_n2714), .A4(div_DP_OP_279J39_124_314_n2536), 
        .A5(div_DP_OP_279J39_124_314_n2719), .Y(div_DP_OP_279J39_124_314_n2537) );
  AO221X1_LVT div_DP_OP_279J39_124_314_U1874 ( .A1(1'b1), .A2(
        div_DP_OP_279J39_124_314_n2547), .A3(div_DP_OP_279J39_124_314_n2761), 
        .A4(div_DP_OP_279J39_124_314_n2759), .A5(
        div_DP_OP_279J39_124_314_n2758), .Y(div_DP_OP_279J39_124_314_n2549) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1211 ( .A0(div_n_T_51_65_), .B0(
        div_DP_OP_279J39_124_314_n2235), .C1(div_DP_OP_279J39_124_314_n1649), 
        .SO(div_DP_OP_279J39_124_314_n1650) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1210 ( .A0(div_n_T_51_66_), .B0(
        div_DP_OP_279J39_124_314_n2234), .C1(div_DP_OP_279J39_124_314_n1647), 
        .SO(div_DP_OP_279J39_124_314_n1648) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1209 ( .A(
        div_DP_OP_279J39_124_314_n2170), .B(div_DP_OP_279J39_124_314_n2106), 
        .CI(div_DP_OP_279J39_124_314_n1649), .CO(
        div_DP_OP_279J39_124_314_n1645), .S(div_DP_OP_279J39_124_314_n1646) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1208 ( .A0(div_n_T_51_67_), .B0(
        div_DP_OP_279J39_124_314_n2105), .C1(div_DP_OP_279J39_124_314_n1643), 
        .SO(div_DP_OP_279J39_124_314_n1644) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1207 ( .A(
        div_DP_OP_279J39_124_314_n2233), .B(div_DP_OP_279J39_124_314_n2041), 
        .CI(div_DP_OP_279J39_124_314_n2169), .CO(
        div_DP_OP_279J39_124_314_n1641), .S(div_DP_OP_279J39_124_314_n1642) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1206 ( .A(
        div_DP_OP_279J39_124_314_n1647), .B(div_DP_OP_279J39_124_314_n1644), 
        .CI(div_DP_OP_279J39_124_314_n1642), .CO(
        div_DP_OP_279J39_124_314_n1639), .S(div_DP_OP_279J39_124_314_n1640) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1205 ( .A0(div_n_T_51_68_), .B0(
        div_DP_OP_279J39_124_314_n2040), .C1(div_DP_OP_279J39_124_314_n1637), 
        .SO(div_DP_OP_279J39_124_314_n1638) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1204 ( .A(
        div_DP_OP_279J39_124_314_n2232), .B(div_DP_OP_279J39_124_314_n1976), 
        .CI(div_DP_OP_279J39_124_314_n2104), .CO(
        div_DP_OP_279J39_124_314_n1635), .S(div_DP_OP_279J39_124_314_n1636) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1203 ( .A(
        div_DP_OP_279J39_124_314_n2168), .B(div_DP_OP_279J39_124_314_n1643), 
        .CI(div_DP_OP_279J39_124_314_n1638), .CO(
        div_DP_OP_279J39_124_314_n1633), .S(div_DP_OP_279J39_124_314_n1634) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1202 ( .A(
        div_DP_OP_279J39_124_314_n1641), .B(div_DP_OP_279J39_124_314_n1636), 
        .CI(div_DP_OP_279J39_124_314_n1634), .CO(
        div_DP_OP_279J39_124_314_n1631), .S(div_DP_OP_279J39_124_314_n1632) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1201 ( .A0(div_n_T_51_69_), .B0(
        div_DP_OP_279J39_124_314_n1975), .C1(div_DP_OP_279J39_124_314_n1629), 
        .SO(div_DP_OP_279J39_124_314_n1630) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1200 ( .A(
        div_DP_OP_279J39_124_314_n2231), .B(div_DP_OP_279J39_124_314_n1911), 
        .CI(div_DP_OP_279J39_124_314_n2167), .CO(
        div_DP_OP_279J39_124_314_n1627), .S(div_DP_OP_279J39_124_314_n1628) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1199 ( .A(
        div_DP_OP_279J39_124_314_n2103), .B(div_DP_OP_279J39_124_314_n2039), 
        .CI(div_DP_OP_279J39_124_314_n1637), .CO(
        div_DP_OP_279J39_124_314_n1625), .S(div_DP_OP_279J39_124_314_n1626) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1198 ( .A(
        div_DP_OP_279J39_124_314_n1630), .B(div_DP_OP_279J39_124_314_n1635), 
        .CI(div_DP_OP_279J39_124_314_n1628), .CO(
        div_DP_OP_279J39_124_314_n1623), .S(div_DP_OP_279J39_124_314_n1624) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1197 ( .A(
        div_DP_OP_279J39_124_314_n1633), .B(div_DP_OP_279J39_124_314_n1626), 
        .CI(div_DP_OP_279J39_124_314_n1624), .CO(
        div_DP_OP_279J39_124_314_n1621), .S(div_DP_OP_279J39_124_314_n1622) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1196 ( .A0(div_n_T_51_70_), .B0(
        div_DP_OP_279J39_124_314_n1910), .C1(div_DP_OP_279J39_124_314_n1619), 
        .SO(div_DP_OP_279J39_124_314_n1620) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1195 ( .A(
        div_DP_OP_279J39_124_314_n2230), .B(div_DP_OP_279J39_124_314_n1846), 
        .CI(div_DP_OP_279J39_124_314_n2166), .CO(
        div_DP_OP_279J39_124_314_n1617), .S(div_DP_OP_279J39_124_314_n1618) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1194 ( .A(
        div_DP_OP_279J39_124_314_n2102), .B(div_DP_OP_279J39_124_314_n1974), 
        .CI(div_DP_OP_279J39_124_314_n2038), .CO(
        div_DP_OP_279J39_124_314_n1615), .S(div_DP_OP_279J39_124_314_n1616) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1193 ( .A(
        div_DP_OP_279J39_124_314_n1629), .B(div_DP_OP_279J39_124_314_n1620), 
        .CI(div_DP_OP_279J39_124_314_n1627), .CO(
        div_DP_OP_279J39_124_314_n1613), .S(div_DP_OP_279J39_124_314_n1614) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1192 ( .A(
        div_DP_OP_279J39_124_314_n1616), .B(div_DP_OP_279J39_124_314_n1618), 
        .CI(div_DP_OP_279J39_124_314_n1625), .CO(
        div_DP_OP_279J39_124_314_n1611), .S(div_DP_OP_279J39_124_314_n1612) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1191 ( .A(
        div_DP_OP_279J39_124_314_n1623), .B(div_DP_OP_279J39_124_314_n1614), 
        .CI(div_DP_OP_279J39_124_314_n1612), .CO(
        div_DP_OP_279J39_124_314_n1609), .S(div_DP_OP_279J39_124_314_n1610) );
  HADDX1_LVT div_DP_OP_279J39_124_314_U1190 ( .A0(div_n_T_51_71_), .B0(
        div_DP_OP_279J39_124_314_n1845), .C1(div_DP_OP_279J39_124_314_n1607), 
        .SO(div_DP_OP_279J39_124_314_n1608) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1189 ( .A(
        div_DP_OP_279J39_124_314_n2229), .B(div_DP_OP_279J39_124_314_n1781), 
        .CI(div_DP_OP_279J39_124_314_n2165), .CO(
        div_DP_OP_279J39_124_314_n1605), .S(div_DP_OP_279J39_124_314_n1606) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1188 ( .A(
        div_DP_OP_279J39_124_314_n1973), .B(div_DP_OP_279J39_124_314_n2101), 
        .CI(div_DP_OP_279J39_124_314_n1909), .CO(
        div_DP_OP_279J39_124_314_n1603), .S(div_DP_OP_279J39_124_314_n1604) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1187 ( .A(
        div_DP_OP_279J39_124_314_n2037), .B(div_DP_OP_279J39_124_314_n1619), 
        .CI(div_DP_OP_279J39_124_314_n1608), .CO(
        div_DP_OP_279J39_124_314_n1601), .S(div_DP_OP_279J39_124_314_n1602) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1186 ( .A(
        div_DP_OP_279J39_124_314_n1617), .B(div_DP_OP_279J39_124_314_n1615), 
        .CI(div_DP_OP_279J39_124_314_n1604), .CO(
        div_DP_OP_279J39_124_314_n1599), .S(div_DP_OP_279J39_124_314_n1600) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1185 ( .A(
        div_DP_OP_279J39_124_314_n1606), .B(div_DP_OP_279J39_124_314_n1613), 
        .CI(div_DP_OP_279J39_124_314_n1602), .CO(
        div_DP_OP_279J39_124_314_n1597), .S(div_DP_OP_279J39_124_314_n1598) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1184 ( .A(
        div_DP_OP_279J39_124_314_n1611), .B(div_DP_OP_279J39_124_314_n1600), 
        .CI(div_DP_OP_279J39_124_314_n1598), .CO(
        div_DP_OP_279J39_124_314_n1595), .S(div_DP_OP_279J39_124_314_n1596) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1181 ( .A(
        div_DP_OP_279J39_124_314_n2228), .B(div_DP_OP_279J39_124_314_n1780), 
        .CI(div_DP_OP_279J39_124_314_n1844), .CO(
        div_DP_OP_279J39_124_314_n1591), .S(div_DP_OP_279J39_124_314_n1592) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1180 ( .A(
        div_DP_OP_279J39_124_314_n2164), .B(div_DP_OP_279J39_124_314_n1908), 
        .CI(div_DP_OP_279J39_124_314_n1972), .CO(
        div_DP_OP_279J39_124_314_n1589), .S(div_DP_OP_279J39_124_314_n1590) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1179 ( .A(
        div_DP_OP_279J39_124_314_n2100), .B(div_DP_OP_279J39_124_314_n2036), 
        .CI(div_DP_OP_279J39_124_314_n1607), .CO(
        div_DP_OP_279J39_124_314_n1587), .S(div_DP_OP_279J39_124_314_n1588) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1178 ( .A(
        div_DP_OP_279J39_124_314_n1605), .B(div_DP_OP_279J39_124_314_n1603), 
        .CI(div_DP_OP_279J39_124_314_n1594), .CO(
        div_DP_OP_279J39_124_314_n1585), .S(div_DP_OP_279J39_124_314_n1586) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1177 ( .A(
        div_DP_OP_279J39_124_314_n1590), .B(div_DP_OP_279J39_124_314_n1592), 
        .CI(div_DP_OP_279J39_124_314_n1601), .CO(
        div_DP_OP_279J39_124_314_n1583), .S(div_DP_OP_279J39_124_314_n1584) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1176 ( .A(
        div_DP_OP_279J39_124_314_n1588), .B(div_DP_OP_279J39_124_314_n1599), 
        .CI(div_DP_OP_279J39_124_314_n1586), .CO(
        div_DP_OP_279J39_124_314_n1581), .S(div_DP_OP_279J39_124_314_n1582) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1175 ( .A(
        div_DP_OP_279J39_124_314_n1597), .B(div_DP_OP_279J39_124_314_n1584), 
        .CI(div_DP_OP_279J39_124_314_n1582), .CO(
        div_DP_OP_279J39_124_314_n1579), .S(div_DP_OP_279J39_124_314_n1580) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1174 ( .A(div_n_T_51_73_), .B(
        div_DP_OP_279J39_124_314_n1715), .CI(div_DP_OP_279J39_124_314_n2227), 
        .CO(div_DP_OP_279J39_124_314_n1577), .S(div_DP_OP_279J39_124_314_n1578) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1173 ( .A(
        div_DP_OP_279J39_124_314_n2163), .B(div_DP_OP_279J39_124_314_n1779), 
        .CI(div_DP_OP_279J39_124_314_n1843), .CO(
        div_DP_OP_279J39_124_314_n1575), .S(div_DP_OP_279J39_124_314_n1576) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1172 ( .A(
        div_DP_OP_279J39_124_314_n2099), .B(div_DP_OP_279J39_124_314_n1907), 
        .CI(div_DP_OP_279J39_124_314_n1971), .CO(
        div_DP_OP_279J39_124_314_n1573), .S(div_DP_OP_279J39_124_314_n1574) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1171 ( .A(
        div_DP_OP_279J39_124_314_n2035), .B(div_DP_OP_279J39_124_314_n1593), 
        .CI(div_DP_OP_279J39_124_314_n1591), .CO(
        div_DP_OP_279J39_124_314_n1571), .S(div_DP_OP_279J39_124_314_n1572) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1170 ( .A(
        div_DP_OP_279J39_124_314_n1589), .B(div_DP_OP_279J39_124_314_n1578), 
        .CI(div_DP_OP_279J39_124_314_n1574), .CO(
        div_DP_OP_279J39_124_314_n1569), .S(div_DP_OP_279J39_124_314_n1570) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1169 ( .A(
        div_DP_OP_279J39_124_314_n1576), .B(div_DP_OP_279J39_124_314_n1587), 
        .CI(div_DP_OP_279J39_124_314_n1585), .CO(
        div_DP_OP_279J39_124_314_n1567), .S(div_DP_OP_279J39_124_314_n1568) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1168 ( .A(
        div_DP_OP_279J39_124_314_n1572), .B(div_DP_OP_279J39_124_314_n1583), 
        .CI(div_DP_OP_279J39_124_314_n1570), .CO(
        div_DP_OP_279J39_124_314_n1565), .S(div_DP_OP_279J39_124_314_n1566) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1167 ( .A(
        div_DP_OP_279J39_124_314_n1581), .B(div_DP_OP_279J39_124_314_n1568), 
        .CI(div_DP_OP_279J39_124_314_n1566), .CO(
        div_DP_OP_279J39_124_314_n1563), .S(div_DP_OP_279J39_124_314_n1564) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1166 ( .A(div_n_T_51_74_), .B(
        div_DP_OP_279J39_124_314_n1714), .CI(div_DP_OP_279J39_124_314_n2226), 
        .CO(div_DP_OP_279J39_124_314_n1561), .S(div_DP_OP_279J39_124_314_n1562) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1165 ( .A(
        div_DP_OP_279J39_124_314_n2162), .B(div_DP_OP_279J39_124_314_n1778), 
        .CI(div_DP_OP_279J39_124_314_n1842), .CO(
        div_DP_OP_279J39_124_314_n1559), .S(div_DP_OP_279J39_124_314_n1560) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1164 ( .A(
        div_DP_OP_279J39_124_314_n2098), .B(div_DP_OP_279J39_124_314_n1906), 
        .CI(div_DP_OP_279J39_124_314_n1970), .CO(
        div_DP_OP_279J39_124_314_n1557), .S(div_DP_OP_279J39_124_314_n1558) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1163 ( .A(
        div_DP_OP_279J39_124_314_n2034), .B(div_DP_OP_279J39_124_314_n1577), 
        .CI(div_DP_OP_279J39_124_314_n1575), .CO(
        div_DP_OP_279J39_124_314_n1555), .S(div_DP_OP_279J39_124_314_n1556) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1162 ( .A(
        div_DP_OP_279J39_124_314_n1573), .B(div_DP_OP_279J39_124_314_n1562), 
        .CI(div_DP_OP_279J39_124_314_n1558), .CO(
        div_DP_OP_279J39_124_314_n1553), .S(div_DP_OP_279J39_124_314_n1554) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1161 ( .A(
        div_DP_OP_279J39_124_314_n1560), .B(div_DP_OP_279J39_124_314_n1571), 
        .CI(div_DP_OP_279J39_124_314_n1569), .CO(
        div_DP_OP_279J39_124_314_n1551), .S(div_DP_OP_279J39_124_314_n1552) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1160 ( .A(
        div_DP_OP_279J39_124_314_n1556), .B(div_DP_OP_279J39_124_314_n1554), 
        .CI(div_DP_OP_279J39_124_314_n1567), .CO(
        div_DP_OP_279J39_124_314_n1549), .S(div_DP_OP_279J39_124_314_n1550) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1159 ( .A(
        div_DP_OP_279J39_124_314_n1565), .B(div_DP_OP_279J39_124_314_n1552), 
        .CI(div_DP_OP_279J39_124_314_n1550), .CO(
        div_DP_OP_279J39_124_314_n1547), .S(div_DP_OP_279J39_124_314_n1548) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1158 ( .A(div_n_T_51_75_), .B(
        div_DP_OP_279J39_124_314_n1713), .CI(div_DP_OP_279J39_124_314_n2225), 
        .CO(div_DP_OP_279J39_124_314_n1545), .S(div_DP_OP_279J39_124_314_n1546) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1157 ( .A(
        div_DP_OP_279J39_124_314_n2161), .B(div_DP_OP_279J39_124_314_n1777), 
        .CI(div_DP_OP_279J39_124_314_n1841), .CO(
        div_DP_OP_279J39_124_314_n1543), .S(div_DP_OP_279J39_124_314_n1544) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1156 ( .A(
        div_DP_OP_279J39_124_314_n2097), .B(div_DP_OP_279J39_124_314_n1905), 
        .CI(div_DP_OP_279J39_124_314_n1969), .CO(
        div_DP_OP_279J39_124_314_n1541), .S(div_DP_OP_279J39_124_314_n1542) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1155 ( .A(
        div_DP_OP_279J39_124_314_n2033), .B(div_DP_OP_279J39_124_314_n1561), 
        .CI(div_DP_OP_279J39_124_314_n1559), .CO(
        div_DP_OP_279J39_124_314_n1539), .S(div_DP_OP_279J39_124_314_n1540) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1154 ( .A(
        div_DP_OP_279J39_124_314_n1557), .B(div_DP_OP_279J39_124_314_n1546), 
        .CI(div_DP_OP_279J39_124_314_n1542), .CO(
        div_DP_OP_279J39_124_314_n1537), .S(div_DP_OP_279J39_124_314_n1538) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1153 ( .A(
        div_DP_OP_279J39_124_314_n1544), .B(div_DP_OP_279J39_124_314_n1555), 
        .CI(div_DP_OP_279J39_124_314_n1553), .CO(
        div_DP_OP_279J39_124_314_n1535), .S(div_DP_OP_279J39_124_314_n1536) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1152 ( .A(
        div_DP_OP_279J39_124_314_n1540), .B(div_DP_OP_279J39_124_314_n1538), 
        .CI(div_DP_OP_279J39_124_314_n1551), .CO(
        div_DP_OP_279J39_124_314_n1533), .S(div_DP_OP_279J39_124_314_n1534) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1151 ( .A(
        div_DP_OP_279J39_124_314_n1536), .B(div_DP_OP_279J39_124_314_n1549), 
        .CI(div_DP_OP_279J39_124_314_n1534), .CO(
        div_DP_OP_279J39_124_314_n1531), .S(div_DP_OP_279J39_124_314_n1532) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1150 ( .A(div_n_T_51_76_), .B(
        div_DP_OP_279J39_124_314_n1712), .CI(div_DP_OP_279J39_124_314_n2224), 
        .CO(div_DP_OP_279J39_124_314_n1529), .S(div_DP_OP_279J39_124_314_n1530) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1149 ( .A(
        div_DP_OP_279J39_124_314_n2160), .B(div_DP_OP_279J39_124_314_n1776), 
        .CI(div_DP_OP_279J39_124_314_n1840), .CO(
        div_DP_OP_279J39_124_314_n1527), .S(div_DP_OP_279J39_124_314_n1528) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1148 ( .A(
        div_DP_OP_279J39_124_314_n2096), .B(div_DP_OP_279J39_124_314_n1904), 
        .CI(div_DP_OP_279J39_124_314_n1968), .CO(
        div_DP_OP_279J39_124_314_n1525), .S(div_DP_OP_279J39_124_314_n1526) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1147 ( .A(
        div_DP_OP_279J39_124_314_n2032), .B(div_DP_OP_279J39_124_314_n1545), 
        .CI(div_DP_OP_279J39_124_314_n1543), .CO(
        div_DP_OP_279J39_124_314_n1523), .S(div_DP_OP_279J39_124_314_n1524) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1146 ( .A(
        div_DP_OP_279J39_124_314_n1541), .B(div_DP_OP_279J39_124_314_n1530), 
        .CI(div_DP_OP_279J39_124_314_n1526), .CO(
        div_DP_OP_279J39_124_314_n1521), .S(div_DP_OP_279J39_124_314_n1522) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1145 ( .A(
        div_DP_OP_279J39_124_314_n1528), .B(div_DP_OP_279J39_124_314_n1539), 
        .CI(div_DP_OP_279J39_124_314_n1537), .CO(
        div_DP_OP_279J39_124_314_n1519), .S(div_DP_OP_279J39_124_314_n1520) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1144 ( .A(
        div_DP_OP_279J39_124_314_n1524), .B(div_DP_OP_279J39_124_314_n1522), 
        .CI(div_DP_OP_279J39_124_314_n1535), .CO(
        div_DP_OP_279J39_124_314_n1517), .S(div_DP_OP_279J39_124_314_n1518) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1143 ( .A(
        div_DP_OP_279J39_124_314_n1520), .B(div_DP_OP_279J39_124_314_n1533), 
        .CI(div_DP_OP_279J39_124_314_n1518), .CO(
        div_DP_OP_279J39_124_314_n1515), .S(div_DP_OP_279J39_124_314_n1516) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1142 ( .A(div_n_T_51_77_), .B(
        div_DP_OP_279J39_124_314_n1711), .CI(div_DP_OP_279J39_124_314_n2223), 
        .CO(div_DP_OP_279J39_124_314_n1513), .S(div_DP_OP_279J39_124_314_n1514) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1141 ( .A(
        div_DP_OP_279J39_124_314_n2159), .B(div_DP_OP_279J39_124_314_n1775), 
        .CI(div_DP_OP_279J39_124_314_n1839), .CO(
        div_DP_OP_279J39_124_314_n1511), .S(div_DP_OP_279J39_124_314_n1512) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1140 ( .A(
        div_DP_OP_279J39_124_314_n2095), .B(div_DP_OP_279J39_124_314_n1903), 
        .CI(div_DP_OP_279J39_124_314_n1967), .CO(
        div_DP_OP_279J39_124_314_n1509), .S(div_DP_OP_279J39_124_314_n1510) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1139 ( .A(
        div_DP_OP_279J39_124_314_n2031), .B(div_DP_OP_279J39_124_314_n1529), 
        .CI(div_DP_OP_279J39_124_314_n1527), .CO(
        div_DP_OP_279J39_124_314_n1507), .S(div_DP_OP_279J39_124_314_n1508) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1138 ( .A(
        div_DP_OP_279J39_124_314_n1525), .B(div_DP_OP_279J39_124_314_n1514), 
        .CI(div_DP_OP_279J39_124_314_n1510), .CO(
        div_DP_OP_279J39_124_314_n1505), .S(div_DP_OP_279J39_124_314_n1506) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1137 ( .A(
        div_DP_OP_279J39_124_314_n1512), .B(div_DP_OP_279J39_124_314_n1523), 
        .CI(div_DP_OP_279J39_124_314_n1521), .CO(
        div_DP_OP_279J39_124_314_n1503), .S(div_DP_OP_279J39_124_314_n1504) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1136 ( .A(
        div_DP_OP_279J39_124_314_n1508), .B(div_DP_OP_279J39_124_314_n1506), 
        .CI(div_DP_OP_279J39_124_314_n1519), .CO(
        div_DP_OP_279J39_124_314_n1501), .S(div_DP_OP_279J39_124_314_n1502) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1135 ( .A(
        div_DP_OP_279J39_124_314_n1504), .B(div_DP_OP_279J39_124_314_n1517), 
        .CI(div_DP_OP_279J39_124_314_n1502), .CO(
        div_DP_OP_279J39_124_314_n1499), .S(div_DP_OP_279J39_124_314_n1500) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1134 ( .A(div_n_T_51_78_), .B(
        div_DP_OP_279J39_124_314_n1710), .CI(div_DP_OP_279J39_124_314_n2222), 
        .CO(div_DP_OP_279J39_124_314_n1497), .S(div_DP_OP_279J39_124_314_n1498) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1133 ( .A(
        div_DP_OP_279J39_124_314_n2158), .B(div_DP_OP_279J39_124_314_n1774), 
        .CI(div_DP_OP_279J39_124_314_n1838), .CO(
        div_DP_OP_279J39_124_314_n1495), .S(div_DP_OP_279J39_124_314_n1496) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1132 ( .A(
        div_DP_OP_279J39_124_314_n2094), .B(div_DP_OP_279J39_124_314_n1902), 
        .CI(div_DP_OP_279J39_124_314_n1966), .CO(
        div_DP_OP_279J39_124_314_n1493), .S(div_DP_OP_279J39_124_314_n1494) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1131 ( .A(
        div_DP_OP_279J39_124_314_n2030), .B(div_DP_OP_279J39_124_314_n1513), 
        .CI(div_DP_OP_279J39_124_314_n1511), .CO(
        div_DP_OP_279J39_124_314_n1491), .S(div_DP_OP_279J39_124_314_n1492) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1130 ( .A(
        div_DP_OP_279J39_124_314_n1509), .B(div_DP_OP_279J39_124_314_n1498), 
        .CI(div_DP_OP_279J39_124_314_n1494), .CO(
        div_DP_OP_279J39_124_314_n1489), .S(div_DP_OP_279J39_124_314_n1490) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1129 ( .A(
        div_DP_OP_279J39_124_314_n1496), .B(div_DP_OP_279J39_124_314_n1507), 
        .CI(div_DP_OP_279J39_124_314_n1505), .CO(
        div_DP_OP_279J39_124_314_n1487), .S(div_DP_OP_279J39_124_314_n1488) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1128 ( .A(
        div_DP_OP_279J39_124_314_n1492), .B(div_DP_OP_279J39_124_314_n1490), 
        .CI(div_DP_OP_279J39_124_314_n1503), .CO(
        div_DP_OP_279J39_124_314_n1485), .S(div_DP_OP_279J39_124_314_n1486) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1127 ( .A(
        div_DP_OP_279J39_124_314_n1488), .B(div_DP_OP_279J39_124_314_n1501), 
        .CI(div_DP_OP_279J39_124_314_n1486), .CO(
        div_DP_OP_279J39_124_314_n1483), .S(div_DP_OP_279J39_124_314_n1484) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1126 ( .A(div_n_T_51_79_), .B(
        div_DP_OP_279J39_124_314_n1709), .CI(div_DP_OP_279J39_124_314_n2221), 
        .CO(div_DP_OP_279J39_124_314_n1481), .S(div_DP_OP_279J39_124_314_n1482) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1125 ( .A(
        div_DP_OP_279J39_124_314_n2157), .B(div_DP_OP_279J39_124_314_n1773), 
        .CI(div_DP_OP_279J39_124_314_n1837), .CO(
        div_DP_OP_279J39_124_314_n1479), .S(div_DP_OP_279J39_124_314_n1480) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1124 ( .A(
        div_DP_OP_279J39_124_314_n2093), .B(div_DP_OP_279J39_124_314_n1901), 
        .CI(div_DP_OP_279J39_124_314_n1965), .CO(
        div_DP_OP_279J39_124_314_n1477), .S(div_DP_OP_279J39_124_314_n1478) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1123 ( .A(
        div_DP_OP_279J39_124_314_n2029), .B(div_DP_OP_279J39_124_314_n1497), 
        .CI(div_DP_OP_279J39_124_314_n1495), .CO(
        div_DP_OP_279J39_124_314_n1475), .S(div_DP_OP_279J39_124_314_n1476) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1122 ( .A(
        div_DP_OP_279J39_124_314_n1493), .B(div_DP_OP_279J39_124_314_n1482), 
        .CI(div_DP_OP_279J39_124_314_n1478), .CO(
        div_DP_OP_279J39_124_314_n1473), .S(div_DP_OP_279J39_124_314_n1474) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1121 ( .A(
        div_DP_OP_279J39_124_314_n1480), .B(div_DP_OP_279J39_124_314_n1491), 
        .CI(div_DP_OP_279J39_124_314_n1489), .CO(
        div_DP_OP_279J39_124_314_n1471), .S(div_DP_OP_279J39_124_314_n1472) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1120 ( .A(
        div_DP_OP_279J39_124_314_n1476), .B(div_DP_OP_279J39_124_314_n1474), 
        .CI(div_DP_OP_279J39_124_314_n1487), .CO(
        div_DP_OP_279J39_124_314_n1469), .S(div_DP_OP_279J39_124_314_n1470) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1119 ( .A(
        div_DP_OP_279J39_124_314_n1472), .B(div_DP_OP_279J39_124_314_n1485), 
        .CI(div_DP_OP_279J39_124_314_n1470), .CO(
        div_DP_OP_279J39_124_314_n1467), .S(div_DP_OP_279J39_124_314_n1468) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1118 ( .A(div_n_T_51_80_), .B(
        div_DP_OP_279J39_124_314_n1708), .CI(div_DP_OP_279J39_124_314_n2220), 
        .CO(div_DP_OP_279J39_124_314_n1465), .S(div_DP_OP_279J39_124_314_n1466) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1117 ( .A(
        div_DP_OP_279J39_124_314_n2156), .B(div_DP_OP_279J39_124_314_n1772), 
        .CI(div_DP_OP_279J39_124_314_n1836), .CO(
        div_DP_OP_279J39_124_314_n1463), .S(div_DP_OP_279J39_124_314_n1464) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1116 ( .A(
        div_DP_OP_279J39_124_314_n2092), .B(div_DP_OP_279J39_124_314_n1900), 
        .CI(div_DP_OP_279J39_124_314_n1964), .CO(
        div_DP_OP_279J39_124_314_n1461), .S(div_DP_OP_279J39_124_314_n1462) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1115 ( .A(
        div_DP_OP_279J39_124_314_n2028), .B(div_DP_OP_279J39_124_314_n1481), 
        .CI(div_DP_OP_279J39_124_314_n1479), .CO(
        div_DP_OP_279J39_124_314_n1459), .S(div_DP_OP_279J39_124_314_n1460) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1114 ( .A(
        div_DP_OP_279J39_124_314_n1477), .B(div_DP_OP_279J39_124_314_n1466), 
        .CI(div_DP_OP_279J39_124_314_n1462), .CO(
        div_DP_OP_279J39_124_314_n1457), .S(div_DP_OP_279J39_124_314_n1458) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1113 ( .A(
        div_DP_OP_279J39_124_314_n1464), .B(div_DP_OP_279J39_124_314_n1475), 
        .CI(div_DP_OP_279J39_124_314_n1473), .CO(
        div_DP_OP_279J39_124_314_n1455), .S(div_DP_OP_279J39_124_314_n1456) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1112 ( .A(
        div_DP_OP_279J39_124_314_n1460), .B(div_DP_OP_279J39_124_314_n1458), 
        .CI(div_DP_OP_279J39_124_314_n1471), .CO(
        div_DP_OP_279J39_124_314_n1453), .S(div_DP_OP_279J39_124_314_n1454) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1111 ( .A(
        div_DP_OP_279J39_124_314_n1456), .B(div_DP_OP_279J39_124_314_n1469), 
        .CI(div_DP_OP_279J39_124_314_n1454), .CO(
        div_DP_OP_279J39_124_314_n1451), .S(div_DP_OP_279J39_124_314_n1452) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1110 ( .A(div_n_T_51_81_), .B(
        div_DP_OP_279J39_124_314_n1707), .CI(div_DP_OP_279J39_124_314_n2219), 
        .CO(div_DP_OP_279J39_124_314_n1449), .S(div_DP_OP_279J39_124_314_n1450) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1109 ( .A(
        div_DP_OP_279J39_124_314_n2155), .B(div_DP_OP_279J39_124_314_n1771), 
        .CI(div_DP_OP_279J39_124_314_n1835), .CO(
        div_DP_OP_279J39_124_314_n1447), .S(div_DP_OP_279J39_124_314_n1448) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1108 ( .A(
        div_DP_OP_279J39_124_314_n2091), .B(div_DP_OP_279J39_124_314_n1899), 
        .CI(div_DP_OP_279J39_124_314_n1963), .CO(
        div_DP_OP_279J39_124_314_n1445), .S(div_DP_OP_279J39_124_314_n1446) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1107 ( .A(
        div_DP_OP_279J39_124_314_n2027), .B(div_DP_OP_279J39_124_314_n1465), 
        .CI(div_DP_OP_279J39_124_314_n1463), .CO(
        div_DP_OP_279J39_124_314_n1443), .S(div_DP_OP_279J39_124_314_n1444) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1106 ( .A(
        div_DP_OP_279J39_124_314_n1461), .B(div_DP_OP_279J39_124_314_n1450), 
        .CI(div_DP_OP_279J39_124_314_n1446), .CO(
        div_DP_OP_279J39_124_314_n1441), .S(div_DP_OP_279J39_124_314_n1442) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1105 ( .A(
        div_DP_OP_279J39_124_314_n1448), .B(div_DP_OP_279J39_124_314_n1459), 
        .CI(div_DP_OP_279J39_124_314_n1457), .CO(
        div_DP_OP_279J39_124_314_n1439), .S(div_DP_OP_279J39_124_314_n1440) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1104 ( .A(
        div_DP_OP_279J39_124_314_n1444), .B(div_DP_OP_279J39_124_314_n1442), 
        .CI(div_DP_OP_279J39_124_314_n1455), .CO(
        div_DP_OP_279J39_124_314_n1437), .S(div_DP_OP_279J39_124_314_n1438) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1103 ( .A(
        div_DP_OP_279J39_124_314_n1440), .B(div_DP_OP_279J39_124_314_n1453), 
        .CI(div_DP_OP_279J39_124_314_n1438), .CO(
        div_DP_OP_279J39_124_314_n1435), .S(div_DP_OP_279J39_124_314_n1436) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1102 ( .A(div_n_T_51_82_), .B(
        div_DP_OP_279J39_124_314_n1706), .CI(div_DP_OP_279J39_124_314_n2218), 
        .CO(div_DP_OP_279J39_124_314_n1433), .S(div_DP_OP_279J39_124_314_n1434) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1101 ( .A(
        div_DP_OP_279J39_124_314_n2154), .B(div_DP_OP_279J39_124_314_n1770), 
        .CI(div_DP_OP_279J39_124_314_n1834), .CO(
        div_DP_OP_279J39_124_314_n1431), .S(div_DP_OP_279J39_124_314_n1432) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1100 ( .A(
        div_DP_OP_279J39_124_314_n2090), .B(div_DP_OP_279J39_124_314_n1898), 
        .CI(div_DP_OP_279J39_124_314_n1962), .CO(
        div_DP_OP_279J39_124_314_n1429), .S(div_DP_OP_279J39_124_314_n1430) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1099 ( .A(
        div_DP_OP_279J39_124_314_n2026), .B(div_DP_OP_279J39_124_314_n1449), 
        .CI(div_DP_OP_279J39_124_314_n1447), .CO(
        div_DP_OP_279J39_124_314_n1427), .S(div_DP_OP_279J39_124_314_n1428) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1098 ( .A(
        div_DP_OP_279J39_124_314_n1445), .B(div_DP_OP_279J39_124_314_n1434), 
        .CI(div_DP_OP_279J39_124_314_n1430), .CO(
        div_DP_OP_279J39_124_314_n1425), .S(div_DP_OP_279J39_124_314_n1426) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1097 ( .A(
        div_DP_OP_279J39_124_314_n1432), .B(div_DP_OP_279J39_124_314_n1443), 
        .CI(div_DP_OP_279J39_124_314_n1441), .CO(
        div_DP_OP_279J39_124_314_n1423), .S(div_DP_OP_279J39_124_314_n1424) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1096 ( .A(
        div_DP_OP_279J39_124_314_n1428), .B(div_DP_OP_279J39_124_314_n1426), 
        .CI(div_DP_OP_279J39_124_314_n1439), .CO(
        div_DP_OP_279J39_124_314_n1421), .S(div_DP_OP_279J39_124_314_n1422) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1095 ( .A(
        div_DP_OP_279J39_124_314_n1424), .B(div_DP_OP_279J39_124_314_n1437), 
        .CI(div_DP_OP_279J39_124_314_n1422), .CO(
        div_DP_OP_279J39_124_314_n1419), .S(div_DP_OP_279J39_124_314_n1420) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1094 ( .A(div_n_T_51_83_), .B(
        div_DP_OP_279J39_124_314_n1705), .CI(div_DP_OP_279J39_124_314_n2217), 
        .CO(div_DP_OP_279J39_124_314_n1417), .S(div_DP_OP_279J39_124_314_n1418) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1093 ( .A(
        div_DP_OP_279J39_124_314_n2153), .B(div_DP_OP_279J39_124_314_n1769), 
        .CI(div_DP_OP_279J39_124_314_n1833), .CO(
        div_DP_OP_279J39_124_314_n1415), .S(div_DP_OP_279J39_124_314_n1416) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1092 ( .A(
        div_DP_OP_279J39_124_314_n2089), .B(div_DP_OP_279J39_124_314_n1897), 
        .CI(div_DP_OP_279J39_124_314_n1961), .CO(
        div_DP_OP_279J39_124_314_n1413), .S(div_DP_OP_279J39_124_314_n1414) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1091 ( .A(
        div_DP_OP_279J39_124_314_n2025), .B(div_DP_OP_279J39_124_314_n1433), 
        .CI(div_DP_OP_279J39_124_314_n1431), .CO(
        div_DP_OP_279J39_124_314_n1411), .S(div_DP_OP_279J39_124_314_n1412) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1090 ( .A(
        div_DP_OP_279J39_124_314_n1429), .B(div_DP_OP_279J39_124_314_n1418), 
        .CI(div_DP_OP_279J39_124_314_n1414), .CO(
        div_DP_OP_279J39_124_314_n1409), .S(div_DP_OP_279J39_124_314_n1410) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1089 ( .A(
        div_DP_OP_279J39_124_314_n1416), .B(div_DP_OP_279J39_124_314_n1427), 
        .CI(div_DP_OP_279J39_124_314_n1425), .CO(
        div_DP_OP_279J39_124_314_n1407), .S(div_DP_OP_279J39_124_314_n1408) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1088 ( .A(
        div_DP_OP_279J39_124_314_n1412), .B(div_DP_OP_279J39_124_314_n1410), 
        .CI(div_DP_OP_279J39_124_314_n1423), .CO(
        div_DP_OP_279J39_124_314_n1405), .S(div_DP_OP_279J39_124_314_n1406) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1087 ( .A(
        div_DP_OP_279J39_124_314_n1408), .B(div_DP_OP_279J39_124_314_n1421), 
        .CI(div_DP_OP_279J39_124_314_n1406), .CO(
        div_DP_OP_279J39_124_314_n1403), .S(div_DP_OP_279J39_124_314_n1404) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1086 ( .A(div_n_T_51_84_), .B(
        div_DP_OP_279J39_124_314_n1704), .CI(div_DP_OP_279J39_124_314_n2216), 
        .CO(div_DP_OP_279J39_124_314_n1401), .S(div_DP_OP_279J39_124_314_n1402) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1085 ( .A(
        div_DP_OP_279J39_124_314_n2152), .B(div_DP_OP_279J39_124_314_n1768), 
        .CI(div_DP_OP_279J39_124_314_n1832), .CO(
        div_DP_OP_279J39_124_314_n1399), .S(div_DP_OP_279J39_124_314_n1400) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1084 ( .A(
        div_DP_OP_279J39_124_314_n2088), .B(div_DP_OP_279J39_124_314_n1896), 
        .CI(div_DP_OP_279J39_124_314_n1960), .CO(
        div_DP_OP_279J39_124_314_n1397), .S(div_DP_OP_279J39_124_314_n1398) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1083 ( .A(
        div_DP_OP_279J39_124_314_n2024), .B(div_DP_OP_279J39_124_314_n1417), 
        .CI(div_DP_OP_279J39_124_314_n1415), .CO(
        div_DP_OP_279J39_124_314_n1395), .S(div_DP_OP_279J39_124_314_n1396) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1082 ( .A(
        div_DP_OP_279J39_124_314_n1413), .B(div_DP_OP_279J39_124_314_n1402), 
        .CI(div_DP_OP_279J39_124_314_n1398), .CO(
        div_DP_OP_279J39_124_314_n1393), .S(div_DP_OP_279J39_124_314_n1394) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1081 ( .A(
        div_DP_OP_279J39_124_314_n1400), .B(div_DP_OP_279J39_124_314_n1411), 
        .CI(div_DP_OP_279J39_124_314_n1409), .CO(
        div_DP_OP_279J39_124_314_n1391), .S(div_DP_OP_279J39_124_314_n1392) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1080 ( .A(
        div_DP_OP_279J39_124_314_n1396), .B(div_DP_OP_279J39_124_314_n1394), 
        .CI(div_DP_OP_279J39_124_314_n1407), .CO(
        div_DP_OP_279J39_124_314_n1389), .S(div_DP_OP_279J39_124_314_n1390) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1079 ( .A(
        div_DP_OP_279J39_124_314_n1392), .B(div_DP_OP_279J39_124_314_n1405), 
        .CI(div_DP_OP_279J39_124_314_n1390), .CO(
        div_DP_OP_279J39_124_314_n1387), .S(div_DP_OP_279J39_124_314_n1388) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1078 ( .A(div_n_T_51_85_), .B(
        div_DP_OP_279J39_124_314_n1703), .CI(div_DP_OP_279J39_124_314_n2215), 
        .CO(div_DP_OP_279J39_124_314_n1385), .S(div_DP_OP_279J39_124_314_n1386) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1077 ( .A(
        div_DP_OP_279J39_124_314_n2151), .B(div_DP_OP_279J39_124_314_n1767), 
        .CI(div_DP_OP_279J39_124_314_n1831), .CO(
        div_DP_OP_279J39_124_314_n1383), .S(div_DP_OP_279J39_124_314_n1384) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1076 ( .A(
        div_DP_OP_279J39_124_314_n2087), .B(div_DP_OP_279J39_124_314_n1895), 
        .CI(div_DP_OP_279J39_124_314_n1959), .CO(
        div_DP_OP_279J39_124_314_n1381), .S(div_DP_OP_279J39_124_314_n1382) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1075 ( .A(
        div_DP_OP_279J39_124_314_n2023), .B(div_DP_OP_279J39_124_314_n1401), 
        .CI(div_DP_OP_279J39_124_314_n1399), .CO(
        div_DP_OP_279J39_124_314_n1379), .S(div_DP_OP_279J39_124_314_n1380) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1074 ( .A(
        div_DP_OP_279J39_124_314_n1397), .B(div_DP_OP_279J39_124_314_n1386), 
        .CI(div_DP_OP_279J39_124_314_n1382), .CO(
        div_DP_OP_279J39_124_314_n1377), .S(div_DP_OP_279J39_124_314_n1378) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1073 ( .A(
        div_DP_OP_279J39_124_314_n1384), .B(div_DP_OP_279J39_124_314_n1395), 
        .CI(div_DP_OP_279J39_124_314_n1393), .CO(
        div_DP_OP_279J39_124_314_n1375), .S(div_DP_OP_279J39_124_314_n1376) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1072 ( .A(
        div_DP_OP_279J39_124_314_n1380), .B(div_DP_OP_279J39_124_314_n1378), 
        .CI(div_DP_OP_279J39_124_314_n1391), .CO(
        div_DP_OP_279J39_124_314_n1373), .S(div_DP_OP_279J39_124_314_n1374) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1071 ( .A(
        div_DP_OP_279J39_124_314_n1376), .B(div_DP_OP_279J39_124_314_n1389), 
        .CI(div_DP_OP_279J39_124_314_n1374), .CO(
        div_DP_OP_279J39_124_314_n1371), .S(div_DP_OP_279J39_124_314_n1372) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1070 ( .A(div_n_T_51_86_), .B(
        div_DP_OP_279J39_124_314_n1702), .CI(div_DP_OP_279J39_124_314_n2214), 
        .CO(div_DP_OP_279J39_124_314_n1369), .S(div_DP_OP_279J39_124_314_n1370) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1069 ( .A(
        div_DP_OP_279J39_124_314_n2150), .B(div_DP_OP_279J39_124_314_n1766), 
        .CI(div_DP_OP_279J39_124_314_n1830), .CO(
        div_DP_OP_279J39_124_314_n1367), .S(div_DP_OP_279J39_124_314_n1368) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1068 ( .A(
        div_DP_OP_279J39_124_314_n2086), .B(div_DP_OP_279J39_124_314_n1894), 
        .CI(div_DP_OP_279J39_124_314_n1958), .CO(
        div_DP_OP_279J39_124_314_n1365), .S(div_DP_OP_279J39_124_314_n1366) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1067 ( .A(
        div_DP_OP_279J39_124_314_n2022), .B(div_DP_OP_279J39_124_314_n1385), 
        .CI(div_DP_OP_279J39_124_314_n1383), .CO(
        div_DP_OP_279J39_124_314_n1363), .S(div_DP_OP_279J39_124_314_n1364) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1066 ( .A(
        div_DP_OP_279J39_124_314_n1381), .B(div_DP_OP_279J39_124_314_n1370), 
        .CI(div_DP_OP_279J39_124_314_n1366), .CO(
        div_DP_OP_279J39_124_314_n1361), .S(div_DP_OP_279J39_124_314_n1362) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1065 ( .A(
        div_DP_OP_279J39_124_314_n1368), .B(div_DP_OP_279J39_124_314_n1379), 
        .CI(div_DP_OP_279J39_124_314_n1377), .CO(
        div_DP_OP_279J39_124_314_n1359), .S(div_DP_OP_279J39_124_314_n1360) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1064 ( .A(
        div_DP_OP_279J39_124_314_n1364), .B(div_DP_OP_279J39_124_314_n1362), 
        .CI(div_DP_OP_279J39_124_314_n1375), .CO(
        div_DP_OP_279J39_124_314_n1357), .S(div_DP_OP_279J39_124_314_n1358) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1063 ( .A(
        div_DP_OP_279J39_124_314_n1360), .B(div_DP_OP_279J39_124_314_n1373), 
        .CI(div_DP_OP_279J39_124_314_n1358), .CO(
        div_DP_OP_279J39_124_314_n1355), .S(div_DP_OP_279J39_124_314_n1356) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1062 ( .A(div_n_T_51_87_), .B(
        div_DP_OP_279J39_124_314_n1701), .CI(div_DP_OP_279J39_124_314_n2213), 
        .CO(div_DP_OP_279J39_124_314_n1353), .S(div_DP_OP_279J39_124_314_n1354) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1061 ( .A(
        div_DP_OP_279J39_124_314_n2149), .B(div_DP_OP_279J39_124_314_n1765), 
        .CI(div_DP_OP_279J39_124_314_n1829), .CO(
        div_DP_OP_279J39_124_314_n1351), .S(div_DP_OP_279J39_124_314_n1352) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1060 ( .A(
        div_DP_OP_279J39_124_314_n2085), .B(div_DP_OP_279J39_124_314_n1893), 
        .CI(div_DP_OP_279J39_124_314_n1957), .CO(
        div_DP_OP_279J39_124_314_n1349), .S(div_DP_OP_279J39_124_314_n1350) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1059 ( .A(
        div_DP_OP_279J39_124_314_n2021), .B(div_DP_OP_279J39_124_314_n1369), 
        .CI(div_DP_OP_279J39_124_314_n1367), .CO(
        div_DP_OP_279J39_124_314_n1347), .S(div_DP_OP_279J39_124_314_n1348) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1058 ( .A(
        div_DP_OP_279J39_124_314_n1365), .B(div_DP_OP_279J39_124_314_n1354), 
        .CI(div_DP_OP_279J39_124_314_n1350), .CO(
        div_DP_OP_279J39_124_314_n1345), .S(div_DP_OP_279J39_124_314_n1346) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1057 ( .A(
        div_DP_OP_279J39_124_314_n1352), .B(div_DP_OP_279J39_124_314_n1363), 
        .CI(div_DP_OP_279J39_124_314_n1361), .CO(
        div_DP_OP_279J39_124_314_n1343), .S(div_DP_OP_279J39_124_314_n1344) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1056 ( .A(
        div_DP_OP_279J39_124_314_n1348), .B(div_DP_OP_279J39_124_314_n1346), 
        .CI(div_DP_OP_279J39_124_314_n1359), .CO(
        div_DP_OP_279J39_124_314_n1341), .S(div_DP_OP_279J39_124_314_n1342) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1055 ( .A(
        div_DP_OP_279J39_124_314_n1344), .B(div_DP_OP_279J39_124_314_n1357), 
        .CI(div_DP_OP_279J39_124_314_n1342), .CO(
        div_DP_OP_279J39_124_314_n1339), .S(div_DP_OP_279J39_124_314_n1340) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1054 ( .A(div_n_T_51_88_), .B(
        div_DP_OP_279J39_124_314_n1700), .CI(div_DP_OP_279J39_124_314_n2212), 
        .CO(div_DP_OP_279J39_124_314_n1337), .S(div_DP_OP_279J39_124_314_n1338) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1053 ( .A(
        div_DP_OP_279J39_124_314_n2148), .B(div_DP_OP_279J39_124_314_n1764), 
        .CI(div_DP_OP_279J39_124_314_n1828), .CO(
        div_DP_OP_279J39_124_314_n1335), .S(div_DP_OP_279J39_124_314_n1336) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1052 ( .A(
        div_DP_OP_279J39_124_314_n2084), .B(div_DP_OP_279J39_124_314_n1892), 
        .CI(div_DP_OP_279J39_124_314_n1956), .CO(
        div_DP_OP_279J39_124_314_n1333), .S(div_DP_OP_279J39_124_314_n1334) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1051 ( .A(
        div_DP_OP_279J39_124_314_n2020), .B(div_DP_OP_279J39_124_314_n1353), 
        .CI(div_DP_OP_279J39_124_314_n1351), .CO(
        div_DP_OP_279J39_124_314_n1331), .S(div_DP_OP_279J39_124_314_n1332) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1050 ( .A(
        div_DP_OP_279J39_124_314_n1349), .B(div_DP_OP_279J39_124_314_n1338), 
        .CI(div_DP_OP_279J39_124_314_n1334), .CO(
        div_DP_OP_279J39_124_314_n1329), .S(div_DP_OP_279J39_124_314_n1330) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1049 ( .A(
        div_DP_OP_279J39_124_314_n1336), .B(div_DP_OP_279J39_124_314_n1347), 
        .CI(div_DP_OP_279J39_124_314_n1345), .CO(
        div_DP_OP_279J39_124_314_n1327), .S(div_DP_OP_279J39_124_314_n1328) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1048 ( .A(
        div_DP_OP_279J39_124_314_n1332), .B(div_DP_OP_279J39_124_314_n1330), 
        .CI(div_DP_OP_279J39_124_314_n1343), .CO(
        div_DP_OP_279J39_124_314_n1325), .S(div_DP_OP_279J39_124_314_n1326) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1047 ( .A(
        div_DP_OP_279J39_124_314_n1328), .B(div_DP_OP_279J39_124_314_n1341), 
        .CI(div_DP_OP_279J39_124_314_n1326), .CO(
        div_DP_OP_279J39_124_314_n1323), .S(div_DP_OP_279J39_124_314_n1324) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1046 ( .A(div_n_T_51_89_), .B(
        div_DP_OP_279J39_124_314_n1699), .CI(div_DP_OP_279J39_124_314_n2211), 
        .CO(div_DP_OP_279J39_124_314_n1321), .S(div_DP_OP_279J39_124_314_n1322) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1045 ( .A(
        div_DP_OP_279J39_124_314_n2147), .B(div_DP_OP_279J39_124_314_n1763), 
        .CI(div_DP_OP_279J39_124_314_n1827), .CO(
        div_DP_OP_279J39_124_314_n1319), .S(div_DP_OP_279J39_124_314_n1320) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1044 ( .A(
        div_DP_OP_279J39_124_314_n2083), .B(div_DP_OP_279J39_124_314_n1891), 
        .CI(div_DP_OP_279J39_124_314_n1955), .CO(
        div_DP_OP_279J39_124_314_n1317), .S(div_DP_OP_279J39_124_314_n1318) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1043 ( .A(
        div_DP_OP_279J39_124_314_n2019), .B(div_DP_OP_279J39_124_314_n1337), 
        .CI(div_DP_OP_279J39_124_314_n1335), .CO(
        div_DP_OP_279J39_124_314_n1315), .S(div_DP_OP_279J39_124_314_n1316) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1042 ( .A(
        div_DP_OP_279J39_124_314_n1333), .B(div_DP_OP_279J39_124_314_n1322), 
        .CI(div_DP_OP_279J39_124_314_n1318), .CO(
        div_DP_OP_279J39_124_314_n1313), .S(div_DP_OP_279J39_124_314_n1314) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1041 ( .A(
        div_DP_OP_279J39_124_314_n1320), .B(div_DP_OP_279J39_124_314_n1331), 
        .CI(div_DP_OP_279J39_124_314_n1329), .CO(
        div_DP_OP_279J39_124_314_n1311), .S(div_DP_OP_279J39_124_314_n1312) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1040 ( .A(
        div_DP_OP_279J39_124_314_n1316), .B(div_DP_OP_279J39_124_314_n1314), 
        .CI(div_DP_OP_279J39_124_314_n1327), .CO(
        div_DP_OP_279J39_124_314_n1309), .S(div_DP_OP_279J39_124_314_n1310) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1039 ( .A(
        div_DP_OP_279J39_124_314_n1312), .B(div_DP_OP_279J39_124_314_n1325), 
        .CI(div_DP_OP_279J39_124_314_n1310), .CO(
        div_DP_OP_279J39_124_314_n1307), .S(div_DP_OP_279J39_124_314_n1308) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1038 ( .A(div_n_T_51_90_), .B(
        div_DP_OP_279J39_124_314_n1698), .CI(div_DP_OP_279J39_124_314_n2210), 
        .CO(div_DP_OP_279J39_124_314_n1305), .S(div_DP_OP_279J39_124_314_n1306) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1037 ( .A(
        div_DP_OP_279J39_124_314_n2146), .B(div_DP_OP_279J39_124_314_n1762), 
        .CI(div_DP_OP_279J39_124_314_n1826), .CO(
        div_DP_OP_279J39_124_314_n1303), .S(div_DP_OP_279J39_124_314_n1304) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1036 ( .A(
        div_DP_OP_279J39_124_314_n2082), .B(div_DP_OP_279J39_124_314_n1890), 
        .CI(div_DP_OP_279J39_124_314_n1954), .CO(
        div_DP_OP_279J39_124_314_n1301), .S(div_DP_OP_279J39_124_314_n1302) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1035 ( .A(
        div_DP_OP_279J39_124_314_n2018), .B(div_DP_OP_279J39_124_314_n1321), 
        .CI(div_DP_OP_279J39_124_314_n1319), .CO(
        div_DP_OP_279J39_124_314_n1299), .S(div_DP_OP_279J39_124_314_n1300) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1034 ( .A(
        div_DP_OP_279J39_124_314_n1317), .B(div_DP_OP_279J39_124_314_n1306), 
        .CI(div_DP_OP_279J39_124_314_n1302), .CO(
        div_DP_OP_279J39_124_314_n1297), .S(div_DP_OP_279J39_124_314_n1298) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1033 ( .A(
        div_DP_OP_279J39_124_314_n1304), .B(div_DP_OP_279J39_124_314_n1315), 
        .CI(div_DP_OP_279J39_124_314_n1313), .CO(
        div_DP_OP_279J39_124_314_n1295), .S(div_DP_OP_279J39_124_314_n1296) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1032 ( .A(
        div_DP_OP_279J39_124_314_n1300), .B(div_DP_OP_279J39_124_314_n1298), 
        .CI(div_DP_OP_279J39_124_314_n1311), .CO(
        div_DP_OP_279J39_124_314_n1293), .S(div_DP_OP_279J39_124_314_n1294) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1031 ( .A(
        div_DP_OP_279J39_124_314_n1296), .B(div_DP_OP_279J39_124_314_n1309), 
        .CI(div_DP_OP_279J39_124_314_n1294), .CO(
        div_DP_OP_279J39_124_314_n1291), .S(div_DP_OP_279J39_124_314_n1292) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1030 ( .A(div_n_T_51_91_), .B(
        div_DP_OP_279J39_124_314_n1697), .CI(div_DP_OP_279J39_124_314_n2209), 
        .CO(div_DP_OP_279J39_124_314_n1289), .S(div_DP_OP_279J39_124_314_n1290) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1029 ( .A(
        div_DP_OP_279J39_124_314_n2145), .B(div_DP_OP_279J39_124_314_n1761), 
        .CI(div_DP_OP_279J39_124_314_n1825), .CO(
        div_DP_OP_279J39_124_314_n1287), .S(div_DP_OP_279J39_124_314_n1288) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1028 ( .A(
        div_DP_OP_279J39_124_314_n2081), .B(div_DP_OP_279J39_124_314_n1889), 
        .CI(div_DP_OP_279J39_124_314_n1953), .CO(
        div_DP_OP_279J39_124_314_n1285), .S(div_DP_OP_279J39_124_314_n1286) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1027 ( .A(
        div_DP_OP_279J39_124_314_n2017), .B(div_DP_OP_279J39_124_314_n1305), 
        .CI(div_DP_OP_279J39_124_314_n1303), .CO(
        div_DP_OP_279J39_124_314_n1283), .S(div_DP_OP_279J39_124_314_n1284) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1026 ( .A(
        div_DP_OP_279J39_124_314_n1301), .B(div_DP_OP_279J39_124_314_n1290), 
        .CI(div_DP_OP_279J39_124_314_n1286), .CO(
        div_DP_OP_279J39_124_314_n1281), .S(div_DP_OP_279J39_124_314_n1282) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1025 ( .A(
        div_DP_OP_279J39_124_314_n1288), .B(div_DP_OP_279J39_124_314_n1299), 
        .CI(div_DP_OP_279J39_124_314_n1297), .CO(
        div_DP_OP_279J39_124_314_n1279), .S(div_DP_OP_279J39_124_314_n1280) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1024 ( .A(
        div_DP_OP_279J39_124_314_n1284), .B(div_DP_OP_279J39_124_314_n1282), 
        .CI(div_DP_OP_279J39_124_314_n1295), .CO(
        div_DP_OP_279J39_124_314_n1277), .S(div_DP_OP_279J39_124_314_n1278) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1023 ( .A(
        div_DP_OP_279J39_124_314_n1280), .B(div_DP_OP_279J39_124_314_n1293), 
        .CI(div_DP_OP_279J39_124_314_n1278), .CO(
        div_DP_OP_279J39_124_314_n1275), .S(div_DP_OP_279J39_124_314_n1276) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1022 ( .A(div_n_T_51_92_), .B(
        div_DP_OP_279J39_124_314_n1696), .CI(div_DP_OP_279J39_124_314_n2208), 
        .CO(div_DP_OP_279J39_124_314_n1273), .S(div_DP_OP_279J39_124_314_n1274) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1021 ( .A(
        div_DP_OP_279J39_124_314_n2144), .B(div_DP_OP_279J39_124_314_n1760), 
        .CI(div_DP_OP_279J39_124_314_n1824), .CO(
        div_DP_OP_279J39_124_314_n1271), .S(div_DP_OP_279J39_124_314_n1272) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1020 ( .A(
        div_DP_OP_279J39_124_314_n2080), .B(div_DP_OP_279J39_124_314_n1888), 
        .CI(div_DP_OP_279J39_124_314_n1952), .CO(
        div_DP_OP_279J39_124_314_n1269), .S(div_DP_OP_279J39_124_314_n1270) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1019 ( .A(
        div_DP_OP_279J39_124_314_n2016), .B(div_DP_OP_279J39_124_314_n1289), 
        .CI(div_DP_OP_279J39_124_314_n1287), .CO(
        div_DP_OP_279J39_124_314_n1267), .S(div_DP_OP_279J39_124_314_n1268) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1018 ( .A(
        div_DP_OP_279J39_124_314_n1285), .B(div_DP_OP_279J39_124_314_n1274), 
        .CI(div_DP_OP_279J39_124_314_n1270), .CO(
        div_DP_OP_279J39_124_314_n1265), .S(div_DP_OP_279J39_124_314_n1266) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1017 ( .A(
        div_DP_OP_279J39_124_314_n1272), .B(div_DP_OP_279J39_124_314_n1283), 
        .CI(div_DP_OP_279J39_124_314_n1281), .CO(
        div_DP_OP_279J39_124_314_n1263), .S(div_DP_OP_279J39_124_314_n1264) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1016 ( .A(
        div_DP_OP_279J39_124_314_n1268), .B(div_DP_OP_279J39_124_314_n1266), 
        .CI(div_DP_OP_279J39_124_314_n1279), .CO(
        div_DP_OP_279J39_124_314_n1261), .S(div_DP_OP_279J39_124_314_n1262) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1015 ( .A(
        div_DP_OP_279J39_124_314_n1264), .B(div_DP_OP_279J39_124_314_n1277), 
        .CI(div_DP_OP_279J39_124_314_n1262), .CO(
        div_DP_OP_279J39_124_314_n1259), .S(div_DP_OP_279J39_124_314_n1260) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1014 ( .A(div_n_T_51_93_), .B(
        div_DP_OP_279J39_124_314_n1695), .CI(div_DP_OP_279J39_124_314_n2207), 
        .CO(div_DP_OP_279J39_124_314_n1257), .S(div_DP_OP_279J39_124_314_n1258) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1013 ( .A(
        div_DP_OP_279J39_124_314_n2143), .B(div_DP_OP_279J39_124_314_n1759), 
        .CI(div_DP_OP_279J39_124_314_n1823), .CO(
        div_DP_OP_279J39_124_314_n1255), .S(div_DP_OP_279J39_124_314_n1256) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1012 ( .A(
        div_DP_OP_279J39_124_314_n2079), .B(div_DP_OP_279J39_124_314_n1887), 
        .CI(div_DP_OP_279J39_124_314_n1951), .CO(
        div_DP_OP_279J39_124_314_n1253), .S(div_DP_OP_279J39_124_314_n1254) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1011 ( .A(
        div_DP_OP_279J39_124_314_n2015), .B(div_DP_OP_279J39_124_314_n1273), 
        .CI(div_DP_OP_279J39_124_314_n1271), .CO(
        div_DP_OP_279J39_124_314_n1251), .S(div_DP_OP_279J39_124_314_n1252) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1010 ( .A(
        div_DP_OP_279J39_124_314_n1269), .B(div_DP_OP_279J39_124_314_n1258), 
        .CI(div_DP_OP_279J39_124_314_n1254), .CO(
        div_DP_OP_279J39_124_314_n1249), .S(div_DP_OP_279J39_124_314_n1250) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1009 ( .A(
        div_DP_OP_279J39_124_314_n1256), .B(div_DP_OP_279J39_124_314_n1267), 
        .CI(div_DP_OP_279J39_124_314_n1265), .CO(
        div_DP_OP_279J39_124_314_n1247), .S(div_DP_OP_279J39_124_314_n1248) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1008 ( .A(
        div_DP_OP_279J39_124_314_n1252), .B(div_DP_OP_279J39_124_314_n1250), 
        .CI(div_DP_OP_279J39_124_314_n1263), .CO(
        div_DP_OP_279J39_124_314_n1245), .S(div_DP_OP_279J39_124_314_n1246) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1007 ( .A(
        div_DP_OP_279J39_124_314_n1248), .B(div_DP_OP_279J39_124_314_n1261), 
        .CI(div_DP_OP_279J39_124_314_n1246), .CO(
        div_DP_OP_279J39_124_314_n1243), .S(div_DP_OP_279J39_124_314_n1244) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1006 ( .A(div_n_T_51_94_), .B(
        div_DP_OP_279J39_124_314_n1694), .CI(div_DP_OP_279J39_124_314_n2206), 
        .CO(div_DP_OP_279J39_124_314_n1241), .S(div_DP_OP_279J39_124_314_n1242) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1005 ( .A(
        div_DP_OP_279J39_124_314_n2142), .B(div_DP_OP_279J39_124_314_n1758), 
        .CI(div_DP_OP_279J39_124_314_n1822), .CO(
        div_DP_OP_279J39_124_314_n1239), .S(div_DP_OP_279J39_124_314_n1240) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1004 ( .A(
        div_DP_OP_279J39_124_314_n2078), .B(div_DP_OP_279J39_124_314_n1886), 
        .CI(div_DP_OP_279J39_124_314_n1950), .CO(
        div_DP_OP_279J39_124_314_n1237), .S(div_DP_OP_279J39_124_314_n1238) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1003 ( .A(
        div_DP_OP_279J39_124_314_n2014), .B(div_DP_OP_279J39_124_314_n1257), 
        .CI(div_DP_OP_279J39_124_314_n1255), .CO(
        div_DP_OP_279J39_124_314_n1235), .S(div_DP_OP_279J39_124_314_n1236) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1002 ( .A(
        div_DP_OP_279J39_124_314_n1253), .B(div_DP_OP_279J39_124_314_n1242), 
        .CI(div_DP_OP_279J39_124_314_n1238), .CO(
        div_DP_OP_279J39_124_314_n1233), .S(div_DP_OP_279J39_124_314_n1234) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1001 ( .A(
        div_DP_OP_279J39_124_314_n1240), .B(div_DP_OP_279J39_124_314_n1251), 
        .CI(div_DP_OP_279J39_124_314_n1249), .CO(
        div_DP_OP_279J39_124_314_n1231), .S(div_DP_OP_279J39_124_314_n1232) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U1000 ( .A(
        div_DP_OP_279J39_124_314_n1236), .B(div_DP_OP_279J39_124_314_n1234), 
        .CI(div_DP_OP_279J39_124_314_n1247), .CO(
        div_DP_OP_279J39_124_314_n1229), .S(div_DP_OP_279J39_124_314_n1230) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U999 ( .A(div_DP_OP_279J39_124_314_n1232), .B(div_DP_OP_279J39_124_314_n1245), .CI(div_DP_OP_279J39_124_314_n1230), 
        .CO(div_DP_OP_279J39_124_314_n1227), .S(div_DP_OP_279J39_124_314_n1228) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U998 ( .A(div_n_T_51_95_), .B(
        div_DP_OP_279J39_124_314_n1693), .CI(div_DP_OP_279J39_124_314_n2205), 
        .CO(div_DP_OP_279J39_124_314_n1225), .S(div_DP_OP_279J39_124_314_n1226) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U997 ( .A(div_DP_OP_279J39_124_314_n2141), .B(div_DP_OP_279J39_124_314_n1757), .CI(div_DP_OP_279J39_124_314_n1821), 
        .CO(div_DP_OP_279J39_124_314_n1223), .S(div_DP_OP_279J39_124_314_n1224) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U996 ( .A(div_DP_OP_279J39_124_314_n2077), .B(div_DP_OP_279J39_124_314_n1885), .CI(div_DP_OP_279J39_124_314_n1949), 
        .CO(div_DP_OP_279J39_124_314_n1221), .S(div_DP_OP_279J39_124_314_n1222) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U995 ( .A(div_DP_OP_279J39_124_314_n2013), .B(div_DP_OP_279J39_124_314_n1241), .CI(div_DP_OP_279J39_124_314_n1239), 
        .CO(div_DP_OP_279J39_124_314_n1219), .S(div_DP_OP_279J39_124_314_n1220) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U994 ( .A(div_DP_OP_279J39_124_314_n1237), .B(div_DP_OP_279J39_124_314_n1226), .CI(div_DP_OP_279J39_124_314_n1222), 
        .CO(div_DP_OP_279J39_124_314_n1217), .S(div_DP_OP_279J39_124_314_n1218) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U993 ( .A(div_DP_OP_279J39_124_314_n1224), .B(div_DP_OP_279J39_124_314_n1235), .CI(div_DP_OP_279J39_124_314_n1233), 
        .CO(div_DP_OP_279J39_124_314_n1215), .S(div_DP_OP_279J39_124_314_n1216) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U992 ( .A(div_DP_OP_279J39_124_314_n1220), .B(div_DP_OP_279J39_124_314_n1218), .CI(div_DP_OP_279J39_124_314_n1231), 
        .CO(div_DP_OP_279J39_124_314_n1213), .S(div_DP_OP_279J39_124_314_n1214) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U991 ( .A(div_DP_OP_279J39_124_314_n1216), .B(div_DP_OP_279J39_124_314_n1229), .CI(div_DP_OP_279J39_124_314_n1214), 
        .CO(div_DP_OP_279J39_124_314_n1211), .S(div_DP_OP_279J39_124_314_n1212) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U990 ( .A(div_n_T_51_96_), .B(
        div_DP_OP_279J39_124_314_n1692), .CI(div_DP_OP_279J39_124_314_n2204), 
        .CO(div_DP_OP_279J39_124_314_n1209), .S(div_DP_OP_279J39_124_314_n1210) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U989 ( .A(div_DP_OP_279J39_124_314_n2140), .B(div_DP_OP_279J39_124_314_n1756), .CI(div_DP_OP_279J39_124_314_n1820), 
        .CO(div_DP_OP_279J39_124_314_n1207), .S(div_DP_OP_279J39_124_314_n1208) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U988 ( .A(div_DP_OP_279J39_124_314_n2076), .B(div_DP_OP_279J39_124_314_n1884), .CI(div_DP_OP_279J39_124_314_n1948), 
        .CO(div_DP_OP_279J39_124_314_n1205), .S(div_DP_OP_279J39_124_314_n1206) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U987 ( .A(div_DP_OP_279J39_124_314_n2012), .B(div_DP_OP_279J39_124_314_n1225), .CI(div_DP_OP_279J39_124_314_n1223), 
        .CO(div_DP_OP_279J39_124_314_n1203), .S(div_DP_OP_279J39_124_314_n1204) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U986 ( .A(div_DP_OP_279J39_124_314_n1221), .B(div_DP_OP_279J39_124_314_n1210), .CI(div_DP_OP_279J39_124_314_n1206), 
        .CO(div_DP_OP_279J39_124_314_n1201), .S(div_DP_OP_279J39_124_314_n1202) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U985 ( .A(div_DP_OP_279J39_124_314_n1208), .B(div_DP_OP_279J39_124_314_n1219), .CI(div_DP_OP_279J39_124_314_n1217), 
        .CO(div_DP_OP_279J39_124_314_n1199), .S(div_DP_OP_279J39_124_314_n1200) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U984 ( .A(div_DP_OP_279J39_124_314_n1204), .B(div_DP_OP_279J39_124_314_n1202), .CI(div_DP_OP_279J39_124_314_n1215), 
        .CO(div_DP_OP_279J39_124_314_n1197), .S(div_DP_OP_279J39_124_314_n1198) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U983 ( .A(div_DP_OP_279J39_124_314_n1200), .B(div_DP_OP_279J39_124_314_n1213), .CI(div_DP_OP_279J39_124_314_n1198), 
        .CO(div_DP_OP_279J39_124_314_n1195), .S(div_DP_OP_279J39_124_314_n1196) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U982 ( .A(div_n_T_51_97_), .B(
        div_DP_OP_279J39_124_314_n1691), .CI(div_DP_OP_279J39_124_314_n2203), 
        .CO(div_DP_OP_279J39_124_314_n1193), .S(div_DP_OP_279J39_124_314_n1194) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U981 ( .A(div_DP_OP_279J39_124_314_n2139), .B(div_DP_OP_279J39_124_314_n1755), .CI(div_DP_OP_279J39_124_314_n1819), 
        .CO(div_DP_OP_279J39_124_314_n1191), .S(div_DP_OP_279J39_124_314_n1192) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U980 ( .A(div_DP_OP_279J39_124_314_n2075), .B(div_DP_OP_279J39_124_314_n1883), .CI(div_DP_OP_279J39_124_314_n1947), 
        .CO(div_DP_OP_279J39_124_314_n1189), .S(div_DP_OP_279J39_124_314_n1190) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U979 ( .A(div_DP_OP_279J39_124_314_n2011), .B(div_DP_OP_279J39_124_314_n1209), .CI(div_DP_OP_279J39_124_314_n1207), 
        .CO(div_DP_OP_279J39_124_314_n1187), .S(div_DP_OP_279J39_124_314_n1188) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U978 ( .A(div_DP_OP_279J39_124_314_n1205), .B(div_DP_OP_279J39_124_314_n1194), .CI(div_DP_OP_279J39_124_314_n1190), 
        .CO(div_DP_OP_279J39_124_314_n1185), .S(div_DP_OP_279J39_124_314_n1186) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U977 ( .A(div_DP_OP_279J39_124_314_n1192), .B(div_DP_OP_279J39_124_314_n1203), .CI(div_DP_OP_279J39_124_314_n1201), 
        .CO(div_DP_OP_279J39_124_314_n1183), .S(div_DP_OP_279J39_124_314_n1184) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U976 ( .A(div_DP_OP_279J39_124_314_n1188), .B(div_DP_OP_279J39_124_314_n1186), .CI(div_DP_OP_279J39_124_314_n1199), 
        .CO(div_DP_OP_279J39_124_314_n1181), .S(div_DP_OP_279J39_124_314_n1182) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U975 ( .A(div_DP_OP_279J39_124_314_n1184), .B(div_DP_OP_279J39_124_314_n1197), .CI(div_DP_OP_279J39_124_314_n1182), 
        .CO(div_DP_OP_279J39_124_314_n1179), .S(div_DP_OP_279J39_124_314_n1180) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U974 ( .A(div_n_T_51_98_), .B(
        div_DP_OP_279J39_124_314_n1690), .CI(div_DP_OP_279J39_124_314_n2202), 
        .CO(div_DP_OP_279J39_124_314_n1177), .S(div_DP_OP_279J39_124_314_n1178) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U973 ( .A(div_DP_OP_279J39_124_314_n2138), .B(div_DP_OP_279J39_124_314_n1754), .CI(div_DP_OP_279J39_124_314_n1818), 
        .CO(div_DP_OP_279J39_124_314_n1175), .S(div_DP_OP_279J39_124_314_n1176) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U972 ( .A(div_DP_OP_279J39_124_314_n2074), .B(div_DP_OP_279J39_124_314_n1882), .CI(div_DP_OP_279J39_124_314_n1946), 
        .CO(div_DP_OP_279J39_124_314_n1173), .S(div_DP_OP_279J39_124_314_n1174) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U971 ( .A(div_DP_OP_279J39_124_314_n2010), .B(div_DP_OP_279J39_124_314_n1193), .CI(div_DP_OP_279J39_124_314_n1191), 
        .CO(div_DP_OP_279J39_124_314_n1171), .S(div_DP_OP_279J39_124_314_n1172) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U970 ( .A(div_DP_OP_279J39_124_314_n1189), .B(div_DP_OP_279J39_124_314_n1178), .CI(div_DP_OP_279J39_124_314_n1174), 
        .CO(div_DP_OP_279J39_124_314_n1169), .S(div_DP_OP_279J39_124_314_n1170) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U969 ( .A(div_DP_OP_279J39_124_314_n1176), .B(div_DP_OP_279J39_124_314_n1187), .CI(div_DP_OP_279J39_124_314_n1185), 
        .CO(div_DP_OP_279J39_124_314_n1167), .S(div_DP_OP_279J39_124_314_n1168) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U968 ( .A(div_DP_OP_279J39_124_314_n1172), .B(div_DP_OP_279J39_124_314_n1170), .CI(div_DP_OP_279J39_124_314_n1183), 
        .CO(div_DP_OP_279J39_124_314_n1165), .S(div_DP_OP_279J39_124_314_n1166) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U967 ( .A(div_DP_OP_279J39_124_314_n1168), .B(div_DP_OP_279J39_124_314_n1181), .CI(div_DP_OP_279J39_124_314_n1166), 
        .CO(div_DP_OP_279J39_124_314_n1163), .S(div_DP_OP_279J39_124_314_n1164) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U966 ( .A(div_n_T_51_99_), .B(
        div_DP_OP_279J39_124_314_n1689), .CI(div_DP_OP_279J39_124_314_n2201), 
        .CO(div_DP_OP_279J39_124_314_n1161), .S(div_DP_OP_279J39_124_314_n1162) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U965 ( .A(div_DP_OP_279J39_124_314_n2137), .B(div_DP_OP_279J39_124_314_n1753), .CI(div_DP_OP_279J39_124_314_n1817), 
        .CO(div_DP_OP_279J39_124_314_n1159), .S(div_DP_OP_279J39_124_314_n1160) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U964 ( .A(div_DP_OP_279J39_124_314_n2073), .B(div_DP_OP_279J39_124_314_n1881), .CI(div_DP_OP_279J39_124_314_n1945), 
        .CO(div_DP_OP_279J39_124_314_n1157), .S(div_DP_OP_279J39_124_314_n1158) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U963 ( .A(div_DP_OP_279J39_124_314_n2009), .B(div_DP_OP_279J39_124_314_n1177), .CI(div_DP_OP_279J39_124_314_n1175), 
        .CO(div_DP_OP_279J39_124_314_n1155), .S(div_DP_OP_279J39_124_314_n1156) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U962 ( .A(div_DP_OP_279J39_124_314_n1173), .B(div_DP_OP_279J39_124_314_n1162), .CI(div_DP_OP_279J39_124_314_n1158), 
        .CO(div_DP_OP_279J39_124_314_n1153), .S(div_DP_OP_279J39_124_314_n1154) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U961 ( .A(div_DP_OP_279J39_124_314_n1160), .B(div_DP_OP_279J39_124_314_n1171), .CI(div_DP_OP_279J39_124_314_n1169), 
        .CO(div_DP_OP_279J39_124_314_n1151), .S(div_DP_OP_279J39_124_314_n1152) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U960 ( .A(div_DP_OP_279J39_124_314_n1156), .B(div_DP_OP_279J39_124_314_n1154), .CI(div_DP_OP_279J39_124_314_n1167), 
        .CO(div_DP_OP_279J39_124_314_n1149), .S(div_DP_OP_279J39_124_314_n1150) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U959 ( .A(div_DP_OP_279J39_124_314_n1152), .B(div_DP_OP_279J39_124_314_n1165), .CI(div_DP_OP_279J39_124_314_n1150), 
        .CO(div_DP_OP_279J39_124_314_n1147), .S(div_DP_OP_279J39_124_314_n1148) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U958 ( .A(div_n_T_51_100_), .B(
        div_DP_OP_279J39_124_314_n1688), .CI(div_DP_OP_279J39_124_314_n2200), 
        .CO(div_DP_OP_279J39_124_314_n1145), .S(div_DP_OP_279J39_124_314_n1146) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U957 ( .A(div_DP_OP_279J39_124_314_n2136), .B(div_DP_OP_279J39_124_314_n1752), .CI(div_DP_OP_279J39_124_314_n1816), 
        .CO(div_DP_OP_279J39_124_314_n1143), .S(div_DP_OP_279J39_124_314_n1144) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U956 ( .A(div_DP_OP_279J39_124_314_n2072), .B(div_DP_OP_279J39_124_314_n1880), .CI(div_DP_OP_279J39_124_314_n1944), 
        .CO(div_DP_OP_279J39_124_314_n1141), .S(div_DP_OP_279J39_124_314_n1142) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U955 ( .A(div_DP_OP_279J39_124_314_n2008), .B(div_DP_OP_279J39_124_314_n1161), .CI(div_DP_OP_279J39_124_314_n1159), 
        .CO(div_DP_OP_279J39_124_314_n1139), .S(div_DP_OP_279J39_124_314_n1140) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U954 ( .A(div_DP_OP_279J39_124_314_n1157), .B(div_DP_OP_279J39_124_314_n1146), .CI(div_DP_OP_279J39_124_314_n1142), 
        .CO(div_DP_OP_279J39_124_314_n1137), .S(div_DP_OP_279J39_124_314_n1138) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U953 ( .A(div_DP_OP_279J39_124_314_n1144), .B(div_DP_OP_279J39_124_314_n1155), .CI(div_DP_OP_279J39_124_314_n1153), 
        .CO(div_DP_OP_279J39_124_314_n1135), .S(div_DP_OP_279J39_124_314_n1136) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U952 ( .A(div_DP_OP_279J39_124_314_n1140), .B(div_DP_OP_279J39_124_314_n1138), .CI(div_DP_OP_279J39_124_314_n1151), 
        .CO(div_DP_OP_279J39_124_314_n1133), .S(div_DP_OP_279J39_124_314_n1134) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U951 ( .A(div_DP_OP_279J39_124_314_n1136), .B(div_DP_OP_279J39_124_314_n1149), .CI(div_DP_OP_279J39_124_314_n1134), 
        .CO(div_DP_OP_279J39_124_314_n1131), .S(div_DP_OP_279J39_124_314_n1132) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U950 ( .A(div_n_T_51_101_), .B(
        div_DP_OP_279J39_124_314_n1687), .CI(div_DP_OP_279J39_124_314_n2199), 
        .CO(div_DP_OP_279J39_124_314_n1129), .S(div_DP_OP_279J39_124_314_n1130) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U949 ( .A(div_DP_OP_279J39_124_314_n2135), .B(div_DP_OP_279J39_124_314_n1751), .CI(div_DP_OP_279J39_124_314_n1815), 
        .CO(div_DP_OP_279J39_124_314_n1127), .S(div_DP_OP_279J39_124_314_n1128) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U948 ( .A(div_DP_OP_279J39_124_314_n2071), .B(div_DP_OP_279J39_124_314_n1879), .CI(div_DP_OP_279J39_124_314_n1943), 
        .CO(div_DP_OP_279J39_124_314_n1125), .S(div_DP_OP_279J39_124_314_n1126) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U947 ( .A(div_DP_OP_279J39_124_314_n2007), .B(div_DP_OP_279J39_124_314_n1145), .CI(div_DP_OP_279J39_124_314_n1143), 
        .CO(div_DP_OP_279J39_124_314_n1123), .S(div_DP_OP_279J39_124_314_n1124) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U946 ( .A(div_DP_OP_279J39_124_314_n1141), .B(div_DP_OP_279J39_124_314_n1130), .CI(div_DP_OP_279J39_124_314_n1126), 
        .CO(div_DP_OP_279J39_124_314_n1121), .S(div_DP_OP_279J39_124_314_n1122) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U945 ( .A(div_DP_OP_279J39_124_314_n1128), .B(div_DP_OP_279J39_124_314_n1139), .CI(div_DP_OP_279J39_124_314_n1137), 
        .CO(div_DP_OP_279J39_124_314_n1119), .S(div_DP_OP_279J39_124_314_n1120) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U944 ( .A(div_DP_OP_279J39_124_314_n1124), .B(div_DP_OP_279J39_124_314_n1122), .CI(div_DP_OP_279J39_124_314_n1135), 
        .CO(div_DP_OP_279J39_124_314_n1117), .S(div_DP_OP_279J39_124_314_n1118) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U943 ( .A(div_DP_OP_279J39_124_314_n1120), .B(div_DP_OP_279J39_124_314_n1133), .CI(div_DP_OP_279J39_124_314_n1118), 
        .CO(div_DP_OP_279J39_124_314_n1115), .S(div_DP_OP_279J39_124_314_n1116) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U942 ( .A(div_n_T_51_102_), .B(
        div_DP_OP_279J39_124_314_n1686), .CI(div_DP_OP_279J39_124_314_n2198), 
        .CO(div_DP_OP_279J39_124_314_n1113), .S(div_DP_OP_279J39_124_314_n1114) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U941 ( .A(div_DP_OP_279J39_124_314_n2134), .B(div_DP_OP_279J39_124_314_n1750), .CI(div_DP_OP_279J39_124_314_n1814), 
        .CO(div_DP_OP_279J39_124_314_n1111), .S(div_DP_OP_279J39_124_314_n1112) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U940 ( .A(div_DP_OP_279J39_124_314_n2070), .B(div_DP_OP_279J39_124_314_n1878), .CI(div_DP_OP_279J39_124_314_n1942), 
        .CO(div_DP_OP_279J39_124_314_n1109), .S(div_DP_OP_279J39_124_314_n1110) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U939 ( .A(div_DP_OP_279J39_124_314_n2006), .B(div_DP_OP_279J39_124_314_n1129), .CI(div_DP_OP_279J39_124_314_n1127), 
        .CO(div_DP_OP_279J39_124_314_n1107), .S(div_DP_OP_279J39_124_314_n1108) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U938 ( .A(div_DP_OP_279J39_124_314_n1125), .B(div_DP_OP_279J39_124_314_n1114), .CI(div_DP_OP_279J39_124_314_n1110), 
        .CO(div_DP_OP_279J39_124_314_n1105), .S(div_DP_OP_279J39_124_314_n1106) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U937 ( .A(div_DP_OP_279J39_124_314_n1112), .B(div_DP_OP_279J39_124_314_n1123), .CI(div_DP_OP_279J39_124_314_n1121), 
        .CO(div_DP_OP_279J39_124_314_n1103), .S(div_DP_OP_279J39_124_314_n1104) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U936 ( .A(div_DP_OP_279J39_124_314_n1108), .B(div_DP_OP_279J39_124_314_n1106), .CI(div_DP_OP_279J39_124_314_n1119), 
        .CO(div_DP_OP_279J39_124_314_n1101), .S(div_DP_OP_279J39_124_314_n1102) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U935 ( .A(div_DP_OP_279J39_124_314_n1104), .B(div_DP_OP_279J39_124_314_n1117), .CI(div_DP_OP_279J39_124_314_n1102), 
        .CO(div_DP_OP_279J39_124_314_n1099), .S(div_DP_OP_279J39_124_314_n1100) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U934 ( .A(div_n_T_51_103_), .B(
        div_DP_OP_279J39_124_314_n1685), .CI(div_DP_OP_279J39_124_314_n2197), 
        .CO(div_DP_OP_279J39_124_314_n1097), .S(div_DP_OP_279J39_124_314_n1098) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U933 ( .A(div_DP_OP_279J39_124_314_n2133), .B(div_DP_OP_279J39_124_314_n1749), .CI(div_DP_OP_279J39_124_314_n1813), 
        .CO(div_DP_OP_279J39_124_314_n1095), .S(div_DP_OP_279J39_124_314_n1096) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U932 ( .A(div_DP_OP_279J39_124_314_n2069), .B(div_DP_OP_279J39_124_314_n1877), .CI(div_DP_OP_279J39_124_314_n1941), 
        .CO(div_DP_OP_279J39_124_314_n1093), .S(div_DP_OP_279J39_124_314_n1094) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U931 ( .A(div_DP_OP_279J39_124_314_n2005), .B(div_DP_OP_279J39_124_314_n1113), .CI(div_DP_OP_279J39_124_314_n1111), 
        .CO(div_DP_OP_279J39_124_314_n1091), .S(div_DP_OP_279J39_124_314_n1092) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U930 ( .A(div_DP_OP_279J39_124_314_n1109), .B(div_DP_OP_279J39_124_314_n1098), .CI(div_DP_OP_279J39_124_314_n1094), 
        .CO(div_DP_OP_279J39_124_314_n1089), .S(div_DP_OP_279J39_124_314_n1090) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U929 ( .A(div_DP_OP_279J39_124_314_n1096), .B(div_DP_OP_279J39_124_314_n1107), .CI(div_DP_OP_279J39_124_314_n1105), 
        .CO(div_DP_OP_279J39_124_314_n1087), .S(div_DP_OP_279J39_124_314_n1088) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U928 ( .A(div_DP_OP_279J39_124_314_n1092), .B(div_DP_OP_279J39_124_314_n1090), .CI(div_DP_OP_279J39_124_314_n1103), 
        .CO(div_DP_OP_279J39_124_314_n1085), .S(div_DP_OP_279J39_124_314_n1086) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U927 ( .A(div_DP_OP_279J39_124_314_n1088), .B(div_DP_OP_279J39_124_314_n1101), .CI(div_DP_OP_279J39_124_314_n1086), 
        .CO(div_DP_OP_279J39_124_314_n1083), .S(div_DP_OP_279J39_124_314_n1084) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U926 ( .A(div_n_T_51_104_), .B(
        div_DP_OP_279J39_124_314_n1684), .CI(div_DP_OP_279J39_124_314_n2196), 
        .CO(div_DP_OP_279J39_124_314_n1081), .S(div_DP_OP_279J39_124_314_n1082) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U925 ( .A(div_DP_OP_279J39_124_314_n2132), .B(div_DP_OP_279J39_124_314_n1748), .CI(div_DP_OP_279J39_124_314_n1812), 
        .CO(div_DP_OP_279J39_124_314_n1079), .S(div_DP_OP_279J39_124_314_n1080) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U924 ( .A(div_DP_OP_279J39_124_314_n2068), .B(div_DP_OP_279J39_124_314_n1876), .CI(div_DP_OP_279J39_124_314_n1940), 
        .CO(div_DP_OP_279J39_124_314_n1077), .S(div_DP_OP_279J39_124_314_n1078) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U923 ( .A(div_DP_OP_279J39_124_314_n2004), .B(div_DP_OP_279J39_124_314_n1097), .CI(div_DP_OP_279J39_124_314_n1095), 
        .CO(div_DP_OP_279J39_124_314_n1075), .S(div_DP_OP_279J39_124_314_n1076) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U922 ( .A(div_DP_OP_279J39_124_314_n1093), .B(div_DP_OP_279J39_124_314_n1082), .CI(div_DP_OP_279J39_124_314_n1078), 
        .CO(div_DP_OP_279J39_124_314_n1073), .S(div_DP_OP_279J39_124_314_n1074) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U921 ( .A(div_DP_OP_279J39_124_314_n1080), .B(div_DP_OP_279J39_124_314_n1091), .CI(div_DP_OP_279J39_124_314_n1089), 
        .CO(div_DP_OP_279J39_124_314_n1071), .S(div_DP_OP_279J39_124_314_n1072) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U920 ( .A(div_DP_OP_279J39_124_314_n1076), .B(div_DP_OP_279J39_124_314_n1074), .CI(div_DP_OP_279J39_124_314_n1087), 
        .CO(div_DP_OP_279J39_124_314_n1069), .S(div_DP_OP_279J39_124_314_n1070) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U919 ( .A(div_DP_OP_279J39_124_314_n1072), .B(div_DP_OP_279J39_124_314_n1085), .CI(div_DP_OP_279J39_124_314_n1070), 
        .CO(div_DP_OP_279J39_124_314_n1067), .S(div_DP_OP_279J39_124_314_n1068) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U918 ( .A(div_n_T_51_105_), .B(
        div_DP_OP_279J39_124_314_n1683), .CI(div_DP_OP_279J39_124_314_n2195), 
        .CO(div_DP_OP_279J39_124_314_n1065), .S(div_DP_OP_279J39_124_314_n1066) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U917 ( .A(div_DP_OP_279J39_124_314_n2131), .B(div_DP_OP_279J39_124_314_n1747), .CI(div_DP_OP_279J39_124_314_n1811), 
        .CO(div_DP_OP_279J39_124_314_n1063), .S(div_DP_OP_279J39_124_314_n1064) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U916 ( .A(div_DP_OP_279J39_124_314_n2067), .B(div_DP_OP_279J39_124_314_n1875), .CI(div_DP_OP_279J39_124_314_n1939), 
        .CO(div_DP_OP_279J39_124_314_n1061), .S(div_DP_OP_279J39_124_314_n1062) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U915 ( .A(div_DP_OP_279J39_124_314_n2003), .B(div_DP_OP_279J39_124_314_n1081), .CI(div_DP_OP_279J39_124_314_n1079), 
        .CO(div_DP_OP_279J39_124_314_n1059), .S(div_DP_OP_279J39_124_314_n1060) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U914 ( .A(div_DP_OP_279J39_124_314_n1077), .B(div_DP_OP_279J39_124_314_n1066), .CI(div_DP_OP_279J39_124_314_n1062), 
        .CO(div_DP_OP_279J39_124_314_n1057), .S(div_DP_OP_279J39_124_314_n1058) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U913 ( .A(div_DP_OP_279J39_124_314_n1064), .B(div_DP_OP_279J39_124_314_n1075), .CI(div_DP_OP_279J39_124_314_n1073), 
        .CO(div_DP_OP_279J39_124_314_n1055), .S(div_DP_OP_279J39_124_314_n1056) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U912 ( .A(div_DP_OP_279J39_124_314_n1060), .B(div_DP_OP_279J39_124_314_n1058), .CI(div_DP_OP_279J39_124_314_n1071), 
        .CO(div_DP_OP_279J39_124_314_n1053), .S(div_DP_OP_279J39_124_314_n1054) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U911 ( .A(div_DP_OP_279J39_124_314_n1056), .B(div_DP_OP_279J39_124_314_n1069), .CI(div_DP_OP_279J39_124_314_n1054), 
        .CO(div_DP_OP_279J39_124_314_n1051), .S(div_DP_OP_279J39_124_314_n1052) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U910 ( .A(div_n_T_51_106_), .B(
        div_DP_OP_279J39_124_314_n1682), .CI(div_DP_OP_279J39_124_314_n2194), 
        .CO(div_DP_OP_279J39_124_314_n1049), .S(div_DP_OP_279J39_124_314_n1050) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U909 ( .A(div_DP_OP_279J39_124_314_n2130), .B(div_DP_OP_279J39_124_314_n1746), .CI(div_DP_OP_279J39_124_314_n1810), 
        .CO(div_DP_OP_279J39_124_314_n1047), .S(div_DP_OP_279J39_124_314_n1048) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U908 ( .A(div_DP_OP_279J39_124_314_n2066), .B(div_DP_OP_279J39_124_314_n1874), .CI(div_DP_OP_279J39_124_314_n1938), 
        .CO(div_DP_OP_279J39_124_314_n1045), .S(div_DP_OP_279J39_124_314_n1046) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U907 ( .A(div_DP_OP_279J39_124_314_n2002), .B(div_DP_OP_279J39_124_314_n1065), .CI(div_DP_OP_279J39_124_314_n1063), 
        .CO(div_DP_OP_279J39_124_314_n1043), .S(div_DP_OP_279J39_124_314_n1044) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U906 ( .A(div_DP_OP_279J39_124_314_n1061), .B(div_DP_OP_279J39_124_314_n1050), .CI(div_DP_OP_279J39_124_314_n1046), 
        .CO(div_DP_OP_279J39_124_314_n1041), .S(div_DP_OP_279J39_124_314_n1042) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U905 ( .A(div_DP_OP_279J39_124_314_n1048), .B(div_DP_OP_279J39_124_314_n1059), .CI(div_DP_OP_279J39_124_314_n1057), 
        .CO(div_DP_OP_279J39_124_314_n1039), .S(div_DP_OP_279J39_124_314_n1040) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U904 ( .A(div_DP_OP_279J39_124_314_n1044), .B(div_DP_OP_279J39_124_314_n1042), .CI(div_DP_OP_279J39_124_314_n1055), 
        .CO(div_DP_OP_279J39_124_314_n1037), .S(div_DP_OP_279J39_124_314_n1038) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U903 ( .A(div_DP_OP_279J39_124_314_n1040), .B(div_DP_OP_279J39_124_314_n1053), .CI(div_DP_OP_279J39_124_314_n1038), 
        .CO(div_DP_OP_279J39_124_314_n1035), .S(div_DP_OP_279J39_124_314_n1036) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U902 ( .A(div_n_T_51_107_), .B(
        div_DP_OP_279J39_124_314_n1681), .CI(div_DP_OP_279J39_124_314_n2193), 
        .CO(div_DP_OP_279J39_124_314_n1033), .S(div_DP_OP_279J39_124_314_n1034) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U901 ( .A(div_DP_OP_279J39_124_314_n2129), .B(div_DP_OP_279J39_124_314_n1745), .CI(div_DP_OP_279J39_124_314_n1809), 
        .CO(div_DP_OP_279J39_124_314_n1031), .S(div_DP_OP_279J39_124_314_n1032) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U900 ( .A(div_DP_OP_279J39_124_314_n2065), .B(div_DP_OP_279J39_124_314_n1873), .CI(div_DP_OP_279J39_124_314_n1937), 
        .CO(div_DP_OP_279J39_124_314_n1029), .S(div_DP_OP_279J39_124_314_n1030) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U899 ( .A(div_DP_OP_279J39_124_314_n2001), .B(div_DP_OP_279J39_124_314_n1049), .CI(div_DP_OP_279J39_124_314_n1047), 
        .CO(div_DP_OP_279J39_124_314_n1027), .S(div_DP_OP_279J39_124_314_n1028) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U898 ( .A(div_DP_OP_279J39_124_314_n1045), .B(div_DP_OP_279J39_124_314_n1034), .CI(div_DP_OP_279J39_124_314_n1030), 
        .CO(div_DP_OP_279J39_124_314_n1025), .S(div_DP_OP_279J39_124_314_n1026) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U897 ( .A(div_DP_OP_279J39_124_314_n1032), .B(div_DP_OP_279J39_124_314_n1043), .CI(div_DP_OP_279J39_124_314_n1041), 
        .CO(div_DP_OP_279J39_124_314_n1023), .S(div_DP_OP_279J39_124_314_n1024) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U896 ( .A(div_DP_OP_279J39_124_314_n1028), .B(div_DP_OP_279J39_124_314_n1026), .CI(div_DP_OP_279J39_124_314_n1039), 
        .CO(div_DP_OP_279J39_124_314_n1021), .S(div_DP_OP_279J39_124_314_n1022) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U895 ( .A(div_DP_OP_279J39_124_314_n1024), .B(div_DP_OP_279J39_124_314_n1037), .CI(div_DP_OP_279J39_124_314_n1022), 
        .CO(div_DP_OP_279J39_124_314_n1019), .S(div_DP_OP_279J39_124_314_n1020) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U894 ( .A(div_n_T_51_108_), .B(
        div_DP_OP_279J39_124_314_n1680), .CI(div_DP_OP_279J39_124_314_n2192), 
        .CO(div_DP_OP_279J39_124_314_n1017), .S(div_DP_OP_279J39_124_314_n1018) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U893 ( .A(div_DP_OP_279J39_124_314_n2128), .B(div_DP_OP_279J39_124_314_n1744), .CI(div_DP_OP_279J39_124_314_n1808), 
        .CO(div_DP_OP_279J39_124_314_n1015), .S(div_DP_OP_279J39_124_314_n1016) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U892 ( .A(div_DP_OP_279J39_124_314_n2064), .B(div_DP_OP_279J39_124_314_n1872), .CI(div_DP_OP_279J39_124_314_n1936), 
        .CO(div_DP_OP_279J39_124_314_n1013), .S(div_DP_OP_279J39_124_314_n1014) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U891 ( .A(div_DP_OP_279J39_124_314_n2000), .B(div_DP_OP_279J39_124_314_n1033), .CI(div_DP_OP_279J39_124_314_n1031), 
        .CO(div_DP_OP_279J39_124_314_n1011), .S(div_DP_OP_279J39_124_314_n1012) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U890 ( .A(div_DP_OP_279J39_124_314_n1029), .B(div_DP_OP_279J39_124_314_n1018), .CI(div_DP_OP_279J39_124_314_n1014), 
        .CO(div_DP_OP_279J39_124_314_n1009), .S(div_DP_OP_279J39_124_314_n1010) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U889 ( .A(div_DP_OP_279J39_124_314_n1016), .B(div_DP_OP_279J39_124_314_n1027), .CI(div_DP_OP_279J39_124_314_n1025), 
        .CO(div_DP_OP_279J39_124_314_n1007), .S(div_DP_OP_279J39_124_314_n1008) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U888 ( .A(div_DP_OP_279J39_124_314_n1012), .B(div_DP_OP_279J39_124_314_n1010), .CI(div_DP_OP_279J39_124_314_n1023), 
        .CO(div_DP_OP_279J39_124_314_n1005), .S(div_DP_OP_279J39_124_314_n1006) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U887 ( .A(div_DP_OP_279J39_124_314_n1008), .B(div_DP_OP_279J39_124_314_n1021), .CI(div_DP_OP_279J39_124_314_n1006), 
        .CO(div_DP_OP_279J39_124_314_n1003), .S(div_DP_OP_279J39_124_314_n1004) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U886 ( .A(div_n_T_51_109_), .B(
        div_DP_OP_279J39_124_314_n1679), .CI(div_DP_OP_279J39_124_314_n2191), 
        .CO(div_DP_OP_279J39_124_314_n1001), .S(div_DP_OP_279J39_124_314_n1002) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U885 ( .A(div_DP_OP_279J39_124_314_n2127), .B(div_DP_OP_279J39_124_314_n1743), .CI(div_DP_OP_279J39_124_314_n1807), 
        .CO(div_DP_OP_279J39_124_314_n999), .S(div_DP_OP_279J39_124_314_n1000)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U884 ( .A(div_DP_OP_279J39_124_314_n2063), .B(div_DP_OP_279J39_124_314_n1871), .CI(div_DP_OP_279J39_124_314_n1935), 
        .CO(div_DP_OP_279J39_124_314_n997), .S(div_DP_OP_279J39_124_314_n998)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U883 ( .A(div_DP_OP_279J39_124_314_n1999), .B(div_DP_OP_279J39_124_314_n1017), .CI(div_DP_OP_279J39_124_314_n1015), 
        .CO(div_DP_OP_279J39_124_314_n995), .S(div_DP_OP_279J39_124_314_n996)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U882 ( .A(div_DP_OP_279J39_124_314_n1013), .B(div_DP_OP_279J39_124_314_n1002), .CI(div_DP_OP_279J39_124_314_n998), .CO(
        div_DP_OP_279J39_124_314_n993), .S(div_DP_OP_279J39_124_314_n994) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U881 ( .A(div_DP_OP_279J39_124_314_n1000), .B(div_DP_OP_279J39_124_314_n1011), .CI(div_DP_OP_279J39_124_314_n1009), 
        .CO(div_DP_OP_279J39_124_314_n991), .S(div_DP_OP_279J39_124_314_n992)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U880 ( .A(div_DP_OP_279J39_124_314_n996), 
        .B(div_DP_OP_279J39_124_314_n994), .CI(div_DP_OP_279J39_124_314_n1007), 
        .CO(div_DP_OP_279J39_124_314_n989), .S(div_DP_OP_279J39_124_314_n990)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U879 ( .A(div_DP_OP_279J39_124_314_n992), 
        .B(div_DP_OP_279J39_124_314_n1005), .CI(div_DP_OP_279J39_124_314_n990), 
        .CO(div_DP_OP_279J39_124_314_n987), .S(div_DP_OP_279J39_124_314_n988)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U878 ( .A(div_n_T_51_110_), .B(
        div_DP_OP_279J39_124_314_n1678), .CI(div_DP_OP_279J39_124_314_n2190), 
        .CO(div_DP_OP_279J39_124_314_n985), .S(div_DP_OP_279J39_124_314_n986)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U877 ( .A(div_DP_OP_279J39_124_314_n2126), .B(div_DP_OP_279J39_124_314_n1742), .CI(div_DP_OP_279J39_124_314_n1806), 
        .CO(div_DP_OP_279J39_124_314_n983), .S(div_DP_OP_279J39_124_314_n984)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U876 ( .A(div_DP_OP_279J39_124_314_n2062), .B(div_DP_OP_279J39_124_314_n1870), .CI(div_DP_OP_279J39_124_314_n1934), 
        .CO(div_DP_OP_279J39_124_314_n981), .S(div_DP_OP_279J39_124_314_n982)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U875 ( .A(div_DP_OP_279J39_124_314_n1998), .B(div_DP_OP_279J39_124_314_n1001), .CI(div_DP_OP_279J39_124_314_n999), .CO(
        div_DP_OP_279J39_124_314_n979), .S(div_DP_OP_279J39_124_314_n980) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U874 ( .A(div_DP_OP_279J39_124_314_n997), 
        .B(div_DP_OP_279J39_124_314_n986), .CI(div_DP_OP_279J39_124_314_n982), 
        .CO(div_DP_OP_279J39_124_314_n977), .S(div_DP_OP_279J39_124_314_n978)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U873 ( .A(div_DP_OP_279J39_124_314_n984), 
        .B(div_DP_OP_279J39_124_314_n995), .CI(div_DP_OP_279J39_124_314_n993), 
        .CO(div_DP_OP_279J39_124_314_n975), .S(div_DP_OP_279J39_124_314_n976)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U872 ( .A(div_DP_OP_279J39_124_314_n980), 
        .B(div_DP_OP_279J39_124_314_n978), .CI(div_DP_OP_279J39_124_314_n991), 
        .CO(div_DP_OP_279J39_124_314_n973), .S(div_DP_OP_279J39_124_314_n974)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U871 ( .A(div_DP_OP_279J39_124_314_n976), 
        .B(div_DP_OP_279J39_124_314_n989), .CI(div_DP_OP_279J39_124_314_n974), 
        .CO(div_DP_OP_279J39_124_314_n971), .S(div_DP_OP_279J39_124_314_n972)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U870 ( .A(div_n_T_51_111_), .B(
        div_DP_OP_279J39_124_314_n1677), .CI(div_DP_OP_279J39_124_314_n2189), 
        .CO(div_DP_OP_279J39_124_314_n969), .S(div_DP_OP_279J39_124_314_n970)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U869 ( .A(div_DP_OP_279J39_124_314_n2125), .B(div_DP_OP_279J39_124_314_n1741), .CI(div_DP_OP_279J39_124_314_n1805), 
        .CO(div_DP_OP_279J39_124_314_n967), .S(div_DP_OP_279J39_124_314_n968)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U868 ( .A(div_DP_OP_279J39_124_314_n2061), .B(div_DP_OP_279J39_124_314_n1869), .CI(div_DP_OP_279J39_124_314_n1933), 
        .CO(div_DP_OP_279J39_124_314_n965), .S(div_DP_OP_279J39_124_314_n966)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U867 ( .A(div_DP_OP_279J39_124_314_n1997), .B(div_DP_OP_279J39_124_314_n985), .CI(div_DP_OP_279J39_124_314_n983), .CO(
        div_DP_OP_279J39_124_314_n963), .S(div_DP_OP_279J39_124_314_n964) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U866 ( .A(div_DP_OP_279J39_124_314_n981), 
        .B(div_DP_OP_279J39_124_314_n970), .CI(div_DP_OP_279J39_124_314_n966), 
        .CO(div_DP_OP_279J39_124_314_n961), .S(div_DP_OP_279J39_124_314_n962)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U865 ( .A(div_DP_OP_279J39_124_314_n968), 
        .B(div_DP_OP_279J39_124_314_n979), .CI(div_DP_OP_279J39_124_314_n977), 
        .CO(div_DP_OP_279J39_124_314_n959), .S(div_DP_OP_279J39_124_314_n960)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U864 ( .A(div_DP_OP_279J39_124_314_n964), 
        .B(div_DP_OP_279J39_124_314_n962), .CI(div_DP_OP_279J39_124_314_n975), 
        .CO(div_DP_OP_279J39_124_314_n957), .S(div_DP_OP_279J39_124_314_n958)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U863 ( .A(div_DP_OP_279J39_124_314_n960), 
        .B(div_DP_OP_279J39_124_314_n973), .CI(div_DP_OP_279J39_124_314_n958), 
        .CO(div_DP_OP_279J39_124_314_n955), .S(div_DP_OP_279J39_124_314_n956)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U862 ( .A(div_n_T_51_112_), .B(
        div_DP_OP_279J39_124_314_n1676), .CI(div_DP_OP_279J39_124_314_n2188), 
        .CO(div_DP_OP_279J39_124_314_n953), .S(div_DP_OP_279J39_124_314_n954)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U861 ( .A(div_DP_OP_279J39_124_314_n2124), .B(div_DP_OP_279J39_124_314_n1740), .CI(div_DP_OP_279J39_124_314_n1804), 
        .CO(div_DP_OP_279J39_124_314_n951), .S(div_DP_OP_279J39_124_314_n952)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U860 ( .A(div_DP_OP_279J39_124_314_n2060), .B(div_DP_OP_279J39_124_314_n1868), .CI(div_DP_OP_279J39_124_314_n1932), 
        .CO(div_DP_OP_279J39_124_314_n949), .S(div_DP_OP_279J39_124_314_n950)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U859 ( .A(div_DP_OP_279J39_124_314_n1996), .B(div_DP_OP_279J39_124_314_n969), .CI(div_DP_OP_279J39_124_314_n967), .CO(
        div_DP_OP_279J39_124_314_n947), .S(div_DP_OP_279J39_124_314_n948) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U858 ( .A(div_DP_OP_279J39_124_314_n965), 
        .B(div_DP_OP_279J39_124_314_n954), .CI(div_DP_OP_279J39_124_314_n950), 
        .CO(div_DP_OP_279J39_124_314_n945), .S(div_DP_OP_279J39_124_314_n946)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U857 ( .A(div_DP_OP_279J39_124_314_n952), 
        .B(div_DP_OP_279J39_124_314_n963), .CI(div_DP_OP_279J39_124_314_n961), 
        .CO(div_DP_OP_279J39_124_314_n943), .S(div_DP_OP_279J39_124_314_n944)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U856 ( .A(div_DP_OP_279J39_124_314_n948), 
        .B(div_DP_OP_279J39_124_314_n946), .CI(div_DP_OP_279J39_124_314_n959), 
        .CO(div_DP_OP_279J39_124_314_n941), .S(div_DP_OP_279J39_124_314_n942)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U855 ( .A(div_DP_OP_279J39_124_314_n944), 
        .B(div_DP_OP_279J39_124_314_n957), .CI(div_DP_OP_279J39_124_314_n942), 
        .CO(div_DP_OP_279J39_124_314_n939), .S(div_DP_OP_279J39_124_314_n940)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U854 ( .A(div_n_T_51_113_), .B(
        div_DP_OP_279J39_124_314_n1675), .CI(div_DP_OP_279J39_124_314_n2187), 
        .CO(div_DP_OP_279J39_124_314_n937), .S(div_DP_OP_279J39_124_314_n938)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U853 ( .A(div_DP_OP_279J39_124_314_n2123), .B(div_DP_OP_279J39_124_314_n1739), .CI(div_DP_OP_279J39_124_314_n1803), 
        .CO(div_DP_OP_279J39_124_314_n935), .S(div_DP_OP_279J39_124_314_n936)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U852 ( .A(div_DP_OP_279J39_124_314_n2059), .B(div_DP_OP_279J39_124_314_n1867), .CI(div_DP_OP_279J39_124_314_n1931), 
        .CO(div_DP_OP_279J39_124_314_n933), .S(div_DP_OP_279J39_124_314_n934)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U851 ( .A(div_DP_OP_279J39_124_314_n1995), .B(div_DP_OP_279J39_124_314_n953), .CI(div_DP_OP_279J39_124_314_n951), .CO(
        div_DP_OP_279J39_124_314_n931), .S(div_DP_OP_279J39_124_314_n932) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U850 ( .A(div_DP_OP_279J39_124_314_n949), 
        .B(div_DP_OP_279J39_124_314_n938), .CI(div_DP_OP_279J39_124_314_n934), 
        .CO(div_DP_OP_279J39_124_314_n929), .S(div_DP_OP_279J39_124_314_n930)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U849 ( .A(div_DP_OP_279J39_124_314_n936), 
        .B(div_DP_OP_279J39_124_314_n947), .CI(div_DP_OP_279J39_124_314_n945), 
        .CO(div_DP_OP_279J39_124_314_n927), .S(div_DP_OP_279J39_124_314_n928)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U848 ( .A(div_DP_OP_279J39_124_314_n932), 
        .B(div_DP_OP_279J39_124_314_n930), .CI(div_DP_OP_279J39_124_314_n943), 
        .CO(div_DP_OP_279J39_124_314_n925), .S(div_DP_OP_279J39_124_314_n926)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U847 ( .A(div_DP_OP_279J39_124_314_n928), 
        .B(div_DP_OP_279J39_124_314_n941), .CI(div_DP_OP_279J39_124_314_n926), 
        .CO(div_DP_OP_279J39_124_314_n923), .S(div_DP_OP_279J39_124_314_n924)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U846 ( .A(div_n_T_51_114_), .B(
        div_DP_OP_279J39_124_314_n1674), .CI(div_DP_OP_279J39_124_314_n2186), 
        .CO(div_DP_OP_279J39_124_314_n921), .S(div_DP_OP_279J39_124_314_n922)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U845 ( .A(div_DP_OP_279J39_124_314_n2122), .B(div_DP_OP_279J39_124_314_n1738), .CI(div_DP_OP_279J39_124_314_n1802), 
        .CO(div_DP_OP_279J39_124_314_n919), .S(div_DP_OP_279J39_124_314_n920)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U844 ( .A(div_DP_OP_279J39_124_314_n2058), .B(div_DP_OP_279J39_124_314_n1866), .CI(div_DP_OP_279J39_124_314_n1930), 
        .CO(div_DP_OP_279J39_124_314_n917), .S(div_DP_OP_279J39_124_314_n918)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U843 ( .A(div_DP_OP_279J39_124_314_n1994), .B(div_DP_OP_279J39_124_314_n937), .CI(div_DP_OP_279J39_124_314_n935), .CO(
        div_DP_OP_279J39_124_314_n915), .S(div_DP_OP_279J39_124_314_n916) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U842 ( .A(div_DP_OP_279J39_124_314_n933), 
        .B(div_DP_OP_279J39_124_314_n922), .CI(div_DP_OP_279J39_124_314_n918), 
        .CO(div_DP_OP_279J39_124_314_n913), .S(div_DP_OP_279J39_124_314_n914)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U841 ( .A(div_DP_OP_279J39_124_314_n920), 
        .B(div_DP_OP_279J39_124_314_n931), .CI(div_DP_OP_279J39_124_314_n929), 
        .CO(div_DP_OP_279J39_124_314_n911), .S(div_DP_OP_279J39_124_314_n912)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U840 ( .A(div_DP_OP_279J39_124_314_n916), 
        .B(div_DP_OP_279J39_124_314_n914), .CI(div_DP_OP_279J39_124_314_n927), 
        .CO(div_DP_OP_279J39_124_314_n909), .S(div_DP_OP_279J39_124_314_n910)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U839 ( .A(div_DP_OP_279J39_124_314_n912), 
        .B(div_DP_OP_279J39_124_314_n925), .CI(div_DP_OP_279J39_124_314_n910), 
        .CO(div_DP_OP_279J39_124_314_n907), .S(div_DP_OP_279J39_124_314_n908)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U838 ( .A(div_n_T_51_115_), .B(
        div_DP_OP_279J39_124_314_n1673), .CI(div_DP_OP_279J39_124_314_n2185), 
        .CO(div_DP_OP_279J39_124_314_n905), .S(div_DP_OP_279J39_124_314_n906)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U837 ( .A(div_DP_OP_279J39_124_314_n2121), .B(div_DP_OP_279J39_124_314_n1737), .CI(div_DP_OP_279J39_124_314_n1801), 
        .CO(div_DP_OP_279J39_124_314_n903), .S(div_DP_OP_279J39_124_314_n904)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U836 ( .A(div_DP_OP_279J39_124_314_n2057), .B(div_DP_OP_279J39_124_314_n1865), .CI(div_DP_OP_279J39_124_314_n1929), 
        .CO(div_DP_OP_279J39_124_314_n901), .S(div_DP_OP_279J39_124_314_n902)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U835 ( .A(div_DP_OP_279J39_124_314_n1993), .B(div_DP_OP_279J39_124_314_n921), .CI(div_DP_OP_279J39_124_314_n919), .CO(
        div_DP_OP_279J39_124_314_n899), .S(div_DP_OP_279J39_124_314_n900) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U834 ( .A(div_DP_OP_279J39_124_314_n917), 
        .B(div_DP_OP_279J39_124_314_n906), .CI(div_DP_OP_279J39_124_314_n902), 
        .CO(div_DP_OP_279J39_124_314_n897), .S(div_DP_OP_279J39_124_314_n898)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U833 ( .A(div_DP_OP_279J39_124_314_n904), 
        .B(div_DP_OP_279J39_124_314_n915), .CI(div_DP_OP_279J39_124_314_n913), 
        .CO(div_DP_OP_279J39_124_314_n895), .S(div_DP_OP_279J39_124_314_n896)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U832 ( .A(div_DP_OP_279J39_124_314_n900), 
        .B(div_DP_OP_279J39_124_314_n898), .CI(div_DP_OP_279J39_124_314_n911), 
        .CO(div_DP_OP_279J39_124_314_n893), .S(div_DP_OP_279J39_124_314_n894)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U831 ( .A(div_DP_OP_279J39_124_314_n896), 
        .B(div_DP_OP_279J39_124_314_n909), .CI(div_DP_OP_279J39_124_314_n894), 
        .CO(div_DP_OP_279J39_124_314_n891), .S(div_DP_OP_279J39_124_314_n892)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U830 ( .A(div_n_T_51_116_), .B(
        div_DP_OP_279J39_124_314_n1672), .CI(div_DP_OP_279J39_124_314_n2184), 
        .CO(div_DP_OP_279J39_124_314_n889), .S(div_DP_OP_279J39_124_314_n890)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U829 ( .A(div_DP_OP_279J39_124_314_n2120), .B(div_DP_OP_279J39_124_314_n1736), .CI(div_DP_OP_279J39_124_314_n1800), 
        .CO(div_DP_OP_279J39_124_314_n887), .S(div_DP_OP_279J39_124_314_n888)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U828 ( .A(div_DP_OP_279J39_124_314_n2056), .B(div_DP_OP_279J39_124_314_n1864), .CI(div_DP_OP_279J39_124_314_n1928), 
        .CO(div_DP_OP_279J39_124_314_n885), .S(div_DP_OP_279J39_124_314_n886)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U827 ( .A(div_DP_OP_279J39_124_314_n1992), .B(div_DP_OP_279J39_124_314_n905), .CI(div_DP_OP_279J39_124_314_n903), .CO(
        div_DP_OP_279J39_124_314_n883), .S(div_DP_OP_279J39_124_314_n884) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U826 ( .A(div_DP_OP_279J39_124_314_n901), 
        .B(div_DP_OP_279J39_124_314_n890), .CI(div_DP_OP_279J39_124_314_n886), 
        .CO(div_DP_OP_279J39_124_314_n881), .S(div_DP_OP_279J39_124_314_n882)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U825 ( .A(div_DP_OP_279J39_124_314_n888), 
        .B(div_DP_OP_279J39_124_314_n899), .CI(div_DP_OP_279J39_124_314_n897), 
        .CO(div_DP_OP_279J39_124_314_n879), .S(div_DP_OP_279J39_124_314_n880)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U824 ( .A(div_DP_OP_279J39_124_314_n884), 
        .B(div_DP_OP_279J39_124_314_n882), .CI(div_DP_OP_279J39_124_314_n895), 
        .CO(div_DP_OP_279J39_124_314_n877), .S(div_DP_OP_279J39_124_314_n878)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U823 ( .A(div_DP_OP_279J39_124_314_n880), 
        .B(div_DP_OP_279J39_124_314_n893), .CI(div_DP_OP_279J39_124_314_n878), 
        .CO(div_DP_OP_279J39_124_314_n875), .S(div_DP_OP_279J39_124_314_n876)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U822 ( .A(div_n_T_51_117_), .B(
        div_DP_OP_279J39_124_314_n1671), .CI(div_DP_OP_279J39_124_314_n2183), 
        .CO(div_DP_OP_279J39_124_314_n873), .S(div_DP_OP_279J39_124_314_n874)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U821 ( .A(div_DP_OP_279J39_124_314_n2119), .B(div_DP_OP_279J39_124_314_n1735), .CI(div_DP_OP_279J39_124_314_n1799), 
        .CO(div_DP_OP_279J39_124_314_n871), .S(div_DP_OP_279J39_124_314_n872)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U820 ( .A(div_DP_OP_279J39_124_314_n2055), .B(div_DP_OP_279J39_124_314_n1863), .CI(div_DP_OP_279J39_124_314_n1927), 
        .CO(div_DP_OP_279J39_124_314_n869), .S(div_DP_OP_279J39_124_314_n870)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U819 ( .A(div_DP_OP_279J39_124_314_n1991), .B(div_DP_OP_279J39_124_314_n889), .CI(div_DP_OP_279J39_124_314_n887), .CO(
        div_DP_OP_279J39_124_314_n867), .S(div_DP_OP_279J39_124_314_n868) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U818 ( .A(div_DP_OP_279J39_124_314_n885), 
        .B(div_DP_OP_279J39_124_314_n874), .CI(div_DP_OP_279J39_124_314_n870), 
        .CO(div_DP_OP_279J39_124_314_n865), .S(div_DP_OP_279J39_124_314_n866)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U817 ( .A(div_DP_OP_279J39_124_314_n872), 
        .B(div_DP_OP_279J39_124_314_n883), .CI(div_DP_OP_279J39_124_314_n881), 
        .CO(div_DP_OP_279J39_124_314_n863), .S(div_DP_OP_279J39_124_314_n864)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U816 ( .A(div_DP_OP_279J39_124_314_n868), 
        .B(div_DP_OP_279J39_124_314_n866), .CI(div_DP_OP_279J39_124_314_n879), 
        .CO(div_DP_OP_279J39_124_314_n861), .S(div_DP_OP_279J39_124_314_n862)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U815 ( .A(div_DP_OP_279J39_124_314_n864), 
        .B(div_DP_OP_279J39_124_314_n877), .CI(div_DP_OP_279J39_124_314_n862), 
        .CO(div_DP_OP_279J39_124_314_n859), .S(div_DP_OP_279J39_124_314_n860)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U814 ( .A(div_n_T_51_118_), .B(
        div_DP_OP_279J39_124_314_n1670), .CI(div_DP_OP_279J39_124_314_n2182), 
        .CO(div_DP_OP_279J39_124_314_n857), .S(div_DP_OP_279J39_124_314_n858)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U813 ( .A(div_DP_OP_279J39_124_314_n2118), .B(div_DP_OP_279J39_124_314_n1734), .CI(div_DP_OP_279J39_124_314_n1798), 
        .CO(div_DP_OP_279J39_124_314_n855), .S(div_DP_OP_279J39_124_314_n856)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U812 ( .A(div_DP_OP_279J39_124_314_n2054), .B(div_DP_OP_279J39_124_314_n1862), .CI(div_DP_OP_279J39_124_314_n1926), 
        .CO(div_DP_OP_279J39_124_314_n853), .S(div_DP_OP_279J39_124_314_n854)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U811 ( .A(div_DP_OP_279J39_124_314_n1990), .B(div_DP_OP_279J39_124_314_n873), .CI(div_DP_OP_279J39_124_314_n871), .CO(
        div_DP_OP_279J39_124_314_n851), .S(div_DP_OP_279J39_124_314_n852) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U810 ( .A(div_DP_OP_279J39_124_314_n869), 
        .B(div_DP_OP_279J39_124_314_n858), .CI(div_DP_OP_279J39_124_314_n854), 
        .CO(div_DP_OP_279J39_124_314_n849), .S(div_DP_OP_279J39_124_314_n850)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U809 ( .A(div_DP_OP_279J39_124_314_n856), 
        .B(div_DP_OP_279J39_124_314_n867), .CI(div_DP_OP_279J39_124_314_n865), 
        .CO(div_DP_OP_279J39_124_314_n847), .S(div_DP_OP_279J39_124_314_n848)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U808 ( .A(div_DP_OP_279J39_124_314_n852), 
        .B(div_DP_OP_279J39_124_314_n850), .CI(div_DP_OP_279J39_124_314_n863), 
        .CO(div_DP_OP_279J39_124_314_n845), .S(div_DP_OP_279J39_124_314_n846)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U807 ( .A(div_DP_OP_279J39_124_314_n848), 
        .B(div_DP_OP_279J39_124_314_n861), .CI(div_DP_OP_279J39_124_314_n846), 
        .CO(div_DP_OP_279J39_124_314_n843), .S(div_DP_OP_279J39_124_314_n844)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U806 ( .A(div_n_T_51_119_), .B(
        div_DP_OP_279J39_124_314_n1669), .CI(div_DP_OP_279J39_124_314_n2181), 
        .CO(div_DP_OP_279J39_124_314_n841), .S(div_DP_OP_279J39_124_314_n842)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U805 ( .A(div_DP_OP_279J39_124_314_n2117), .B(div_DP_OP_279J39_124_314_n1733), .CI(div_DP_OP_279J39_124_314_n1797), 
        .CO(div_DP_OP_279J39_124_314_n839), .S(div_DP_OP_279J39_124_314_n840)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U804 ( .A(div_DP_OP_279J39_124_314_n2053), .B(div_DP_OP_279J39_124_314_n1861), .CI(div_DP_OP_279J39_124_314_n1925), 
        .CO(div_DP_OP_279J39_124_314_n837), .S(div_DP_OP_279J39_124_314_n838)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U803 ( .A(div_DP_OP_279J39_124_314_n1989), .B(div_DP_OP_279J39_124_314_n857), .CI(div_DP_OP_279J39_124_314_n855), .CO(
        div_DP_OP_279J39_124_314_n835), .S(div_DP_OP_279J39_124_314_n836) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U802 ( .A(div_DP_OP_279J39_124_314_n853), 
        .B(div_DP_OP_279J39_124_314_n842), .CI(div_DP_OP_279J39_124_314_n838), 
        .CO(div_DP_OP_279J39_124_314_n833), .S(div_DP_OP_279J39_124_314_n834)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U801 ( .A(div_DP_OP_279J39_124_314_n840), 
        .B(div_DP_OP_279J39_124_314_n851), .CI(div_DP_OP_279J39_124_314_n849), 
        .CO(div_DP_OP_279J39_124_314_n831), .S(div_DP_OP_279J39_124_314_n832)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U800 ( .A(div_DP_OP_279J39_124_314_n836), 
        .B(div_DP_OP_279J39_124_314_n834), .CI(div_DP_OP_279J39_124_314_n847), 
        .CO(div_DP_OP_279J39_124_314_n829), .S(div_DP_OP_279J39_124_314_n830)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U799 ( .A(div_DP_OP_279J39_124_314_n832), 
        .B(div_DP_OP_279J39_124_314_n845), .CI(div_DP_OP_279J39_124_314_n830), 
        .CO(div_DP_OP_279J39_124_314_n827), .S(div_DP_OP_279J39_124_314_n828)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U798 ( .A(div_n_T_51_120_), .B(
        div_DP_OP_279J39_124_314_n1668), .CI(div_DP_OP_279J39_124_314_n2180), 
        .CO(div_DP_OP_279J39_124_314_n825), .S(div_DP_OP_279J39_124_314_n826)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U797 ( .A(div_DP_OP_279J39_124_314_n2116), .B(div_DP_OP_279J39_124_314_n1732), .CI(div_DP_OP_279J39_124_314_n1796), 
        .CO(div_DP_OP_279J39_124_314_n823), .S(div_DP_OP_279J39_124_314_n824)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U796 ( .A(div_DP_OP_279J39_124_314_n2052), .B(div_DP_OP_279J39_124_314_n1860), .CI(div_DP_OP_279J39_124_314_n1924), 
        .CO(div_DP_OP_279J39_124_314_n821), .S(div_DP_OP_279J39_124_314_n822)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U795 ( .A(div_DP_OP_279J39_124_314_n1988), .B(div_DP_OP_279J39_124_314_n841), .CI(div_DP_OP_279J39_124_314_n839), .CO(
        div_DP_OP_279J39_124_314_n819), .S(div_DP_OP_279J39_124_314_n820) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U794 ( .A(div_DP_OP_279J39_124_314_n837), 
        .B(div_DP_OP_279J39_124_314_n826), .CI(div_DP_OP_279J39_124_314_n822), 
        .CO(div_DP_OP_279J39_124_314_n817), .S(div_DP_OP_279J39_124_314_n818)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U793 ( .A(div_DP_OP_279J39_124_314_n824), 
        .B(div_DP_OP_279J39_124_314_n835), .CI(div_DP_OP_279J39_124_314_n833), 
        .CO(div_DP_OP_279J39_124_314_n815), .S(div_DP_OP_279J39_124_314_n816)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U792 ( .A(div_DP_OP_279J39_124_314_n820), 
        .B(div_DP_OP_279J39_124_314_n818), .CI(div_DP_OP_279J39_124_314_n831), 
        .CO(div_DP_OP_279J39_124_314_n813), .S(div_DP_OP_279J39_124_314_n814)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U791 ( .A(div_DP_OP_279J39_124_314_n816), 
        .B(div_DP_OP_279J39_124_314_n829), .CI(div_DP_OP_279J39_124_314_n814), 
        .CO(div_DP_OP_279J39_124_314_n811), .S(div_DP_OP_279J39_124_314_n812)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U790 ( .A(div_n_T_51_121_), .B(
        div_DP_OP_279J39_124_314_n1667), .CI(div_DP_OP_279J39_124_314_n2179), 
        .CO(div_DP_OP_279J39_124_314_n809), .S(div_DP_OP_279J39_124_314_n810)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U789 ( .A(div_DP_OP_279J39_124_314_n2115), .B(div_DP_OP_279J39_124_314_n1731), .CI(div_DP_OP_279J39_124_314_n1795), 
        .CO(div_DP_OP_279J39_124_314_n807), .S(div_DP_OP_279J39_124_314_n808)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U788 ( .A(div_DP_OP_279J39_124_314_n2051), .B(div_DP_OP_279J39_124_314_n1859), .CI(div_DP_OP_279J39_124_314_n1923), 
        .CO(div_DP_OP_279J39_124_314_n805), .S(div_DP_OP_279J39_124_314_n806)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U787 ( .A(div_DP_OP_279J39_124_314_n1987), .B(div_DP_OP_279J39_124_314_n825), .CI(div_DP_OP_279J39_124_314_n823), .CO(
        div_DP_OP_279J39_124_314_n803), .S(div_DP_OP_279J39_124_314_n804) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U786 ( .A(div_DP_OP_279J39_124_314_n821), 
        .B(div_DP_OP_279J39_124_314_n810), .CI(div_DP_OP_279J39_124_314_n806), 
        .CO(div_DP_OP_279J39_124_314_n801), .S(div_DP_OP_279J39_124_314_n802)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U785 ( .A(div_DP_OP_279J39_124_314_n808), 
        .B(div_DP_OP_279J39_124_314_n819), .CI(div_DP_OP_279J39_124_314_n817), 
        .CO(div_DP_OP_279J39_124_314_n799), .S(div_DP_OP_279J39_124_314_n800)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U784 ( .A(div_DP_OP_279J39_124_314_n804), 
        .B(div_DP_OP_279J39_124_314_n802), .CI(div_DP_OP_279J39_124_314_n815), 
        .CO(div_DP_OP_279J39_124_314_n797), .S(div_DP_OP_279J39_124_314_n798)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U783 ( .A(div_DP_OP_279J39_124_314_n800), 
        .B(div_DP_OP_279J39_124_314_n813), .CI(div_DP_OP_279J39_124_314_n798), 
        .CO(div_DP_OP_279J39_124_314_n795), .S(div_DP_OP_279J39_124_314_n796)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U782 ( .A(div_n_T_51_122_), .B(
        div_DP_OP_279J39_124_314_n1666), .CI(div_DP_OP_279J39_124_314_n2178), 
        .CO(div_DP_OP_279J39_124_314_n793), .S(div_DP_OP_279J39_124_314_n794)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U781 ( .A(div_DP_OP_279J39_124_314_n2114), .B(div_DP_OP_279J39_124_314_n1730), .CI(div_DP_OP_279J39_124_314_n1794), 
        .CO(div_DP_OP_279J39_124_314_n791), .S(div_DP_OP_279J39_124_314_n792)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U780 ( .A(div_DP_OP_279J39_124_314_n2050), .B(div_DP_OP_279J39_124_314_n1858), .CI(div_DP_OP_279J39_124_314_n1922), 
        .CO(div_DP_OP_279J39_124_314_n789), .S(div_DP_OP_279J39_124_314_n790)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U779 ( .A(div_DP_OP_279J39_124_314_n1986), .B(div_DP_OP_279J39_124_314_n809), .CI(div_DP_OP_279J39_124_314_n807), .CO(
        div_DP_OP_279J39_124_314_n787), .S(div_DP_OP_279J39_124_314_n788) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U778 ( .A(div_DP_OP_279J39_124_314_n805), 
        .B(div_DP_OP_279J39_124_314_n794), .CI(div_DP_OP_279J39_124_314_n790), 
        .CO(div_DP_OP_279J39_124_314_n785), .S(div_DP_OP_279J39_124_314_n786)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U777 ( .A(div_DP_OP_279J39_124_314_n792), 
        .B(div_DP_OP_279J39_124_314_n803), .CI(div_DP_OP_279J39_124_314_n801), 
        .CO(div_DP_OP_279J39_124_314_n783), .S(div_DP_OP_279J39_124_314_n784)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U776 ( .A(div_DP_OP_279J39_124_314_n788), 
        .B(div_DP_OP_279J39_124_314_n786), .CI(div_DP_OP_279J39_124_314_n799), 
        .CO(div_DP_OP_279J39_124_314_n781), .S(div_DP_OP_279J39_124_314_n782)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U775 ( .A(div_DP_OP_279J39_124_314_n784), 
        .B(div_DP_OP_279J39_124_314_n797), .CI(div_DP_OP_279J39_124_314_n782), 
        .CO(div_DP_OP_279J39_124_314_n779), .S(div_DP_OP_279J39_124_314_n780)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U774 ( .A(div_n_T_51_123_), .B(
        div_DP_OP_279J39_124_314_n1665), .CI(div_DP_OP_279J39_124_314_n2177), 
        .CO(div_DP_OP_279J39_124_314_n777), .S(div_DP_OP_279J39_124_314_n778)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U773 ( .A(div_DP_OP_279J39_124_314_n2113), .B(div_DP_OP_279J39_124_314_n1729), .CI(div_DP_OP_279J39_124_314_n1793), 
        .CO(div_DP_OP_279J39_124_314_n775), .S(div_DP_OP_279J39_124_314_n776)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U772 ( .A(div_DP_OP_279J39_124_314_n2049), .B(div_DP_OP_279J39_124_314_n1857), .CI(div_DP_OP_279J39_124_314_n1921), 
        .CO(div_DP_OP_279J39_124_314_n773), .S(div_DP_OP_279J39_124_314_n774)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U771 ( .A(div_DP_OP_279J39_124_314_n1985), .B(div_DP_OP_279J39_124_314_n793), .CI(div_DP_OP_279J39_124_314_n791), .CO(
        div_DP_OP_279J39_124_314_n771), .S(div_DP_OP_279J39_124_314_n772) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U770 ( .A(div_DP_OP_279J39_124_314_n789), 
        .B(div_DP_OP_279J39_124_314_n778), .CI(div_DP_OP_279J39_124_314_n774), 
        .CO(div_DP_OP_279J39_124_314_n769), .S(div_DP_OP_279J39_124_314_n770)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U769 ( .A(div_DP_OP_279J39_124_314_n776), 
        .B(div_DP_OP_279J39_124_314_n787), .CI(div_DP_OP_279J39_124_314_n785), 
        .CO(div_DP_OP_279J39_124_314_n767), .S(div_DP_OP_279J39_124_314_n768)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U768 ( .A(div_DP_OP_279J39_124_314_n772), 
        .B(div_DP_OP_279J39_124_314_n770), .CI(div_DP_OP_279J39_124_314_n783), 
        .CO(div_DP_OP_279J39_124_314_n765), .S(div_DP_OP_279J39_124_314_n766)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U767 ( .A(div_DP_OP_279J39_124_314_n768), 
        .B(div_DP_OP_279J39_124_314_n781), .CI(div_DP_OP_279J39_124_314_n766), 
        .CO(div_DP_OP_279J39_124_314_n763), .S(div_DP_OP_279J39_124_314_n764)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U766 ( .A(div_n_T_51_124_), .B(
        div_DP_OP_279J39_124_314_n1664), .CI(div_DP_OP_279J39_124_314_n2176), 
        .CO(div_DP_OP_279J39_124_314_n761), .S(div_DP_OP_279J39_124_314_n762)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U765 ( .A(div_DP_OP_279J39_124_314_n2112), .B(div_DP_OP_279J39_124_314_n1728), .CI(div_DP_OP_279J39_124_314_n1792), 
        .CO(div_DP_OP_279J39_124_314_n759), .S(div_DP_OP_279J39_124_314_n760)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U764 ( .A(div_DP_OP_279J39_124_314_n2048), .B(div_DP_OP_279J39_124_314_n1856), .CI(div_DP_OP_279J39_124_314_n1920), 
        .CO(div_DP_OP_279J39_124_314_n757), .S(div_DP_OP_279J39_124_314_n758)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U763 ( .A(div_DP_OP_279J39_124_314_n1984), .B(div_DP_OP_279J39_124_314_n777), .CI(div_DP_OP_279J39_124_314_n775), .CO(
        div_DP_OP_279J39_124_314_n755), .S(div_DP_OP_279J39_124_314_n756) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U762 ( .A(div_DP_OP_279J39_124_314_n773), 
        .B(div_DP_OP_279J39_124_314_n762), .CI(div_DP_OP_279J39_124_314_n758), 
        .CO(div_DP_OP_279J39_124_314_n753), .S(div_DP_OP_279J39_124_314_n754)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U761 ( .A(div_DP_OP_279J39_124_314_n760), 
        .B(div_DP_OP_279J39_124_314_n771), .CI(div_DP_OP_279J39_124_314_n769), 
        .CO(div_DP_OP_279J39_124_314_n751), .S(div_DP_OP_279J39_124_314_n752)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U760 ( .A(div_DP_OP_279J39_124_314_n756), 
        .B(div_DP_OP_279J39_124_314_n754), .CI(div_DP_OP_279J39_124_314_n767), 
        .CO(div_DP_OP_279J39_124_314_n749), .S(div_DP_OP_279J39_124_314_n750)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U759 ( .A(div_DP_OP_279J39_124_314_n752), 
        .B(div_DP_OP_279J39_124_314_n765), .CI(div_DP_OP_279J39_124_314_n750), 
        .CO(div_DP_OP_279J39_124_314_n747), .S(div_DP_OP_279J39_124_314_n748)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U758 ( .A(div_n_T_51_125_), .B(
        div_DP_OP_279J39_124_314_n1663), .CI(div_DP_OP_279J39_124_314_n2175), 
        .CO(div_DP_OP_279J39_124_314_n745), .S(div_DP_OP_279J39_124_314_n746)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U757 ( .A(div_DP_OP_279J39_124_314_n2111), .B(div_DP_OP_279J39_124_314_n1727), .CI(div_DP_OP_279J39_124_314_n1791), 
        .CO(div_DP_OP_279J39_124_314_n743), .S(div_DP_OP_279J39_124_314_n744)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U756 ( .A(div_DP_OP_279J39_124_314_n2047), .B(div_DP_OP_279J39_124_314_n1855), .CI(div_DP_OP_279J39_124_314_n1919), 
        .CO(div_DP_OP_279J39_124_314_n741), .S(div_DP_OP_279J39_124_314_n742)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U755 ( .A(div_DP_OP_279J39_124_314_n1983), .B(div_DP_OP_279J39_124_314_n761), .CI(div_DP_OP_279J39_124_314_n759), .CO(
        div_DP_OP_279J39_124_314_n739), .S(div_DP_OP_279J39_124_314_n740) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U754 ( .A(div_DP_OP_279J39_124_314_n757), 
        .B(div_DP_OP_279J39_124_314_n746), .CI(div_DP_OP_279J39_124_314_n742), 
        .CO(div_DP_OP_279J39_124_314_n737), .S(div_DP_OP_279J39_124_314_n738)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U753 ( .A(div_DP_OP_279J39_124_314_n744), 
        .B(div_DP_OP_279J39_124_314_n755), .CI(div_DP_OP_279J39_124_314_n753), 
        .CO(div_DP_OP_279J39_124_314_n735), .S(div_DP_OP_279J39_124_314_n736)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U752 ( .A(div_DP_OP_279J39_124_314_n740), 
        .B(div_DP_OP_279J39_124_314_n738), .CI(div_DP_OP_279J39_124_314_n751), 
        .CO(div_DP_OP_279J39_124_314_n733), .S(div_DP_OP_279J39_124_314_n734)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U751 ( .A(div_DP_OP_279J39_124_314_n736), 
        .B(div_DP_OP_279J39_124_314_n749), .CI(div_DP_OP_279J39_124_314_n734), 
        .CO(div_DP_OP_279J39_124_314_n731), .S(div_DP_OP_279J39_124_314_n732)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U750 ( .A(div_n_T_51_126_), .B(
        div_DP_OP_279J39_124_314_n1662), .CI(div_DP_OP_279J39_124_314_n2174), 
        .CO(div_DP_OP_279J39_124_314_n729), .S(div_DP_OP_279J39_124_314_n730)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U749 ( .A(div_DP_OP_279J39_124_314_n2110), .B(div_DP_OP_279J39_124_314_n1726), .CI(div_DP_OP_279J39_124_314_n1790), 
        .CO(div_DP_OP_279J39_124_314_n727), .S(div_DP_OP_279J39_124_314_n728)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U748 ( .A(div_DP_OP_279J39_124_314_n2046), .B(div_DP_OP_279J39_124_314_n1854), .CI(div_DP_OP_279J39_124_314_n1918), 
        .CO(div_DP_OP_279J39_124_314_n725), .S(div_DP_OP_279J39_124_314_n726)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U747 ( .A(div_DP_OP_279J39_124_314_n1982), .B(div_DP_OP_279J39_124_314_n745), .CI(div_DP_OP_279J39_124_314_n743), .CO(
        div_DP_OP_279J39_124_314_n723), .S(div_DP_OP_279J39_124_314_n724) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U746 ( .A(div_DP_OP_279J39_124_314_n741), 
        .B(div_DP_OP_279J39_124_314_n730), .CI(div_DP_OP_279J39_124_314_n726), 
        .CO(div_DP_OP_279J39_124_314_n721), .S(div_DP_OP_279J39_124_314_n722)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U745 ( .A(div_DP_OP_279J39_124_314_n728), 
        .B(div_DP_OP_279J39_124_314_n739), .CI(div_DP_OP_279J39_124_314_n737), 
        .CO(div_DP_OP_279J39_124_314_n719), .S(div_DP_OP_279J39_124_314_n720)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U744 ( .A(div_DP_OP_279J39_124_314_n724), 
        .B(div_DP_OP_279J39_124_314_n722), .CI(div_DP_OP_279J39_124_314_n735), 
        .CO(div_DP_OP_279J39_124_314_n717), .S(div_DP_OP_279J39_124_314_n718)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U743 ( .A(div_DP_OP_279J39_124_314_n720), 
        .B(div_DP_OP_279J39_124_314_n733), .CI(div_DP_OP_279J39_124_314_n718), 
        .CO(div_DP_OP_279J39_124_314_n715), .S(div_DP_OP_279J39_124_314_n716)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U742 ( .A(div_n_T_51_127_), .B(
        div_DP_OP_279J39_124_314_n1661), .CI(div_DP_OP_279J39_124_314_n2173), 
        .CO(div_DP_OP_279J39_124_314_n713), .S(div_DP_OP_279J39_124_314_n714)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U741 ( .A(div_DP_OP_279J39_124_314_n2109), .B(div_DP_OP_279J39_124_314_n1725), .CI(div_DP_OP_279J39_124_314_n1789), 
        .CO(div_DP_OP_279J39_124_314_n711), .S(div_DP_OP_279J39_124_314_n712)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U740 ( .A(div_DP_OP_279J39_124_314_n2045), .B(div_DP_OP_279J39_124_314_n1853), .CI(div_DP_OP_279J39_124_314_n1917), 
        .CO(div_DP_OP_279J39_124_314_n709), .S(div_DP_OP_279J39_124_314_n710)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U739 ( .A(div_DP_OP_279J39_124_314_n1981), .B(div_DP_OP_279J39_124_314_n729), .CI(div_DP_OP_279J39_124_314_n727), .CO(
        div_DP_OP_279J39_124_314_n707), .S(div_DP_OP_279J39_124_314_n708) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U738 ( .A(div_DP_OP_279J39_124_314_n725), 
        .B(div_DP_OP_279J39_124_314_n714), .CI(div_DP_OP_279J39_124_314_n710), 
        .CO(div_DP_OP_279J39_124_314_n705), .S(div_DP_OP_279J39_124_314_n706)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U737 ( .A(div_DP_OP_279J39_124_314_n712), 
        .B(div_DP_OP_279J39_124_314_n723), .CI(div_DP_OP_279J39_124_314_n721), 
        .CO(div_DP_OP_279J39_124_314_n703), .S(div_DP_OP_279J39_124_314_n704)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U736 ( .A(div_DP_OP_279J39_124_314_n708), 
        .B(div_DP_OP_279J39_124_314_n706), .CI(div_DP_OP_279J39_124_314_n719), 
        .CO(div_DP_OP_279J39_124_314_n701), .S(div_DP_OP_279J39_124_314_n702)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U735 ( .A(div_DP_OP_279J39_124_314_n704), 
        .B(div_DP_OP_279J39_124_314_n717), .CI(div_DP_OP_279J39_124_314_n702), 
        .CO(div_DP_OP_279J39_124_314_n699), .S(div_DP_OP_279J39_124_314_n700)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U734 ( .A(div_DP_OP_279J39_124_314_n2587), .B(div_DP_OP_279J39_124_314_n1660), .CI(div_DP_OP_279J39_124_314_n2172), 
        .CO(div_DP_OP_279J39_124_314_n697), .S(div_DP_OP_279J39_124_314_n698)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U733 ( .A(div_DP_OP_279J39_124_314_n2108), .B(div_DP_OP_279J39_124_314_n1724), .CI(div_DP_OP_279J39_124_314_n1788), 
        .CO(div_DP_OP_279J39_124_314_n695), .S(div_DP_OP_279J39_124_314_n696)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U732 ( .A(div_DP_OP_279J39_124_314_n2044), .B(div_DP_OP_279J39_124_314_n1852), .CI(div_DP_OP_279J39_124_314_n1916), 
        .CO(div_DP_OP_279J39_124_314_n693), .S(div_DP_OP_279J39_124_314_n694)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U731 ( .A(div_DP_OP_279J39_124_314_n1980), .B(div_DP_OP_279J39_124_314_n713), .CI(div_DP_OP_279J39_124_314_n711), .CO(
        div_DP_OP_279J39_124_314_n691), .S(div_DP_OP_279J39_124_314_n692) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U730 ( .A(div_DP_OP_279J39_124_314_n709), 
        .B(div_DP_OP_279J39_124_314_n698), .CI(div_DP_OP_279J39_124_314_n694), 
        .CO(div_DP_OP_279J39_124_314_n689), .S(div_DP_OP_279J39_124_314_n690)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U729 ( .A(div_DP_OP_279J39_124_314_n696), 
        .B(div_DP_OP_279J39_124_314_n707), .CI(div_DP_OP_279J39_124_314_n705), 
        .CO(div_DP_OP_279J39_124_314_n687), .S(div_DP_OP_279J39_124_314_n688)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U728 ( .A(div_DP_OP_279J39_124_314_n692), 
        .B(div_DP_OP_279J39_124_314_n690), .CI(div_DP_OP_279J39_124_314_n703), 
        .CO(div_DP_OP_279J39_124_314_n685), .S(div_DP_OP_279J39_124_314_n686)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U727 ( .A(div_DP_OP_279J39_124_314_n688), 
        .B(div_DP_OP_279J39_124_314_n701), .CI(div_DP_OP_279J39_124_314_n686), 
        .CO(div_DP_OP_279J39_124_314_n683), .S(div_DP_OP_279J39_124_314_n684)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U726 ( .A(div_DP_OP_279J39_124_314_n2107), .B(div_DP_OP_279J39_124_314_n1659), .CI(div_DP_OP_279J39_124_314_n2043), 
        .CO(div_DP_OP_279J39_124_314_n681), .S(div_DP_OP_279J39_124_314_n682)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U725 ( .A(div_DP_OP_279J39_124_314_n1979), .B(div_DP_OP_279J39_124_314_n1723), .CI(div_DP_OP_279J39_124_314_n1787), 
        .CO(div_DP_OP_279J39_124_314_n679), .S(div_DP_OP_279J39_124_314_n680)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U724 ( .A(div_DP_OP_279J39_124_314_n1915), .B(div_DP_OP_279J39_124_314_n1851), .CI(div_DP_OP_279J39_124_314_n697), .CO(
        div_DP_OP_279J39_124_314_n677), .S(div_DP_OP_279J39_124_314_n678) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U723 ( .A(div_DP_OP_279J39_124_314_n695), 
        .B(div_DP_OP_279J39_124_314_n693), .CI(div_DP_OP_279J39_124_314_n682), 
        .CO(div_DP_OP_279J39_124_314_n675), .S(div_DP_OP_279J39_124_314_n676)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U722 ( .A(div_DP_OP_279J39_124_314_n680), 
        .B(div_DP_OP_279J39_124_314_n691), .CI(div_DP_OP_279J39_124_314_n678), 
        .CO(div_DP_OP_279J39_124_314_n673), .S(div_DP_OP_279J39_124_314_n674)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U721 ( .A(div_DP_OP_279J39_124_314_n689), 
        .B(div_DP_OP_279J39_124_314_n676), .CI(div_DP_OP_279J39_124_314_n687), 
        .CO(div_DP_OP_279J39_124_314_n671), .S(div_DP_OP_279J39_124_314_n672)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U720 ( .A(div_DP_OP_279J39_124_314_n674), 
        .B(div_DP_OP_279J39_124_314_n685), .CI(div_DP_OP_279J39_124_314_n672), 
        .CO(div_DP_OP_279J39_124_314_n669), .S(div_DP_OP_279J39_124_314_n670)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U719 ( .A(div_DP_OP_279J39_124_314_n2042), .B(div_DP_OP_279J39_124_314_n1658), .CI(div_DP_OP_279J39_124_314_n1978), 
        .CO(div_DP_OP_279J39_124_314_n667), .S(div_DP_OP_279J39_124_314_n668)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U718 ( .A(div_DP_OP_279J39_124_314_n1722), .B(div_DP_OP_279J39_124_314_n1914), .CI(div_DP_OP_279J39_124_314_n1850), 
        .CO(div_DP_OP_279J39_124_314_n665), .S(div_DP_OP_279J39_124_314_n666)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U717 ( .A(div_DP_OP_279J39_124_314_n1786), .B(div_DP_OP_279J39_124_314_n681), .CI(div_DP_OP_279J39_124_314_n679), .CO(
        div_DP_OP_279J39_124_314_n663), .S(div_DP_OP_279J39_124_314_n664) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U716 ( .A(div_DP_OP_279J39_124_314_n668), 
        .B(div_DP_OP_279J39_124_314_n666), .CI(div_DP_OP_279J39_124_314_n677), 
        .CO(div_DP_OP_279J39_124_314_n661), .S(div_DP_OP_279J39_124_314_n662)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U715 ( .A(div_DP_OP_279J39_124_314_n675), 
        .B(div_DP_OP_279J39_124_314_n664), .CI(div_DP_OP_279J39_124_314_n673), 
        .CO(div_DP_OP_279J39_124_314_n659), .S(div_DP_OP_279J39_124_314_n660)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U714 ( .A(div_DP_OP_279J39_124_314_n662), 
        .B(div_DP_OP_279J39_124_314_n671), .CI(div_DP_OP_279J39_124_314_n660), 
        .CO(div_DP_OP_279J39_124_314_n657), .S(div_DP_OP_279J39_124_314_n658)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U713 ( .A(div_DP_OP_279J39_124_314_n1977), .B(div_DP_OP_279J39_124_314_n1657), .CI(div_DP_OP_279J39_124_314_n1913), 
        .CO(div_DP_OP_279J39_124_314_n655), .S(div_DP_OP_279J39_124_314_n656)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U712 ( .A(div_DP_OP_279J39_124_314_n1721), .B(div_DP_OP_279J39_124_314_n1785), .CI(div_DP_OP_279J39_124_314_n1849), 
        .CO(div_DP_OP_279J39_124_314_n653), .S(div_DP_OP_279J39_124_314_n654)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U711 ( .A(div_DP_OP_279J39_124_314_n667), 
        .B(div_DP_OP_279J39_124_314_n665), .CI(div_DP_OP_279J39_124_314_n656), 
        .CO(div_DP_OP_279J39_124_314_n651), .S(div_DP_OP_279J39_124_314_n652)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U710 ( .A(div_DP_OP_279J39_124_314_n654), 
        .B(div_DP_OP_279J39_124_314_n663), .CI(div_DP_OP_279J39_124_314_n661), 
        .CO(div_DP_OP_279J39_124_314_n649), .S(div_DP_OP_279J39_124_314_n650)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U709 ( .A(div_DP_OP_279J39_124_314_n652), 
        .B(div_DP_OP_279J39_124_314_n659), .CI(div_DP_OP_279J39_124_314_n650), 
        .CO(div_DP_OP_279J39_124_314_n647), .S(div_DP_OP_279J39_124_314_n648)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U708 ( .A(div_DP_OP_279J39_124_314_n1912), .B(div_DP_OP_279J39_124_314_n1656), .CI(div_DP_OP_279J39_124_314_n1848), 
        .CO(div_DP_OP_279J39_124_314_n645), .S(div_DP_OP_279J39_124_314_n646)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U707 ( .A(div_DP_OP_279J39_124_314_n1784), .B(div_DP_OP_279J39_124_314_n1720), .CI(div_DP_OP_279J39_124_314_n655), .CO(
        div_DP_OP_279J39_124_314_n643), .S(div_DP_OP_279J39_124_314_n644) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U706 ( .A(div_DP_OP_279J39_124_314_n653), 
        .B(div_DP_OP_279J39_124_314_n646), .CI(div_DP_OP_279J39_124_314_n644), 
        .CO(div_DP_OP_279J39_124_314_n641), .S(div_DP_OP_279J39_124_314_n642)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U705 ( .A(div_DP_OP_279J39_124_314_n651), 
        .B(div_DP_OP_279J39_124_314_n649), .CI(div_DP_OP_279J39_124_314_n642), 
        .CO(div_DP_OP_279J39_124_314_n639), .S(div_DP_OP_279J39_124_314_n640)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U704 ( .A(div_DP_OP_279J39_124_314_n1847), .B(div_DP_OP_279J39_124_314_n1655), .CI(div_DP_OP_279J39_124_314_n1783), 
        .CO(div_DP_OP_279J39_124_314_n637), .S(div_DP_OP_279J39_124_314_n638)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U703 ( .A(div_DP_OP_279J39_124_314_n1719), .B(div_DP_OP_279J39_124_314_n645), .CI(div_DP_OP_279J39_124_314_n638), .CO(
        div_DP_OP_279J39_124_314_n635), .S(div_DP_OP_279J39_124_314_n636) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U702 ( .A(div_DP_OP_279J39_124_314_n643), 
        .B(div_DP_OP_279J39_124_314_n636), .CI(div_DP_OP_279J39_124_314_n641), 
        .CO(div_DP_OP_279J39_124_314_n633), .S(div_DP_OP_279J39_124_314_n634)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U701 ( .A(div_DP_OP_279J39_124_314_n1782), .B(div_DP_OP_279J39_124_314_n1654), .CI(div_DP_OP_279J39_124_314_n1718), 
        .CO(div_DP_OP_279J39_124_314_n631), .S(div_DP_OP_279J39_124_314_n632)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U700 ( .A(div_DP_OP_279J39_124_314_n637), 
        .B(div_DP_OP_279J39_124_314_n632), .CI(div_DP_OP_279J39_124_314_n635), 
        .CO(div_DP_OP_279J39_124_314_n629), .S(div_DP_OP_279J39_124_314_n630)
         );
  FADDX1_LVT div_DP_OP_279J39_124_314_U699 ( .A(div_DP_OP_279J39_124_314_n1717), .B(div_DP_OP_279J39_124_314_n1653), .CI(div_DP_OP_279J39_124_314_n631), .CO(
        div_DP_OP_279J39_124_314_n627), .S(div_DP_OP_279J39_124_314_n628) );
  FADDX1_LVT div_DP_OP_279J39_124_314_U692 ( .A(div_DP_OP_279J39_124_314_n2171), .B(div_DP_OP_279J39_124_314_n2586), .CI(div_DP_OP_279J39_124_314_n1650), 
        .CO(div_DP_OP_279J39_124_314_n551), .S(div_n_T_65[1]) );
  AND4X1_LVT div_ash_111_U1030 ( .A1(div_n302), .A2(div_ash_111_n683), .A3(
        div_ash_111_n684), .A4(div_ash_111_n679), .Y(div_ash_111_n846) );
  AND3X1_LVT div_ash_111_U1029 ( .A1(div_ash_111_n846), .A2(div_ash_111_n681), 
        .A3(div_ash_111_n682), .Y(div_ash_111_n885) );
  AO22X1_LVT div_ash_111_U1028 ( .A1(div_n171), .A2(div_n_T_51_37_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_38_), .Y(div_ash_111_n858) );
  AO22X1_LVT div_ash_111_U1027 ( .A1(div_n171), .A2(div_n_T_51_39_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_40_), .Y(div_ash_111_n1037) );
  AO22X1_LVT div_ash_111_U1026 ( .A1(div_n166), .A2(div_ash_111_n858), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1037), .Y(div_ash_111_n844) );
  AO22X1_LVT div_ash_111_U1025 ( .A1(div_n171), .A2(div_n_T_51_41_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_42_), .Y(div_ash_111_n1038) );
  AO22X1_LVT div_ash_111_U1024 ( .A1(div_n171), .A2(div_n_T_51_43_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_44_), .Y(div_ash_111_n1035) );
  AO22X1_LVT div_ash_111_U1023 ( .A1(div_n166), .A2(div_ash_111_n1038), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1035), .Y(div_ash_111_n1013) );
  AO22X1_LVT div_ash_111_U1022 ( .A1(div_n167), .A2(div_ash_111_n844), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1013), .Y(div_ash_111_n824) );
  AO22X1_LVT div_ash_111_U1021 ( .A1(div_n171), .A2(div_n_T_51_45_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_46_), .Y(div_ash_111_n1036) );
  AO22X1_LVT div_ash_111_U1020 ( .A1(div_n171), .A2(div_n_T_51_47_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_48_), .Y(div_ash_111_n1033) );
  AO22X1_LVT div_ash_111_U1019 ( .A1(div_n166), .A2(div_ash_111_n1036), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1033), .Y(div_ash_111_n1014) );
  AO22X1_LVT div_ash_111_U1018 ( .A1(div_n171), .A2(div_n_T_51_49_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_50_), .Y(div_ash_111_n1034) );
  AO22X1_LVT div_ash_111_U1017 ( .A1(div_n171), .A2(div_n_T_51_51_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_52_), .Y(div_ash_111_n1031) );
  AO22X1_LVT div_ash_111_U1016 ( .A1(div_n166), .A2(div_ash_111_n1034), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1031), .Y(div_ash_111_n1011) );
  AO22X1_LVT div_ash_111_U1015 ( .A1(div_n167), .A2(div_ash_111_n1014), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1011), .Y(div_ash_111_n994) );
  AO22X1_LVT div_ash_111_U1014 ( .A1(div_n168), .A2(div_ash_111_n824), .A3(
        div_ash_111_n682), .A4(div_ash_111_n994), .Y(div_ash_111_n791) );
  AO22X1_LVT div_ash_111_U1013 ( .A1(div_n171), .A2(div_n_T_51_61_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_62_), .Y(div_ash_111_n1028) );
  OA222X1_LVT div_ash_111_U1012 ( .A1(div_n166), .A2(div_n171), .A3(div_n166), 
        .A4(div_n_T_51_63_), .A5(div_ash_111_n684), .A6(div_ash_111_n1028), 
        .Y(div_ash_111_n993) );
  AO22X1_LVT div_ash_111_U1011 ( .A1(div_n171), .A2(div_n_T_51_53_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_54_), .Y(div_ash_111_n1032) );
  AO22X1_LVT div_ash_111_U1010 ( .A1(div_n171), .A2(div_n_T_51_55_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_56_), .Y(div_ash_111_n1029) );
  AO22X1_LVT div_ash_111_U1009 ( .A1(div_n166), .A2(div_ash_111_n1032), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1029), .Y(div_ash_111_n1012) );
  AO22X1_LVT div_ash_111_U1008 ( .A1(div_n171), .A2(div_n_T_51_57_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_58_), .Y(div_ash_111_n1030) );
  AO22X1_LVT div_ash_111_U1007 ( .A1(div_n171), .A2(div_n_T_51_59_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_60_), .Y(div_ash_111_n1027) );
  AO22X1_LVT div_ash_111_U1006 ( .A1(div_n166), .A2(div_ash_111_n1030), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1027), .Y(div_ash_111_n1015) );
  AO22X1_LVT div_ash_111_U1005 ( .A1(div_n167), .A2(div_ash_111_n1012), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1015), .Y(div_ash_111_n995) );
  OA222X1_LVT div_ash_111_U1004 ( .A1(div_n168), .A2(div_n167), .A3(div_n168), 
        .A4(div_ash_111_n993), .A5(div_ash_111_n682), .A6(div_ash_111_n995), 
        .Y(div_ash_111_n712) );
  AO22X1_LVT div_ash_111_U1003 ( .A1(div_n169), .A2(div_ash_111_n791), .A3(
        div_ash_111_n681), .A4(div_ash_111_n712), .Y(div_ash_111_n747) );
  AND2X1_LVT div_ash_111_U1002 ( .A1(div_n170), .A2(div_ash_111_n747), .Y(
        div_n_T_442[100]) );
  AO22X1_LVT div_ash_111_U1001 ( .A1(div_n171), .A2(div_n_T_51_38_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_39_), .Y(div_ash_111_n852) );
  AO22X1_LVT div_ash_111_U1000 ( .A1(div_n171), .A2(div_n_T_51_40_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_41_), .Y(div_ash_111_n1022) );
  AO22X1_LVT div_ash_111_U999 ( .A1(div_n166), .A2(div_ash_111_n852), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1022), .Y(div_ash_111_n838) );
  AO22X1_LVT div_ash_111_U998 ( .A1(div_n171), .A2(div_n_T_51_42_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_43_), .Y(div_ash_111_n1023) );
  AO22X1_LVT div_ash_111_U997 ( .A1(div_n171), .A2(div_n_T_51_44_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_45_), .Y(div_ash_111_n1020) );
  AO22X1_LVT div_ash_111_U996 ( .A1(div_n166), .A2(div_ash_111_n1023), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1020), .Y(div_ash_111_n1007) );
  AO22X1_LVT div_ash_111_U995 ( .A1(div_n167), .A2(div_ash_111_n838), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1007), .Y(div_ash_111_n820) );
  AO22X1_LVT div_ash_111_U994 ( .A1(div_n171), .A2(div_n_T_51_46_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_47_), .Y(div_ash_111_n1021) );
  AO22X1_LVT div_ash_111_U993 ( .A1(div_n171), .A2(div_n_T_51_48_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_49_), .Y(div_ash_111_n1018) );
  AO22X1_LVT div_ash_111_U992 ( .A1(div_n166), .A2(div_ash_111_n1021), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1018), .Y(div_ash_111_n1008) );
  AO22X1_LVT div_ash_111_U991 ( .A1(div_n171), .A2(div_n_T_51_50_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_51_), .Y(div_ash_111_n1019) );
  AO22X1_LVT div_ash_111_U990 ( .A1(div_n171), .A2(div_n_T_51_52_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_53_), .Y(div_ash_111_n1016) );
  AO22X1_LVT div_ash_111_U989 ( .A1(div_n166), .A2(div_ash_111_n1019), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1016), .Y(div_ash_111_n1005) );
  AO22X1_LVT div_ash_111_U988 ( .A1(div_n167), .A2(div_ash_111_n1008), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1005), .Y(div_ash_111_n991) );
  AO22X1_LVT div_ash_111_U987 ( .A1(div_n168), .A2(div_ash_111_n820), .A3(
        div_ash_111_n682), .A4(div_ash_111_n991), .Y(div_ash_111_n788) );
  AO22X1_LVT div_ash_111_U986 ( .A1(div_n171), .A2(div_n_T_51_54_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_55_), .Y(div_ash_111_n1017) );
  AO22X1_LVT div_ash_111_U985 ( .A1(div_n171), .A2(div_n_T_51_56_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_57_), .Y(div_ash_111_n1025) );
  AO22X1_LVT div_ash_111_U984 ( .A1(div_n166), .A2(div_ash_111_n1017), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1025), .Y(div_ash_111_n1006) );
  AO22X1_LVT div_ash_111_U983 ( .A1(div_n171), .A2(div_n_T_51_58_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_59_), .Y(div_ash_111_n1026) );
  AO22X1_LVT div_ash_111_U982 ( .A1(div_n171), .A2(div_n_T_51_60_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_61_), .Y(div_ash_111_n1024) );
  AO22X1_LVT div_ash_111_U981 ( .A1(div_n166), .A2(div_ash_111_n1026), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1024), .Y(div_ash_111_n1010) );
  AO22X1_LVT div_ash_111_U980 ( .A1(div_n167), .A2(div_ash_111_n1006), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1010), .Y(div_ash_111_n992) );
  AO22X1_LVT div_ash_111_U979 ( .A1(div_n171), .A2(div_n_T_51_62_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_63_), .Y(div_ash_111_n1009) );
  AND3X1_LVT div_ash_111_U978 ( .A1(div_n166), .A2(div_n167), .A3(
        div_ash_111_n1009), .Y(div_ash_111_n976) );
  AO22X1_LVT div_ash_111_U977 ( .A1(div_n168), .A2(div_ash_111_n992), .A3(
        div_ash_111_n682), .A4(div_ash_111_n976), .Y(div_ash_111_n710) );
  AO22X1_LVT div_ash_111_U976 ( .A1(div_n169), .A2(div_ash_111_n788), .A3(
        div_ash_111_n681), .A4(div_ash_111_n710), .Y(div_ash_111_n745) );
  AND2X1_LVT div_ash_111_U975 ( .A1(div_n170), .A2(div_ash_111_n745), .Y(
        div_n_T_442[101]) );
  AO22X1_LVT div_ash_111_U974 ( .A1(div_n166), .A2(div_ash_111_n1037), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1038), .Y(div_ash_111_n834) );
  AO22X1_LVT div_ash_111_U973 ( .A1(div_n166), .A2(div_ash_111_n1035), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1036), .Y(div_ash_111_n1002) );
  AO22X1_LVT div_ash_111_U972 ( .A1(div_n167), .A2(div_ash_111_n834), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1002), .Y(div_ash_111_n816) );
  AO22X1_LVT div_ash_111_U971 ( .A1(div_n166), .A2(div_ash_111_n1033), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1034), .Y(div_ash_111_n1003) );
  AO22X1_LVT div_ash_111_U970 ( .A1(div_n166), .A2(div_ash_111_n1031), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1032), .Y(div_ash_111_n1000) );
  AO22X1_LVT div_ash_111_U969 ( .A1(div_n167), .A2(div_ash_111_n1003), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1000), .Y(div_ash_111_n989) );
  AO22X1_LVT div_ash_111_U968 ( .A1(div_n168), .A2(div_ash_111_n816), .A3(
        div_ash_111_n682), .A4(div_ash_111_n989), .Y(div_ash_111_n785) );
  AND3X1_LVT div_ash_111_U967 ( .A1(div_n166), .A2(div_n171), .A3(
        div_n_T_51_63_), .Y(div_ash_111_n988) );
  AO22X1_LVT div_ash_111_U966 ( .A1(div_n166), .A2(div_ash_111_n1029), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1030), .Y(div_ash_111_n1001) );
  AO22X1_LVT div_ash_111_U965 ( .A1(div_n166), .A2(div_ash_111_n1027), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1028), .Y(div_ash_111_n1004) );
  AO22X1_LVT div_ash_111_U964 ( .A1(div_n167), .A2(div_ash_111_n1001), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1004), .Y(div_ash_111_n990) );
  OA222X1_LVT div_ash_111_U963 ( .A1(div_n168), .A2(div_n167), .A3(div_n168), 
        .A4(div_ash_111_n988), .A5(div_ash_111_n682), .A6(div_ash_111_n990), 
        .Y(div_ash_111_n708) );
  AO22X1_LVT div_ash_111_U962 ( .A1(div_n169), .A2(div_ash_111_n785), .A3(
        div_ash_111_n681), .A4(div_ash_111_n708), .Y(div_ash_111_n742) );
  AND2X1_LVT div_ash_111_U961 ( .A1(div_n170), .A2(div_ash_111_n742), .Y(
        div_n_T_442[102]) );
  AO22X1_LVT div_ash_111_U960 ( .A1(div_n166), .A2(div_ash_111_n1025), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1026), .Y(div_ash_111_n997) );
  AO22X1_LVT div_ash_111_U959 ( .A1(div_n166), .A2(div_ash_111_n1024), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1009), .Y(div_ash_111_n982) );
  AO22X1_LVT div_ash_111_U958 ( .A1(div_n167), .A2(div_ash_111_n997), .A3(
        div_ash_111_n683), .A4(div_ash_111_n982), .Y(div_ash_111_n981) );
  AO22X1_LVT div_ash_111_U957 ( .A1(div_n166), .A2(div_ash_111_n1022), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1023), .Y(div_ash_111_n829) );
  AO22X1_LVT div_ash_111_U956 ( .A1(div_n166), .A2(div_ash_111_n1020), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1021), .Y(div_ash_111_n998) );
  AO22X1_LVT div_ash_111_U955 ( .A1(div_n167), .A2(div_ash_111_n829), .A3(
        div_ash_111_n683), .A4(div_ash_111_n998), .Y(div_ash_111_n812) );
  AO22X1_LVT div_ash_111_U954 ( .A1(div_n166), .A2(div_ash_111_n1018), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1019), .Y(div_ash_111_n999) );
  AO22X1_LVT div_ash_111_U953 ( .A1(div_n166), .A2(div_ash_111_n1016), .A3(
        div_ash_111_n684), .A4(div_ash_111_n1017), .Y(div_ash_111_n996) );
  AO22X1_LVT div_ash_111_U952 ( .A1(div_n167), .A2(div_ash_111_n999), .A3(
        div_ash_111_n683), .A4(div_ash_111_n996), .Y(div_ash_111_n987) );
  AO22X1_LVT div_ash_111_U951 ( .A1(div_n168), .A2(div_ash_111_n812), .A3(
        div_ash_111_n682), .A4(div_ash_111_n987), .Y(div_ash_111_n782) );
  OA222X1_LVT div_ash_111_U950 ( .A1(div_n169), .A2(div_n168), .A3(div_n169), 
        .A4(div_ash_111_n981), .A5(div_ash_111_n681), .A6(div_ash_111_n782), 
        .Y(div_ash_111_n740) );
  AND2X1_LVT div_ash_111_U949 ( .A1(div_n170), .A2(div_ash_111_n740), .Y(
        div_n_T_442[103]) );
  AO22X1_LVT div_ash_111_U948 ( .A1(div_n167), .A2(div_ash_111_n1015), .A3(
        div_ash_111_n683), .A4(div_ash_111_n993), .Y(div_ash_111_n979) );
  AO22X1_LVT div_ash_111_U947 ( .A1(div_n167), .A2(div_ash_111_n1013), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1014), .Y(div_ash_111_n808) );
  AO22X1_LVT div_ash_111_U946 ( .A1(div_n167), .A2(div_ash_111_n1011), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1012), .Y(div_ash_111_n986) );
  AO22X1_LVT div_ash_111_U945 ( .A1(div_n168), .A2(div_ash_111_n808), .A3(
        div_ash_111_n682), .A4(div_ash_111_n986), .Y(div_ash_111_n779) );
  OA222X1_LVT div_ash_111_U944 ( .A1(div_n169), .A2(div_n168), .A3(div_n169), 
        .A4(div_ash_111_n979), .A5(div_ash_111_n681), .A6(div_ash_111_n779), 
        .Y(div_ash_111_n738) );
  AND2X1_LVT div_ash_111_U943 ( .A1(div_n170), .A2(div_ash_111_n738), .Y(
        div_n_T_442[104]) );
  OA222X1_LVT div_ash_111_U942 ( .A1(div_n167), .A2(div_n166), .A3(div_n167), 
        .A4(div_ash_111_n1009), .A5(div_ash_111_n683), .A6(div_ash_111_n1010), 
        .Y(div_ash_111_n978) );
  AO22X1_LVT div_ash_111_U941 ( .A1(div_n167), .A2(div_ash_111_n1007), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1008), .Y(div_ash_111_n804) );
  AO22X1_LVT div_ash_111_U940 ( .A1(div_n167), .A2(div_ash_111_n1005), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1006), .Y(div_ash_111_n985) );
  AO22X1_LVT div_ash_111_U939 ( .A1(div_n168), .A2(div_ash_111_n804), .A3(
        div_ash_111_n682), .A4(div_ash_111_n985), .Y(div_ash_111_n776) );
  OA222X1_LVT div_ash_111_U938 ( .A1(div_n169), .A2(div_n168), .A3(div_n169), 
        .A4(div_ash_111_n978), .A5(div_ash_111_n681), .A6(div_ash_111_n776), 
        .Y(div_ash_111_n736) );
  AND2X1_LVT div_ash_111_U937 ( .A1(div_n170), .A2(div_ash_111_n736), .Y(
        div_n_T_442[105]) );
  AO22X1_LVT div_ash_111_U936 ( .A1(div_n167), .A2(div_ash_111_n1004), .A3(
        div_ash_111_n683), .A4(div_ash_111_n988), .Y(div_ash_111_n977) );
  AO22X1_LVT div_ash_111_U935 ( .A1(div_n167), .A2(div_ash_111_n1002), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1003), .Y(div_ash_111_n799) );
  AO22X1_LVT div_ash_111_U934 ( .A1(div_n167), .A2(div_ash_111_n1000), .A3(
        div_ash_111_n683), .A4(div_ash_111_n1001), .Y(div_ash_111_n984) );
  AO22X1_LVT div_ash_111_U933 ( .A1(div_n168), .A2(div_ash_111_n799), .A3(
        div_ash_111_n682), .A4(div_ash_111_n984), .Y(div_ash_111_n773) );
  OA222X1_LVT div_ash_111_U932 ( .A1(div_n169), .A2(div_n168), .A3(div_n169), 
        .A4(div_ash_111_n977), .A5(div_ash_111_n681), .A6(div_ash_111_n773), 
        .Y(div_ash_111_n734) );
  AND2X1_LVT div_ash_111_U931 ( .A1(div_n170), .A2(div_ash_111_n734), .Y(
        div_n_T_442[106]) );
  AO22X1_LVT div_ash_111_U930 ( .A1(div_n167), .A2(div_ash_111_n998), .A3(
        div_ash_111_n683), .A4(div_ash_111_n999), .Y(div_ash_111_n795) );
  AO22X1_LVT div_ash_111_U929 ( .A1(div_n167), .A2(div_ash_111_n996), .A3(
        div_ash_111_n683), .A4(div_ash_111_n997), .Y(div_ash_111_n983) );
  AO22X1_LVT div_ash_111_U928 ( .A1(div_n168), .A2(div_ash_111_n795), .A3(
        div_ash_111_n682), .A4(div_ash_111_n983), .Y(div_ash_111_n770) );
  AND3X1_LVT div_ash_111_U927 ( .A1(div_n167), .A2(div_n168), .A3(
        div_ash_111_n982), .Y(div_ash_111_n697) );
  AO22X1_LVT div_ash_111_U926 ( .A1(div_n169), .A2(div_ash_111_n770), .A3(
        div_ash_111_n681), .A4(div_ash_111_n697), .Y(div_ash_111_n732) );
  AND2X1_LVT div_ash_111_U925 ( .A1(div_n170), .A2(div_ash_111_n732), .Y(
        div_n_T_442[107]) );
  AO22X1_LVT div_ash_111_U924 ( .A1(div_n168), .A2(div_ash_111_n994), .A3(
        div_ash_111_n682), .A4(div_ash_111_n995), .Y(div_ash_111_n766) );
  AND3X1_LVT div_ash_111_U923 ( .A1(div_n167), .A2(div_n168), .A3(
        div_ash_111_n993), .Y(div_ash_111_n695) );
  AO22X1_LVT div_ash_111_U922 ( .A1(div_n169), .A2(div_ash_111_n766), .A3(
        div_ash_111_n681), .A4(div_ash_111_n695), .Y(div_ash_111_n730) );
  AND2X1_LVT div_ash_111_U921 ( .A1(div_n170), .A2(div_ash_111_n730), .Y(
        div_n_T_442[108]) );
  AO22X1_LVT div_ash_111_U920 ( .A1(div_n168), .A2(div_ash_111_n991), .A3(
        div_ash_111_n682), .A4(div_ash_111_n992), .Y(div_ash_111_n763) );
  OA222X1_LVT div_ash_111_U919 ( .A1(div_n169), .A2(div_n168), .A3(div_n169), 
        .A4(div_ash_111_n976), .A5(div_ash_111_n681), .A6(div_ash_111_n763), 
        .Y(div_ash_111_n728) );
  AND2X1_LVT div_ash_111_U918 ( .A1(div_n170), .A2(div_ash_111_n728), .Y(
        div_n_T_442[109]) );
  AO22X1_LVT div_ash_111_U917 ( .A1(div_n171), .A2(div_n305), .A3(
        div_ash_111_n679), .A4(div_n306), .Y(div_ash_111_n972) );
  AO22X1_LVT div_ash_111_U916 ( .A1(div_n171), .A2(div_n_T_51_5_), .A3(
        div_ash_111_n679), .A4(div_n307), .Y(div_ash_111_n974) );
  AO22X1_LVT div_ash_111_U915 ( .A1(div_n166), .A2(div_ash_111_n972), .A3(
        div_ash_111_n684), .A4(div_ash_111_n974), .Y(div_ash_111_n937) );
  AO22X1_LVT div_ash_111_U914 ( .A1(div_n171), .A2(div_n_T_51_7_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_8_), .Y(div_ash_111_n975) );
  AO22X1_LVT div_ash_111_U913 ( .A1(div_n171), .A2(div_n_T_51_9_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_10_), .Y(div_ash_111_n973) );
  AO22X1_LVT div_ash_111_U912 ( .A1(div_n166), .A2(div_ash_111_n975), .A3(
        div_ash_111_n684), .A4(div_ash_111_n973), .Y(div_ash_111_n962) );
  AO22X1_LVT div_ash_111_U911 ( .A1(div_n167), .A2(div_ash_111_n937), .A3(
        div_ash_111_n683), .A4(div_ash_111_n962), .Y(div_ash_111_n920) );
  AO22X1_LVT div_ash_111_U910 ( .A1(div_n171), .A2(div_n303), .A3(
        div_ash_111_n679), .A4(div_n304), .Y(div_ash_111_n971) );
  OA222X1_LVT div_ash_111_U909 ( .A1(div_ash_111_n684), .A2(div_n302), .A3(
        div_ash_111_n684), .A4(div_ash_111_n679), .A5(div_n166), .A6(
        div_ash_111_n971), .Y(div_ash_111_n938) );
  AND2X1_LVT div_ash_111_U908 ( .A1(div_ash_111_n683), .A2(div_ash_111_n938), 
        .Y(div_ash_111_n919) );
  OA221X1_LVT div_ash_111_U907 ( .A1(div_n168), .A2(div_ash_111_n920), .A3(
        div_ash_111_n682), .A4(div_ash_111_n919), .A5(div_ash_111_n681), .Y(
        div_ash_111_n830) );
  AND2X1_LVT div_ash_111_U906 ( .A1(div_ash_111_n830), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[10]) );
  AO22X1_LVT div_ash_111_U905 ( .A1(div_n168), .A2(div_ash_111_n989), .A3(
        div_ash_111_n682), .A4(div_ash_111_n990), .Y(div_ash_111_n760) );
  AND3X1_LVT div_ash_111_U904 ( .A1(div_n168), .A2(div_n167), .A3(
        div_ash_111_n988), .Y(div_ash_111_n691) );
  AO22X1_LVT div_ash_111_U903 ( .A1(div_n169), .A2(div_ash_111_n760), .A3(
        div_ash_111_n681), .A4(div_ash_111_n691), .Y(div_ash_111_n726) );
  AND2X1_LVT div_ash_111_U902 ( .A1(div_n170), .A2(div_ash_111_n726), .Y(
        div_n_T_442[110]) );
  AO22X1_LVT div_ash_111_U901 ( .A1(div_n168), .A2(div_ash_111_n987), .A3(
        div_ash_111_n682), .A4(div_ash_111_n981), .Y(div_ash_111_n723) );
  AND3X1_LVT div_ash_111_U900 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n723), .Y(div_n_T_442[111]) );
  AO22X1_LVT div_ash_111_U899 ( .A1(div_n168), .A2(div_ash_111_n986), .A3(
        div_ash_111_n682), .A4(div_ash_111_n979), .Y(div_ash_111_n720) );
  AND3X1_LVT div_ash_111_U898 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n720), .Y(div_n_T_442[112]) );
  AO22X1_LVT div_ash_111_U897 ( .A1(div_n168), .A2(div_ash_111_n985), .A3(
        div_ash_111_n682), .A4(div_ash_111_n978), .Y(div_ash_111_n718) );
  AND3X1_LVT div_ash_111_U896 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n718), .Y(div_n_T_442[113]) );
  AO22X1_LVT div_ash_111_U895 ( .A1(div_n168), .A2(div_ash_111_n984), .A3(
        div_ash_111_n682), .A4(div_ash_111_n977), .Y(div_ash_111_n716) );
  AND3X1_LVT div_ash_111_U894 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n716), .Y(div_n_T_442[114]) );
  OA222X1_LVT div_ash_111_U893 ( .A1(div_n168), .A2(div_n167), .A3(div_n168), 
        .A4(div_ash_111_n982), .A5(div_ash_111_n682), .A6(div_ash_111_n983), 
        .Y(div_ash_111_n714) );
  AND3X1_LVT div_ash_111_U892 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n714), .Y(div_n_T_442[115]) );
  AND3X1_LVT div_ash_111_U891 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n712), .Y(div_n_T_442[116]) );
  AND3X1_LVT div_ash_111_U890 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n710), .Y(div_n_T_442[117]) );
  AND3X1_LVT div_ash_111_U889 ( .A1(div_n169), .A2(div_n170), .A3(
        div_ash_111_n708), .Y(div_n_T_442[118]) );
  AND3X1_LVT div_ash_111_U888 ( .A1(div_n168), .A2(div_n169), .A3(
        div_ash_111_n981), .Y(div_ash_111_n707) );
  AND2X1_LVT div_ash_111_U887 ( .A1(div_n170), .A2(div_ash_111_n707), .Y(
        div_n_T_442[119]) );
  AO22X1_LVT div_ash_111_U886 ( .A1(div_n171), .A2(div_n306), .A3(
        div_ash_111_n679), .A4(div_n_T_51_5_), .Y(div_ash_111_n969) );
  AO22X1_LVT div_ash_111_U885 ( .A1(div_n171), .A2(div_n307), .A3(
        div_ash_111_n679), .A4(div_n_T_51_7_), .Y(div_ash_111_n966) );
  AO22X1_LVT div_ash_111_U884 ( .A1(div_n166), .A2(div_ash_111_n969), .A3(
        div_ash_111_n684), .A4(div_ash_111_n966), .Y(div_ash_111_n932) );
  AO22X1_LVT div_ash_111_U883 ( .A1(div_n171), .A2(div_n_T_51_8_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_9_), .Y(div_ash_111_n967) );
  AO22X1_LVT div_ash_111_U882 ( .A1(div_n171), .A2(div_n_T_51_10_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_11_), .Y(div_ash_111_n965) );
  AO22X1_LVT div_ash_111_U881 ( .A1(div_n166), .A2(div_ash_111_n967), .A3(
        div_ash_111_n684), .A4(div_ash_111_n965), .Y(div_ash_111_n959) );
  AO22X1_LVT div_ash_111_U880 ( .A1(div_n167), .A2(div_ash_111_n932), .A3(
        div_ash_111_n683), .A4(div_ash_111_n959), .Y(div_ash_111_n914) );
  AO22X1_LVT div_ash_111_U879 ( .A1(div_n171), .A2(div_n302), .A3(
        div_ash_111_n679), .A4(div_n303), .Y(div_ash_111_n980) );
  AO22X1_LVT div_ash_111_U878 ( .A1(div_n171), .A2(div_n304), .A3(
        div_ash_111_n679), .A4(div_n305), .Y(div_ash_111_n968) );
  AO22X1_LVT div_ash_111_U877 ( .A1(div_n166), .A2(div_ash_111_n980), .A3(
        div_ash_111_n684), .A4(div_ash_111_n968), .Y(div_ash_111_n933) );
  AND2X1_LVT div_ash_111_U876 ( .A1(div_ash_111_n683), .A2(div_ash_111_n933), 
        .Y(div_ash_111_n913) );
  OA221X1_LVT div_ash_111_U875 ( .A1(div_n168), .A2(div_ash_111_n914), .A3(
        div_ash_111_n682), .A4(div_ash_111_n913), .A5(div_ash_111_n681), .Y(
        div_ash_111_n825) );
  AND2X1_LVT div_ash_111_U874 ( .A1(div_ash_111_n825), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[11]) );
  AND3X1_LVT div_ash_111_U873 ( .A1(div_n168), .A2(div_n169), .A3(
        div_ash_111_n979), .Y(div_ash_111_n705) );
  AND2X1_LVT div_ash_111_U872 ( .A1(div_n170), .A2(div_ash_111_n705), .Y(
        div_n_T_442[120]) );
  AND3X1_LVT div_ash_111_U871 ( .A1(div_n168), .A2(div_n169), .A3(
        div_ash_111_n978), .Y(div_ash_111_n703) );
  AND2X1_LVT div_ash_111_U870 ( .A1(div_n170), .A2(div_ash_111_n703), .Y(
        div_n_T_442[121]) );
  AND3X1_LVT div_ash_111_U869 ( .A1(div_n168), .A2(div_n169), .A3(
        div_ash_111_n977), .Y(div_ash_111_n700) );
  AND2X1_LVT div_ash_111_U868 ( .A1(div_n170), .A2(div_ash_111_n700), .Y(
        div_n_T_442[122]) );
  AND3X1_LVT div_ash_111_U867 ( .A1(div_n170), .A2(div_n169), .A3(
        div_ash_111_n697), .Y(div_n_T_442[123]) );
  AND3X1_LVT div_ash_111_U866 ( .A1(div_n170), .A2(div_n169), .A3(
        div_ash_111_n695), .Y(div_n_T_442[124]) );
  AND3X1_LVT div_ash_111_U865 ( .A1(div_n169), .A2(div_n168), .A3(
        div_ash_111_n976), .Y(div_ash_111_n694) );
  AND2X1_LVT div_ash_111_U864 ( .A1(div_n170), .A2(div_ash_111_n694), .Y(
        div_n_T_442[125]) );
  AND3X1_LVT div_ash_111_U863 ( .A1(div_n170), .A2(div_n169), .A3(
        div_ash_111_n691), .Y(div_n_T_442[126]) );
  AO22X1_LVT div_ash_111_U862 ( .A1(div_n166), .A2(div_ash_111_n974), .A3(
        div_ash_111_n684), .A4(div_ash_111_n975), .Y(div_ash_111_n957) );
  AO22X1_LVT div_ash_111_U861 ( .A1(div_n171), .A2(div_n_T_51_11_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_12_), .Y(div_ash_111_n963) );
  AO22X1_LVT div_ash_111_U860 ( .A1(div_n166), .A2(div_ash_111_n973), .A3(
        div_ash_111_n684), .A4(div_ash_111_n963), .Y(div_ash_111_n954) );
  AO22X1_LVT div_ash_111_U859 ( .A1(div_n167), .A2(div_ash_111_n957), .A3(
        div_ash_111_n683), .A4(div_ash_111_n954), .Y(div_ash_111_n908) );
  AND3X1_LVT div_ash_111_U858 ( .A1(div_n302), .A2(div_ash_111_n684), .A3(
        div_ash_111_n679), .Y(div_ash_111_n970) );
  AO22X1_LVT div_ash_111_U857 ( .A1(div_n166), .A2(div_ash_111_n971), .A3(
        div_ash_111_n684), .A4(div_ash_111_n972), .Y(div_ash_111_n956) );
  AO22X1_LVT div_ash_111_U856 ( .A1(div_n167), .A2(div_ash_111_n970), .A3(
        div_ash_111_n683), .A4(div_ash_111_n956), .Y(div_ash_111_n907) );
  OA221X1_LVT div_ash_111_U855 ( .A1(div_n168), .A2(div_ash_111_n908), .A3(
        div_ash_111_n682), .A4(div_ash_111_n907), .A5(div_ash_111_n681), .Y(
        div_ash_111_n821) );
  OA221X1_LVT div_ash_111_U854 ( .A1(div_n171), .A2(div_n303), .A3(
        div_ash_111_n679), .A4(div_n302), .A5(div_ash_111_n684), .Y(
        div_ash_111_n943) );
  AO22X1_LVT div_ash_111_U853 ( .A1(div_n166), .A2(div_ash_111_n968), .A3(
        div_ash_111_n684), .A4(div_ash_111_n969), .Y(div_ash_111_n942) );
  AO22X1_LVT div_ash_111_U852 ( .A1(div_n167), .A2(div_ash_111_n943), .A3(
        div_ash_111_n683), .A4(div_ash_111_n942), .Y(div_ash_111_n964) );
  AO22X1_LVT div_ash_111_U851 ( .A1(div_n166), .A2(div_ash_111_n966), .A3(
        div_ash_111_n684), .A4(div_ash_111_n967), .Y(div_ash_111_n953) );
  AO22X1_LVT div_ash_111_U850 ( .A1(div_n171), .A2(div_n_T_51_12_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_13_), .Y(div_ash_111_n960) );
  AO22X1_LVT div_ash_111_U849 ( .A1(div_n166), .A2(div_ash_111_n965), .A3(
        div_ash_111_n684), .A4(div_ash_111_n960), .Y(div_ash_111_n951) );
  AO22X1_LVT div_ash_111_U848 ( .A1(div_n167), .A2(div_ash_111_n953), .A3(
        div_ash_111_n683), .A4(div_ash_111_n951), .Y(div_ash_111_n939) );
  AO22X1_LVT div_ash_111_U847 ( .A1(div_n168), .A2(div_ash_111_n964), .A3(
        div_ash_111_n682), .A4(div_ash_111_n939), .Y(div_ash_111_n899) );
  AND2X1_LVT div_ash_111_U846 ( .A1(div_ash_111_n681), .A2(div_ash_111_n899), 
        .Y(div_ash_111_n817) );
  AND2X1_LVT div_ash_111_U845 ( .A1(div_ash_111_n817), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[13]) );
  AO22X1_LVT div_ash_111_U844 ( .A1(div_n167), .A2(div_ash_111_n938), .A3(
        div_ash_111_n683), .A4(div_ash_111_n937), .Y(div_ash_111_n961) );
  AO22X1_LVT div_ash_111_U843 ( .A1(div_n171), .A2(div_n_T_51_13_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_14_), .Y(div_ash_111_n955) );
  AO22X1_LVT div_ash_111_U842 ( .A1(div_n166), .A2(div_ash_111_n963), .A3(
        div_ash_111_n684), .A4(div_ash_111_n955), .Y(div_ash_111_n949) );
  AO22X1_LVT div_ash_111_U841 ( .A1(div_n167), .A2(div_ash_111_n962), .A3(
        div_ash_111_n683), .A4(div_ash_111_n949), .Y(div_ash_111_n934) );
  AO22X1_LVT div_ash_111_U840 ( .A1(div_n168), .A2(div_ash_111_n961), .A3(
        div_ash_111_n682), .A4(div_ash_111_n934), .Y(div_ash_111_n894) );
  AND2X1_LVT div_ash_111_U839 ( .A1(div_ash_111_n681), .A2(div_ash_111_n894), 
        .Y(div_ash_111_n813) );
  AND2X1_LVT div_ash_111_U838 ( .A1(div_ash_111_n813), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[14]) );
  AO22X1_LVT div_ash_111_U837 ( .A1(div_n167), .A2(div_ash_111_n933), .A3(
        div_ash_111_n683), .A4(div_ash_111_n932), .Y(div_ash_111_n958) );
  AO22X1_LVT div_ash_111_U836 ( .A1(div_n171), .A2(div_n_T_51_14_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_15_), .Y(div_ash_111_n952) );
  AO22X1_LVT div_ash_111_U835 ( .A1(div_n166), .A2(div_ash_111_n960), .A3(
        div_ash_111_n684), .A4(div_ash_111_n952), .Y(div_ash_111_n947) );
  AO22X1_LVT div_ash_111_U834 ( .A1(div_n167), .A2(div_ash_111_n959), .A3(
        div_ash_111_n683), .A4(div_ash_111_n947), .Y(div_ash_111_n929) );
  AO22X1_LVT div_ash_111_U833 ( .A1(div_n168), .A2(div_ash_111_n958), .A3(
        div_ash_111_n682), .A4(div_ash_111_n929), .Y(div_ash_111_n890) );
  AND2X1_LVT div_ash_111_U832 ( .A1(div_ash_111_n681), .A2(div_ash_111_n890), 
        .Y(div_ash_111_n809) );
  AND2X1_LVT div_ash_111_U831 ( .A1(div_ash_111_n809), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[15]) );
  AO22X1_LVT div_ash_111_U830 ( .A1(div_n167), .A2(div_ash_111_n956), .A3(
        div_ash_111_n683), .A4(div_ash_111_n957), .Y(div_ash_111_n845) );
  AO22X1_LVT div_ash_111_U829 ( .A1(div_n171), .A2(div_n_T_51_15_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_16_), .Y(div_ash_111_n950) );
  AO22X1_LVT div_ash_111_U828 ( .A1(div_n166), .A2(div_ash_111_n955), .A3(
        div_ash_111_n684), .A4(div_ash_111_n950), .Y(div_ash_111_n944) );
  AO22X1_LVT div_ash_111_U827 ( .A1(div_n167), .A2(div_ash_111_n954), .A3(
        div_ash_111_n683), .A4(div_ash_111_n944), .Y(div_ash_111_n926) );
  AO22X1_LVT div_ash_111_U826 ( .A1(div_n168), .A2(div_ash_111_n845), .A3(
        div_ash_111_n682), .A4(div_ash_111_n926), .Y(div_ash_111_n886) );
  OA222X1_LVT div_ash_111_U825 ( .A1(div_ash_111_n681), .A2(div_ash_111_n846), 
        .A3(div_ash_111_n681), .A4(div_ash_111_n682), .A5(div_n169), .A6(
        div_ash_111_n886), .Y(div_ash_111_n805) );
  AND2X1_LVT div_ash_111_U824 ( .A1(div_ash_111_n943), .A2(div_ash_111_n683), 
        .Y(div_ash_111_n840) );
  AND2X1_LVT div_ash_111_U823 ( .A1(div_ash_111_n840), .A2(div_ash_111_n682), 
        .Y(div_ash_111_n946) );
  AO22X1_LVT div_ash_111_U822 ( .A1(div_n167), .A2(div_ash_111_n942), .A3(
        div_ash_111_n683), .A4(div_ash_111_n953), .Y(div_ash_111_n839) );
  AO22X1_LVT div_ash_111_U821 ( .A1(div_n171), .A2(div_n_T_51_16_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_17_), .Y(div_ash_111_n948) );
  AO22X1_LVT div_ash_111_U820 ( .A1(div_n166), .A2(div_ash_111_n952), .A3(
        div_ash_111_n684), .A4(div_ash_111_n948), .Y(div_ash_111_n940) );
  AO22X1_LVT div_ash_111_U819 ( .A1(div_n167), .A2(div_ash_111_n951), .A3(
        div_ash_111_n683), .A4(div_ash_111_n940), .Y(div_ash_111_n922) );
  AO22X1_LVT div_ash_111_U818 ( .A1(div_n168), .A2(div_ash_111_n839), .A3(
        div_ash_111_n682), .A4(div_ash_111_n922), .Y(div_ash_111_n881) );
  AO22X1_LVT div_ash_111_U817 ( .A1(div_n169), .A2(div_ash_111_n946), .A3(
        div_ash_111_n681), .A4(div_ash_111_n881), .Y(div_ash_111_n801) );
  AND2X1_LVT div_ash_111_U816 ( .A1(div_ash_111_n680), .A2(div_ash_111_n801), 
        .Y(div_n_T_442[17]) );
  AND2X1_LVT div_ash_111_U815 ( .A1(div_ash_111_n919), .A2(div_ash_111_n682), 
        .Y(div_ash_111_n898) );
  AO22X1_LVT div_ash_111_U814 ( .A1(div_n171), .A2(div_n_T_51_17_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_18_), .Y(div_ash_111_n945) );
  AO22X1_LVT div_ash_111_U813 ( .A1(div_n166), .A2(div_ash_111_n950), .A3(
        div_ash_111_n684), .A4(div_ash_111_n945), .Y(div_ash_111_n935) );
  AO22X1_LVT div_ash_111_U812 ( .A1(div_n167), .A2(div_ash_111_n949), .A3(
        div_ash_111_n683), .A4(div_ash_111_n935), .Y(div_ash_111_n916) );
  AO22X1_LVT div_ash_111_U811 ( .A1(div_n168), .A2(div_ash_111_n920), .A3(
        div_ash_111_n682), .A4(div_ash_111_n916), .Y(div_ash_111_n876) );
  AO22X1_LVT div_ash_111_U810 ( .A1(div_n169), .A2(div_ash_111_n898), .A3(
        div_ash_111_n681), .A4(div_ash_111_n876), .Y(div_ash_111_n796) );
  AND2X1_LVT div_ash_111_U809 ( .A1(div_ash_111_n680), .A2(div_ash_111_n796), 
        .Y(div_n_T_442[18]) );
  AND2X1_LVT div_ash_111_U808 ( .A1(div_ash_111_n913), .A2(div_ash_111_n682), 
        .Y(div_ash_111_n874) );
  AO22X1_LVT div_ash_111_U807 ( .A1(div_n171), .A2(div_n_T_51_18_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_19_), .Y(div_ash_111_n941) );
  AO22X1_LVT div_ash_111_U806 ( .A1(div_n166), .A2(div_ash_111_n948), .A3(
        div_ash_111_n684), .A4(div_ash_111_n941), .Y(div_ash_111_n930) );
  AO22X1_LVT div_ash_111_U805 ( .A1(div_n167), .A2(div_ash_111_n947), .A3(
        div_ash_111_n683), .A4(div_ash_111_n930), .Y(div_ash_111_n910) );
  AO22X1_LVT div_ash_111_U804 ( .A1(div_n168), .A2(div_ash_111_n914), .A3(
        div_ash_111_n682), .A4(div_ash_111_n910), .Y(div_ash_111_n870) );
  AO22X1_LVT div_ash_111_U803 ( .A1(div_n169), .A2(div_ash_111_n874), .A3(
        div_ash_111_n681), .A4(div_ash_111_n870), .Y(div_ash_111_n792) );
  AND2X1_LVT div_ash_111_U802 ( .A1(div_ash_111_n680), .A2(div_ash_111_n792), 
        .Y(div_n_T_442[19]) );
  AND2X1_LVT div_ash_111_U801 ( .A1(div_ash_111_n946), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n880) );
  AND2X1_LVT div_ash_111_U800 ( .A1(div_ash_111_n682), .A2(div_ash_111_n907), 
        .Y(div_ash_111_n869) );
  AO22X1_LVT div_ash_111_U799 ( .A1(div_n171), .A2(div_n_T_51_19_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_20_), .Y(div_ash_111_n936) );
  AO22X1_LVT div_ash_111_U798 ( .A1(div_n166), .A2(div_ash_111_n945), .A3(
        div_ash_111_n684), .A4(div_ash_111_n936), .Y(div_ash_111_n927) );
  AO22X1_LVT div_ash_111_U797 ( .A1(div_n167), .A2(div_ash_111_n944), .A3(
        div_ash_111_n683), .A4(div_ash_111_n927), .Y(div_ash_111_n904) );
  AO22X1_LVT div_ash_111_U796 ( .A1(div_n168), .A2(div_ash_111_n908), .A3(
        div_ash_111_n682), .A4(div_ash_111_n904), .Y(div_ash_111_n865) );
  AO22X1_LVT div_ash_111_U795 ( .A1(div_n169), .A2(div_ash_111_n869), .A3(
        div_ash_111_n681), .A4(div_ash_111_n865), .Y(div_ash_111_n789) );
  AND2X1_LVT div_ash_111_U794 ( .A1(div_ash_111_n680), .A2(div_ash_111_n789), 
        .Y(div_n_T_442[20]) );
  OA221X1_LVT div_ash_111_U793 ( .A1(div_n167), .A2(div_ash_111_n942), .A3(
        div_ash_111_n683), .A4(div_ash_111_n943), .A5(div_ash_111_n682), .Y(
        div_ash_111_n864) );
  AO22X1_LVT div_ash_111_U792 ( .A1(div_n171), .A2(div_n_T_51_20_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_21_), .Y(div_ash_111_n931) );
  AO22X1_LVT div_ash_111_U791 ( .A1(div_n166), .A2(div_ash_111_n941), .A3(
        div_ash_111_n684), .A4(div_ash_111_n931), .Y(div_ash_111_n923) );
  AO22X1_LVT div_ash_111_U790 ( .A1(div_n167), .A2(div_ash_111_n940), .A3(
        div_ash_111_n683), .A4(div_ash_111_n923), .Y(div_ash_111_n900) );
  AO22X1_LVT div_ash_111_U789 ( .A1(div_n168), .A2(div_ash_111_n939), .A3(
        div_ash_111_n682), .A4(div_ash_111_n900), .Y(div_ash_111_n860) );
  AO22X1_LVT div_ash_111_U788 ( .A1(div_n169), .A2(div_ash_111_n864), .A3(
        div_ash_111_n681), .A4(div_ash_111_n860), .Y(div_ash_111_n786) );
  AND2X1_LVT div_ash_111_U787 ( .A1(div_ash_111_n680), .A2(div_ash_111_n786), 
        .Y(div_n_T_442[21]) );
  OA221X1_LVT div_ash_111_U786 ( .A1(div_n167), .A2(div_ash_111_n937), .A3(
        div_ash_111_n683), .A4(div_ash_111_n938), .A5(div_ash_111_n682), .Y(
        div_ash_111_n859) );
  AO22X1_LVT div_ash_111_U785 ( .A1(div_n171), .A2(div_n_T_51_21_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_22_), .Y(div_ash_111_n928) );
  AO22X1_LVT div_ash_111_U784 ( .A1(div_n166), .A2(div_ash_111_n936), .A3(
        div_ash_111_n684), .A4(div_ash_111_n928), .Y(div_ash_111_n917) );
  AO22X1_LVT div_ash_111_U783 ( .A1(div_n167), .A2(div_ash_111_n935), .A3(
        div_ash_111_n683), .A4(div_ash_111_n917), .Y(div_ash_111_n895) );
  AO22X1_LVT div_ash_111_U782 ( .A1(div_n168), .A2(div_ash_111_n934), .A3(
        div_ash_111_n682), .A4(div_ash_111_n895), .Y(div_ash_111_n854) );
  AO22X1_LVT div_ash_111_U781 ( .A1(div_n169), .A2(div_ash_111_n859), .A3(
        div_ash_111_n681), .A4(div_ash_111_n854), .Y(div_ash_111_n783) );
  AND2X1_LVT div_ash_111_U780 ( .A1(div_ash_111_n680), .A2(div_ash_111_n783), 
        .Y(div_n_T_442[22]) );
  OA221X1_LVT div_ash_111_U779 ( .A1(div_n167), .A2(div_ash_111_n932), .A3(
        div_ash_111_n683), .A4(div_ash_111_n933), .A5(div_ash_111_n682), .Y(
        div_ash_111_n853) );
  AO22X1_LVT div_ash_111_U778 ( .A1(div_n171), .A2(div_n_T_51_22_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_23_), .Y(div_ash_111_n924) );
  AO22X1_LVT div_ash_111_U777 ( .A1(div_n166), .A2(div_ash_111_n931), .A3(
        div_ash_111_n684), .A4(div_ash_111_n924), .Y(div_ash_111_n911) );
  AO22X1_LVT div_ash_111_U776 ( .A1(div_n167), .A2(div_ash_111_n930), .A3(
        div_ash_111_n683), .A4(div_ash_111_n911), .Y(div_ash_111_n891) );
  AO22X1_LVT div_ash_111_U775 ( .A1(div_n168), .A2(div_ash_111_n929), .A3(
        div_ash_111_n682), .A4(div_ash_111_n891), .Y(div_ash_111_n848) );
  AO22X1_LVT div_ash_111_U774 ( .A1(div_n169), .A2(div_ash_111_n853), .A3(
        div_ash_111_n681), .A4(div_ash_111_n848), .Y(div_ash_111_n780) );
  AND2X1_LVT div_ash_111_U773 ( .A1(div_ash_111_n680), .A2(div_ash_111_n780), 
        .Y(div_n_T_442[23]) );
  AO22X1_LVT div_ash_111_U772 ( .A1(div_n168), .A2(div_ash_111_n846), .A3(
        div_ash_111_n682), .A4(div_ash_111_n845), .Y(div_ash_111_n925) );
  AO22X1_LVT div_ash_111_U771 ( .A1(div_n171), .A2(div_n_T_51_23_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_24_), .Y(div_ash_111_n918) );
  AO22X1_LVT div_ash_111_U770 ( .A1(div_n166), .A2(div_ash_111_n928), .A3(
        div_ash_111_n684), .A4(div_ash_111_n918), .Y(div_ash_111_n905) );
  AO22X1_LVT div_ash_111_U769 ( .A1(div_n167), .A2(div_ash_111_n927), .A3(
        div_ash_111_n683), .A4(div_ash_111_n905), .Y(div_ash_111_n887) );
  AO22X1_LVT div_ash_111_U768 ( .A1(div_n168), .A2(div_ash_111_n926), .A3(
        div_ash_111_n682), .A4(div_ash_111_n887), .Y(div_ash_111_n841) );
  AO22X1_LVT div_ash_111_U767 ( .A1(div_n169), .A2(div_ash_111_n925), .A3(
        div_ash_111_n681), .A4(div_ash_111_n841), .Y(div_ash_111_n777) );
  AO22X1_LVT div_ash_111_U766 ( .A1(div_n168), .A2(div_ash_111_n840), .A3(
        div_ash_111_n682), .A4(div_ash_111_n839), .Y(div_ash_111_n921) );
  AO22X1_LVT div_ash_111_U765 ( .A1(div_n171), .A2(div_n_T_51_24_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_25_), .Y(div_ash_111_n912) );
  AO22X1_LVT div_ash_111_U764 ( .A1(div_n166), .A2(div_ash_111_n924), .A3(
        div_ash_111_n684), .A4(div_ash_111_n912), .Y(div_ash_111_n901) );
  AO22X1_LVT div_ash_111_U763 ( .A1(div_n167), .A2(div_ash_111_n923), .A3(
        div_ash_111_n683), .A4(div_ash_111_n901), .Y(div_ash_111_n882) );
  AO22X1_LVT div_ash_111_U762 ( .A1(div_n168), .A2(div_ash_111_n922), .A3(
        div_ash_111_n682), .A4(div_ash_111_n882), .Y(div_ash_111_n835) );
  AO22X1_LVT div_ash_111_U761 ( .A1(div_n169), .A2(div_ash_111_n921), .A3(
        div_ash_111_n681), .A4(div_ash_111_n835), .Y(div_ash_111_n774) );
  AND2X1_LVT div_ash_111_U760 ( .A1(div_ash_111_n680), .A2(div_ash_111_n774), 
        .Y(div_n_T_442[25]) );
  AO22X1_LVT div_ash_111_U759 ( .A1(div_n168), .A2(div_ash_111_n919), .A3(
        div_ash_111_n682), .A4(div_ash_111_n920), .Y(div_ash_111_n915) );
  AO22X1_LVT div_ash_111_U758 ( .A1(div_n171), .A2(div_n_T_51_25_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_26_), .Y(div_ash_111_n906) );
  AO22X1_LVT div_ash_111_U757 ( .A1(div_n166), .A2(div_ash_111_n918), .A3(
        div_ash_111_n684), .A4(div_ash_111_n906), .Y(div_ash_111_n896) );
  AO22X1_LVT div_ash_111_U756 ( .A1(div_n167), .A2(div_ash_111_n917), .A3(
        div_ash_111_n683), .A4(div_ash_111_n896), .Y(div_ash_111_n877) );
  AO22X1_LVT div_ash_111_U755 ( .A1(div_n168), .A2(div_ash_111_n916), .A3(
        div_ash_111_n682), .A4(div_ash_111_n877), .Y(div_ash_111_n831) );
  AO22X1_LVT div_ash_111_U754 ( .A1(div_n169), .A2(div_ash_111_n915), .A3(
        div_ash_111_n681), .A4(div_ash_111_n831), .Y(div_ash_111_n771) );
  AND2X1_LVT div_ash_111_U753 ( .A1(div_ash_111_n680), .A2(div_ash_111_n771), 
        .Y(div_n_T_442[26]) );
  AO22X1_LVT div_ash_111_U752 ( .A1(div_n168), .A2(div_ash_111_n913), .A3(
        div_ash_111_n682), .A4(div_ash_111_n914), .Y(div_ash_111_n909) );
  AO22X1_LVT div_ash_111_U751 ( .A1(div_n171), .A2(div_n_T_51_26_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_27_), .Y(div_ash_111_n902) );
  AO22X1_LVT div_ash_111_U750 ( .A1(div_n166), .A2(div_ash_111_n912), .A3(
        div_ash_111_n684), .A4(div_ash_111_n902), .Y(div_ash_111_n892) );
  AO22X1_LVT div_ash_111_U749 ( .A1(div_n167), .A2(div_ash_111_n911), .A3(
        div_ash_111_n683), .A4(div_ash_111_n892), .Y(div_ash_111_n871) );
  AO22X1_LVT div_ash_111_U748 ( .A1(div_n168), .A2(div_ash_111_n910), .A3(
        div_ash_111_n682), .A4(div_ash_111_n871), .Y(div_ash_111_n826) );
  AO22X1_LVT div_ash_111_U747 ( .A1(div_n169), .A2(div_ash_111_n909), .A3(
        div_ash_111_n681), .A4(div_ash_111_n826), .Y(div_ash_111_n768) );
  AND2X1_LVT div_ash_111_U746 ( .A1(div_ash_111_n680), .A2(div_ash_111_n768), 
        .Y(div_n_T_442[27]) );
  AO22X1_LVT div_ash_111_U745 ( .A1(div_n168), .A2(div_ash_111_n907), .A3(
        div_ash_111_n682), .A4(div_ash_111_n908), .Y(div_ash_111_n903) );
  AO22X1_LVT div_ash_111_U744 ( .A1(div_n171), .A2(div_n_T_51_27_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_28_), .Y(div_ash_111_n897) );
  AO22X1_LVT div_ash_111_U743 ( .A1(div_n166), .A2(div_ash_111_n906), .A3(
        div_ash_111_n684), .A4(div_ash_111_n897), .Y(div_ash_111_n888) );
  AO22X1_LVT div_ash_111_U742 ( .A1(div_n167), .A2(div_ash_111_n905), .A3(
        div_ash_111_n683), .A4(div_ash_111_n888), .Y(div_ash_111_n866) );
  AO22X1_LVT div_ash_111_U741 ( .A1(div_n168), .A2(div_ash_111_n904), .A3(
        div_ash_111_n682), .A4(div_ash_111_n866), .Y(div_ash_111_n822) );
  AO22X1_LVT div_ash_111_U740 ( .A1(div_n169), .A2(div_ash_111_n903), .A3(
        div_ash_111_n681), .A4(div_ash_111_n822), .Y(div_ash_111_n764) );
  AND2X1_LVT div_ash_111_U739 ( .A1(div_ash_111_n680), .A2(div_ash_111_n764), 
        .Y(div_n_T_442[28]) );
  AO22X1_LVT div_ash_111_U738 ( .A1(div_n171), .A2(div_n_T_51_28_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_29_), .Y(div_ash_111_n893) );
  AO22X1_LVT div_ash_111_U737 ( .A1(div_n166), .A2(div_ash_111_n902), .A3(
        div_ash_111_n684), .A4(div_ash_111_n893), .Y(div_ash_111_n883) );
  AO22X1_LVT div_ash_111_U736 ( .A1(div_n167), .A2(div_ash_111_n901), .A3(
        div_ash_111_n683), .A4(div_ash_111_n883), .Y(div_ash_111_n861) );
  AO22X1_LVT div_ash_111_U735 ( .A1(div_n168), .A2(div_ash_111_n900), .A3(
        div_ash_111_n682), .A4(div_ash_111_n861), .Y(div_ash_111_n818) );
  AO22X1_LVT div_ash_111_U734 ( .A1(div_n169), .A2(div_ash_111_n899), .A3(
        div_ash_111_n681), .A4(div_ash_111_n818), .Y(div_ash_111_n761) );
  AND2X1_LVT div_ash_111_U733 ( .A1(div_ash_111_n680), .A2(div_ash_111_n761), 
        .Y(div_n_T_442[29]) );
  AND2X1_LVT div_ash_111_U732 ( .A1(div_ash_111_n898), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n875) );
  AO22X1_LVT div_ash_111_U731 ( .A1(div_n171), .A2(div_n_T_51_29_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_30_), .Y(div_ash_111_n889) );
  AO22X1_LVT div_ash_111_U730 ( .A1(div_n166), .A2(div_ash_111_n897), .A3(
        div_ash_111_n684), .A4(div_ash_111_n889), .Y(div_ash_111_n878) );
  AO22X1_LVT div_ash_111_U729 ( .A1(div_n167), .A2(div_ash_111_n896), .A3(
        div_ash_111_n683), .A4(div_ash_111_n878), .Y(div_ash_111_n855) );
  AO22X1_LVT div_ash_111_U728 ( .A1(div_n168), .A2(div_ash_111_n895), .A3(
        div_ash_111_n682), .A4(div_ash_111_n855), .Y(div_ash_111_n814) );
  AO22X1_LVT div_ash_111_U727 ( .A1(div_n169), .A2(div_ash_111_n894), .A3(
        div_ash_111_n681), .A4(div_ash_111_n814), .Y(div_ash_111_n758) );
  AND2X1_LVT div_ash_111_U726 ( .A1(div_ash_111_n680), .A2(div_ash_111_n758), 
        .Y(div_n_T_442[30]) );
  AO22X1_LVT div_ash_111_U725 ( .A1(div_n171), .A2(div_n_T_51_30_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_31_), .Y(div_ash_111_n884) );
  AO22X1_LVT div_ash_111_U724 ( .A1(div_n166), .A2(div_ash_111_n893), .A3(
        div_ash_111_n684), .A4(div_ash_111_n884), .Y(div_ash_111_n872) );
  AO22X1_LVT div_ash_111_U723 ( .A1(div_n167), .A2(div_ash_111_n892), .A3(
        div_ash_111_n683), .A4(div_ash_111_n872), .Y(div_ash_111_n849) );
  AO22X1_LVT div_ash_111_U722 ( .A1(div_n168), .A2(div_ash_111_n891), .A3(
        div_ash_111_n682), .A4(div_ash_111_n849), .Y(div_ash_111_n810) );
  AO22X1_LVT div_ash_111_U721 ( .A1(div_n169), .A2(div_ash_111_n890), .A3(
        div_ash_111_n681), .A4(div_ash_111_n810), .Y(div_ash_111_n756) );
  AND2X1_LVT div_ash_111_U720 ( .A1(div_ash_111_n680), .A2(div_ash_111_n756), 
        .Y(div_n_T_442[31]) );
  AO22X1_LVT div_ash_111_U719 ( .A1(div_n171), .A2(div_n_T_51_31_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_32_), .Y(div_ash_111_n879) );
  AO22X1_LVT div_ash_111_U718 ( .A1(div_n166), .A2(div_ash_111_n889), .A3(
        div_ash_111_n684), .A4(div_ash_111_n879), .Y(div_ash_111_n867) );
  AO22X1_LVT div_ash_111_U717 ( .A1(div_n167), .A2(div_ash_111_n888), .A3(
        div_ash_111_n683), .A4(div_ash_111_n867), .Y(div_ash_111_n842) );
  AO22X1_LVT div_ash_111_U716 ( .A1(div_n168), .A2(div_ash_111_n887), .A3(
        div_ash_111_n682), .A4(div_ash_111_n842), .Y(div_ash_111_n806) );
  AO22X1_LVT div_ash_111_U715 ( .A1(div_n169), .A2(div_ash_111_n886), .A3(
        div_ash_111_n681), .A4(div_ash_111_n806), .Y(div_ash_111_n754) );
  AO22X1_LVT div_ash_111_U714 ( .A1(div_n171), .A2(div_n_T_51_32_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_33_), .Y(div_ash_111_n873) );
  AO22X1_LVT div_ash_111_U713 ( .A1(div_n166), .A2(div_ash_111_n884), .A3(
        div_ash_111_n684), .A4(div_ash_111_n873), .Y(div_ash_111_n862) );
  AO22X1_LVT div_ash_111_U712 ( .A1(div_n167), .A2(div_ash_111_n883), .A3(
        div_ash_111_n683), .A4(div_ash_111_n862), .Y(div_ash_111_n836) );
  AO22X1_LVT div_ash_111_U711 ( .A1(div_n168), .A2(div_ash_111_n882), .A3(
        div_ash_111_n682), .A4(div_ash_111_n836), .Y(div_ash_111_n802) );
  AO22X1_LVT div_ash_111_U710 ( .A1(div_n169), .A2(div_ash_111_n881), .A3(
        div_ash_111_n681), .A4(div_ash_111_n802), .Y(div_ash_111_n752) );
  AO22X1_LVT div_ash_111_U709 ( .A1(div_n170), .A2(div_ash_111_n880), .A3(
        div_ash_111_n680), .A4(div_ash_111_n752), .Y(div_n_T_442[33]) );
  AO22X1_LVT div_ash_111_U708 ( .A1(div_n171), .A2(div_n_T_51_33_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_34_), .Y(div_ash_111_n868) );
  AO22X1_LVT div_ash_111_U707 ( .A1(div_n166), .A2(div_ash_111_n879), .A3(
        div_ash_111_n684), .A4(div_ash_111_n868), .Y(div_ash_111_n856) );
  AO22X1_LVT div_ash_111_U706 ( .A1(div_n167), .A2(div_ash_111_n878), .A3(
        div_ash_111_n683), .A4(div_ash_111_n856), .Y(div_ash_111_n832) );
  AO22X1_LVT div_ash_111_U705 ( .A1(div_n168), .A2(div_ash_111_n877), .A3(
        div_ash_111_n682), .A4(div_ash_111_n832), .Y(div_ash_111_n797) );
  AO22X1_LVT div_ash_111_U704 ( .A1(div_n169), .A2(div_ash_111_n876), .A3(
        div_ash_111_n681), .A4(div_ash_111_n797), .Y(div_ash_111_n750) );
  AO22X1_LVT div_ash_111_U703 ( .A1(div_n170), .A2(div_ash_111_n875), .A3(
        div_ash_111_n680), .A4(div_ash_111_n750), .Y(div_n_T_442[34]) );
  AND2X1_LVT div_ash_111_U702 ( .A1(div_ash_111_n874), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n847) );
  AO22X1_LVT div_ash_111_U701 ( .A1(div_n171), .A2(div_n_T_51_34_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_35_), .Y(div_ash_111_n863) );
  AO22X1_LVT div_ash_111_U700 ( .A1(div_n166), .A2(div_ash_111_n873), .A3(
        div_ash_111_n684), .A4(div_ash_111_n863), .Y(div_ash_111_n850) );
  AO22X1_LVT div_ash_111_U699 ( .A1(div_n167), .A2(div_ash_111_n872), .A3(
        div_ash_111_n683), .A4(div_ash_111_n850), .Y(div_ash_111_n827) );
  AO22X1_LVT div_ash_111_U698 ( .A1(div_n168), .A2(div_ash_111_n871), .A3(
        div_ash_111_n682), .A4(div_ash_111_n827), .Y(div_ash_111_n793) );
  AO22X1_LVT div_ash_111_U697 ( .A1(div_n169), .A2(div_ash_111_n870), .A3(
        div_ash_111_n681), .A4(div_ash_111_n793), .Y(div_ash_111_n748) );
  AO22X1_LVT div_ash_111_U696 ( .A1(div_n170), .A2(div_ash_111_n847), .A3(
        div_ash_111_n680), .A4(div_ash_111_n748), .Y(div_n_T_442[35]) );
  AND2X1_LVT div_ash_111_U695 ( .A1(div_ash_111_n869), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n800) );
  AO22X1_LVT div_ash_111_U694 ( .A1(div_n171), .A2(div_n_T_51_35_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_36_), .Y(div_ash_111_n857) );
  AO22X1_LVT div_ash_111_U693 ( .A1(div_n166), .A2(div_ash_111_n868), .A3(
        div_ash_111_n684), .A4(div_ash_111_n857), .Y(div_ash_111_n843) );
  AO22X1_LVT div_ash_111_U692 ( .A1(div_n167), .A2(div_ash_111_n867), .A3(
        div_ash_111_n683), .A4(div_ash_111_n843), .Y(div_ash_111_n823) );
  AO22X1_LVT div_ash_111_U691 ( .A1(div_n168), .A2(div_ash_111_n866), .A3(
        div_ash_111_n682), .A4(div_ash_111_n823), .Y(div_ash_111_n790) );
  AO22X1_LVT div_ash_111_U690 ( .A1(div_n169), .A2(div_ash_111_n865), .A3(
        div_ash_111_n681), .A4(div_ash_111_n790), .Y(div_ash_111_n746) );
  AO22X1_LVT div_ash_111_U689 ( .A1(div_n170), .A2(div_ash_111_n800), .A3(
        div_ash_111_n680), .A4(div_ash_111_n746), .Y(div_n_T_442[36]) );
  AND2X1_LVT div_ash_111_U688 ( .A1(div_ash_111_n864), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n767) );
  AO22X1_LVT div_ash_111_U687 ( .A1(div_n171), .A2(div_n_T_51_36_), .A3(
        div_ash_111_n679), .A4(div_n_T_51_37_), .Y(div_ash_111_n851) );
  AO22X1_LVT div_ash_111_U686 ( .A1(div_n166), .A2(div_ash_111_n863), .A3(
        div_ash_111_n684), .A4(div_ash_111_n851), .Y(div_ash_111_n837) );
  AO22X1_LVT div_ash_111_U685 ( .A1(div_n167), .A2(div_ash_111_n862), .A3(
        div_ash_111_n683), .A4(div_ash_111_n837), .Y(div_ash_111_n819) );
  AO22X1_LVT div_ash_111_U684 ( .A1(div_n168), .A2(div_ash_111_n861), .A3(
        div_ash_111_n682), .A4(div_ash_111_n819), .Y(div_ash_111_n787) );
  AO22X1_LVT div_ash_111_U683 ( .A1(div_n169), .A2(div_ash_111_n860), .A3(
        div_ash_111_n681), .A4(div_ash_111_n787), .Y(div_ash_111_n744) );
  AO22X1_LVT div_ash_111_U682 ( .A1(div_n170), .A2(div_ash_111_n767), .A3(
        div_ash_111_n680), .A4(div_ash_111_n744), .Y(div_n_T_442[37]) );
  AND2X1_LVT div_ash_111_U681 ( .A1(div_ash_111_n859), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n743) );
  AO22X1_LVT div_ash_111_U680 ( .A1(div_n166), .A2(div_ash_111_n857), .A3(
        div_ash_111_n684), .A4(div_ash_111_n858), .Y(div_ash_111_n833) );
  AO22X1_LVT div_ash_111_U679 ( .A1(div_n167), .A2(div_ash_111_n856), .A3(
        div_ash_111_n683), .A4(div_ash_111_n833), .Y(div_ash_111_n815) );
  AO22X1_LVT div_ash_111_U678 ( .A1(div_n168), .A2(div_ash_111_n855), .A3(
        div_ash_111_n682), .A4(div_ash_111_n815), .Y(div_ash_111_n784) );
  AO22X1_LVT div_ash_111_U677 ( .A1(div_n169), .A2(div_ash_111_n854), .A3(
        div_ash_111_n681), .A4(div_ash_111_n784), .Y(div_ash_111_n741) );
  AO22X1_LVT div_ash_111_U676 ( .A1(div_n170), .A2(div_ash_111_n743), .A3(
        div_ash_111_n680), .A4(div_ash_111_n741), .Y(div_n_T_442[38]) );
  AND2X1_LVT div_ash_111_U675 ( .A1(div_ash_111_n853), .A2(div_ash_111_n681), 
        .Y(div_ash_111_n722) );
  AO22X1_LVT div_ash_111_U674 ( .A1(div_n166), .A2(div_ash_111_n851), .A3(
        div_ash_111_n684), .A4(div_ash_111_n852), .Y(div_ash_111_n828) );
  AO22X1_LVT div_ash_111_U673 ( .A1(div_n167), .A2(div_ash_111_n850), .A3(
        div_ash_111_n683), .A4(div_ash_111_n828), .Y(div_ash_111_n811) );
  AO22X1_LVT div_ash_111_U672 ( .A1(div_n168), .A2(div_ash_111_n849), .A3(
        div_ash_111_n682), .A4(div_ash_111_n811), .Y(div_ash_111_n781) );
  AO22X1_LVT div_ash_111_U671 ( .A1(div_n169), .A2(div_ash_111_n848), .A3(
        div_ash_111_n681), .A4(div_ash_111_n781), .Y(div_ash_111_n739) );
  AO22X1_LVT div_ash_111_U670 ( .A1(div_n170), .A2(div_ash_111_n722), .A3(
        div_ash_111_n680), .A4(div_ash_111_n739), .Y(div_n_T_442[39]) );
  AND2X1_LVT div_ash_111_U669 ( .A1(div_ash_111_n847), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[3]) );
  OA221X1_LVT div_ash_111_U668 ( .A1(div_n168), .A2(div_ash_111_n845), .A3(
        div_ash_111_n682), .A4(div_ash_111_n846), .A5(div_ash_111_n681), .Y(
        div_ash_111_n701) );
  AO22X1_LVT div_ash_111_U667 ( .A1(div_n167), .A2(div_ash_111_n843), .A3(
        div_ash_111_n683), .A4(div_ash_111_n844), .Y(div_ash_111_n807) );
  AO22X1_LVT div_ash_111_U666 ( .A1(div_n168), .A2(div_ash_111_n842), .A3(
        div_ash_111_n682), .A4(div_ash_111_n807), .Y(div_ash_111_n778) );
  AO22X1_LVT div_ash_111_U665 ( .A1(div_n169), .A2(div_ash_111_n841), .A3(
        div_ash_111_n681), .A4(div_ash_111_n778), .Y(div_ash_111_n737) );
  OA221X1_LVT div_ash_111_U664 ( .A1(div_n168), .A2(div_ash_111_n839), .A3(
        div_ash_111_n682), .A4(div_ash_111_n840), .A5(div_ash_111_n681), .Y(
        div_ash_111_n685) );
  AO22X1_LVT div_ash_111_U663 ( .A1(div_n167), .A2(div_ash_111_n837), .A3(
        div_ash_111_n683), .A4(div_ash_111_n838), .Y(div_ash_111_n803) );
  AO22X1_LVT div_ash_111_U662 ( .A1(div_n168), .A2(div_ash_111_n836), .A3(
        div_ash_111_n682), .A4(div_ash_111_n803), .Y(div_ash_111_n775) );
  AO22X1_LVT div_ash_111_U661 ( .A1(div_n169), .A2(div_ash_111_n835), .A3(
        div_ash_111_n681), .A4(div_ash_111_n775), .Y(div_ash_111_n735) );
  AO22X1_LVT div_ash_111_U660 ( .A1(div_n170), .A2(div_ash_111_n685), .A3(
        div_ash_111_n680), .A4(div_ash_111_n735), .Y(div_n_T_442[41]) );
  AO22X1_LVT div_ash_111_U659 ( .A1(div_n167), .A2(div_ash_111_n833), .A3(
        div_ash_111_n683), .A4(div_ash_111_n834), .Y(div_ash_111_n798) );
  AO22X1_LVT div_ash_111_U658 ( .A1(div_n168), .A2(div_ash_111_n832), .A3(
        div_ash_111_n682), .A4(div_ash_111_n798), .Y(div_ash_111_n772) );
  AO22X1_LVT div_ash_111_U657 ( .A1(div_n169), .A2(div_ash_111_n831), .A3(
        div_ash_111_n681), .A4(div_ash_111_n772), .Y(div_ash_111_n733) );
  AO22X1_LVT div_ash_111_U656 ( .A1(div_n170), .A2(div_ash_111_n830), .A3(
        div_ash_111_n680), .A4(div_ash_111_n733), .Y(div_n_T_442[42]) );
  AO22X1_LVT div_ash_111_U655 ( .A1(div_n167), .A2(div_ash_111_n828), .A3(
        div_ash_111_n683), .A4(div_ash_111_n829), .Y(div_ash_111_n794) );
  AO22X1_LVT div_ash_111_U654 ( .A1(div_n168), .A2(div_ash_111_n827), .A3(
        div_ash_111_n682), .A4(div_ash_111_n794), .Y(div_ash_111_n769) );
  AO22X1_LVT div_ash_111_U653 ( .A1(div_n169), .A2(div_ash_111_n826), .A3(
        div_ash_111_n681), .A4(div_ash_111_n769), .Y(div_ash_111_n731) );
  AO22X1_LVT div_ash_111_U652 ( .A1(div_n170), .A2(div_ash_111_n825), .A3(
        div_ash_111_n680), .A4(div_ash_111_n731), .Y(div_n_T_442[43]) );
  AO22X1_LVT div_ash_111_U651 ( .A1(div_n168), .A2(div_ash_111_n823), .A3(
        div_ash_111_n682), .A4(div_ash_111_n824), .Y(div_ash_111_n765) );
  AO22X1_LVT div_ash_111_U650 ( .A1(div_n169), .A2(div_ash_111_n822), .A3(
        div_ash_111_n681), .A4(div_ash_111_n765), .Y(div_ash_111_n729) );
  AO22X1_LVT div_ash_111_U649 ( .A1(div_n170), .A2(div_ash_111_n821), .A3(
        div_ash_111_n680), .A4(div_ash_111_n729), .Y(div_n_T_442[44]) );
  AO22X1_LVT div_ash_111_U648 ( .A1(div_n168), .A2(div_ash_111_n819), .A3(
        div_ash_111_n682), .A4(div_ash_111_n820), .Y(div_ash_111_n762) );
  AO22X1_LVT div_ash_111_U647 ( .A1(div_n169), .A2(div_ash_111_n818), .A3(
        div_ash_111_n681), .A4(div_ash_111_n762), .Y(div_ash_111_n727) );
  AO22X1_LVT div_ash_111_U646 ( .A1(div_n170), .A2(div_ash_111_n817), .A3(
        div_ash_111_n680), .A4(div_ash_111_n727), .Y(div_n_T_442[45]) );
  AO22X1_LVT div_ash_111_U645 ( .A1(div_n168), .A2(div_ash_111_n815), .A3(
        div_ash_111_n682), .A4(div_ash_111_n816), .Y(div_ash_111_n759) );
  AO22X1_LVT div_ash_111_U644 ( .A1(div_n169), .A2(div_ash_111_n814), .A3(
        div_ash_111_n681), .A4(div_ash_111_n759), .Y(div_ash_111_n725) );
  AO22X1_LVT div_ash_111_U643 ( .A1(div_n170), .A2(div_ash_111_n813), .A3(
        div_ash_111_n680), .A4(div_ash_111_n725), .Y(div_n_T_442[46]) );
  AO22X1_LVT div_ash_111_U642 ( .A1(div_n168), .A2(div_ash_111_n811), .A3(
        div_ash_111_n682), .A4(div_ash_111_n812), .Y(div_ash_111_n757) );
  AO22X1_LVT div_ash_111_U641 ( .A1(div_n169), .A2(div_ash_111_n810), .A3(
        div_ash_111_n681), .A4(div_ash_111_n757), .Y(div_ash_111_n724) );
  AO22X1_LVT div_ash_111_U640 ( .A1(div_n170), .A2(div_ash_111_n809), .A3(
        div_ash_111_n680), .A4(div_ash_111_n724), .Y(div_n_T_442[47]) );
  AO22X1_LVT div_ash_111_U639 ( .A1(div_n168), .A2(div_ash_111_n807), .A3(
        div_ash_111_n682), .A4(div_ash_111_n808), .Y(div_ash_111_n755) );
  AO22X1_LVT div_ash_111_U638 ( .A1(div_n169), .A2(div_ash_111_n806), .A3(
        div_ash_111_n681), .A4(div_ash_111_n755), .Y(div_ash_111_n721) );
  AO22X1_LVT div_ash_111_U637 ( .A1(div_n168), .A2(div_ash_111_n803), .A3(
        div_ash_111_n682), .A4(div_ash_111_n804), .Y(div_ash_111_n753) );
  AO22X1_LVT div_ash_111_U636 ( .A1(div_n169), .A2(div_ash_111_n802), .A3(
        div_ash_111_n681), .A4(div_ash_111_n753), .Y(div_ash_111_n719) );
  AO22X1_LVT div_ash_111_U635 ( .A1(div_n170), .A2(div_ash_111_n801), .A3(
        div_ash_111_n680), .A4(div_ash_111_n719), .Y(div_n_T_442[49]) );
  AO22X1_LVT div_ash_111_U634 ( .A1(div_n168), .A2(div_ash_111_n798), .A3(
        div_ash_111_n682), .A4(div_ash_111_n799), .Y(div_ash_111_n751) );
  AO22X1_LVT div_ash_111_U633 ( .A1(div_n169), .A2(div_ash_111_n797), .A3(
        div_ash_111_n681), .A4(div_ash_111_n751), .Y(div_ash_111_n717) );
  AO22X1_LVT div_ash_111_U632 ( .A1(div_n170), .A2(div_ash_111_n796), .A3(
        div_ash_111_n680), .A4(div_ash_111_n717), .Y(div_n_T_442[50]) );
  AO22X1_LVT div_ash_111_U631 ( .A1(div_n168), .A2(div_ash_111_n794), .A3(
        div_ash_111_n682), .A4(div_ash_111_n795), .Y(div_ash_111_n749) );
  AO22X1_LVT div_ash_111_U630 ( .A1(div_n169), .A2(div_ash_111_n793), .A3(
        div_ash_111_n681), .A4(div_ash_111_n749), .Y(div_ash_111_n715) );
  AO22X1_LVT div_ash_111_U629 ( .A1(div_n170), .A2(div_ash_111_n792), .A3(
        div_ash_111_n680), .A4(div_ash_111_n715), .Y(div_n_T_442[51]) );
  AO22X1_LVT div_ash_111_U628 ( .A1(div_n169), .A2(div_ash_111_n790), .A3(
        div_ash_111_n681), .A4(div_ash_111_n791), .Y(div_ash_111_n713) );
  AO22X1_LVT div_ash_111_U627 ( .A1(div_n169), .A2(div_ash_111_n787), .A3(
        div_ash_111_n681), .A4(div_ash_111_n788), .Y(div_ash_111_n711) );
  AO22X1_LVT div_ash_111_U626 ( .A1(div_n170), .A2(div_ash_111_n786), .A3(
        div_ash_111_n680), .A4(div_ash_111_n711), .Y(div_n_T_442[53]) );
  AO22X1_LVT div_ash_111_U625 ( .A1(div_n169), .A2(div_ash_111_n784), .A3(
        div_ash_111_n681), .A4(div_ash_111_n785), .Y(div_ash_111_n709) );
  AO22X1_LVT div_ash_111_U624 ( .A1(div_n170), .A2(div_ash_111_n783), .A3(
        div_ash_111_n680), .A4(div_ash_111_n709), .Y(div_n_T_442[54]) );
  AO22X1_LVT div_ash_111_U623 ( .A1(div_n169), .A2(div_ash_111_n781), .A3(
        div_ash_111_n681), .A4(div_ash_111_n782), .Y(div_ash_111_n706) );
  AO22X1_LVT div_ash_111_U622 ( .A1(div_n170), .A2(div_ash_111_n780), .A3(
        div_ash_111_n680), .A4(div_ash_111_n706), .Y(div_n_T_442[55]) );
  AO22X1_LVT div_ash_111_U621 ( .A1(div_n169), .A2(div_ash_111_n778), .A3(
        div_ash_111_n681), .A4(div_ash_111_n779), .Y(div_ash_111_n704) );
  AO22X1_LVT div_ash_111_U620 ( .A1(div_n169), .A2(div_ash_111_n775), .A3(
        div_ash_111_n681), .A4(div_ash_111_n776), .Y(div_ash_111_n702) );
  AO22X1_LVT div_ash_111_U619 ( .A1(div_n170), .A2(div_ash_111_n774), .A3(
        div_ash_111_n680), .A4(div_ash_111_n702), .Y(div_n_T_442[57]) );
  AO22X1_LVT div_ash_111_U618 ( .A1(div_n169), .A2(div_ash_111_n772), .A3(
        div_ash_111_n681), .A4(div_ash_111_n773), .Y(div_ash_111_n699) );
  AO22X1_LVT div_ash_111_U617 ( .A1(div_n170), .A2(div_ash_111_n771), .A3(
        div_ash_111_n680), .A4(div_ash_111_n699), .Y(div_n_T_442[58]) );
  AO22X1_LVT div_ash_111_U616 ( .A1(div_n169), .A2(div_ash_111_n769), .A3(
        div_ash_111_n681), .A4(div_ash_111_n770), .Y(div_ash_111_n698) );
  AO22X1_LVT div_ash_111_U615 ( .A1(div_n170), .A2(div_ash_111_n768), .A3(
        div_ash_111_n680), .A4(div_ash_111_n698), .Y(div_n_T_442[59]) );
  AND2X1_LVT div_ash_111_U614 ( .A1(div_ash_111_n767), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[5]) );
  AO22X1_LVT div_ash_111_U613 ( .A1(div_n169), .A2(div_ash_111_n765), .A3(
        div_ash_111_n681), .A4(div_ash_111_n766), .Y(div_ash_111_n696) );
  AO22X1_LVT div_ash_111_U612 ( .A1(div_n170), .A2(div_ash_111_n764), .A3(
        div_ash_111_n680), .A4(div_ash_111_n696), .Y(div_n_T_442[60]) );
  AO22X1_LVT div_ash_111_U611 ( .A1(div_n169), .A2(div_ash_111_n762), .A3(
        div_ash_111_n681), .A4(div_ash_111_n763), .Y(div_ash_111_n693) );
  AO22X1_LVT div_ash_111_U610 ( .A1(div_n170), .A2(div_ash_111_n761), .A3(
        div_ash_111_n680), .A4(div_ash_111_n693), .Y(div_n_T_442[61]) );
  AO22X1_LVT div_ash_111_U609 ( .A1(div_n169), .A2(div_ash_111_n759), .A3(
        div_ash_111_n681), .A4(div_ash_111_n760), .Y(div_ash_111_n692) );
  AO22X1_LVT div_ash_111_U608 ( .A1(div_n170), .A2(div_ash_111_n758), .A3(
        div_ash_111_n680), .A4(div_ash_111_n692), .Y(div_n_T_442[62]) );
  AO22X1_LVT div_ash_111_U607 ( .A1(div_n169), .A2(div_ash_111_n757), .A3(
        div_ash_111_n681), .A4(div_ash_111_n723), .Y(div_ash_111_n690) );
  AO22X1_LVT div_ash_111_U606 ( .A1(div_n170), .A2(div_ash_111_n756), .A3(
        div_ash_111_n680), .A4(div_ash_111_n690), .Y(div_n_T_442[63]) );
  AO22X1_LVT div_ash_111_U605 ( .A1(div_n169), .A2(div_ash_111_n755), .A3(
        div_ash_111_n681), .A4(div_ash_111_n720), .Y(div_ash_111_n689) );
  AO22X1_LVT div_ash_111_U604 ( .A1(div_n169), .A2(div_ash_111_n753), .A3(
        div_ash_111_n681), .A4(div_ash_111_n718), .Y(div_ash_111_n688) );
  AO22X1_LVT div_ash_111_U603 ( .A1(div_n170), .A2(div_ash_111_n752), .A3(
        div_ash_111_n680), .A4(div_ash_111_n688), .Y(div_n_T_442[65]) );
  AO22X1_LVT div_ash_111_U602 ( .A1(div_n169), .A2(div_ash_111_n751), .A3(
        div_ash_111_n681), .A4(div_ash_111_n716), .Y(div_ash_111_n687) );
  AO22X1_LVT div_ash_111_U601 ( .A1(div_n170), .A2(div_ash_111_n750), .A3(
        div_ash_111_n680), .A4(div_ash_111_n687), .Y(div_n_T_442[66]) );
  AO22X1_LVT div_ash_111_U600 ( .A1(div_n169), .A2(div_ash_111_n749), .A3(
        div_ash_111_n681), .A4(div_ash_111_n714), .Y(div_ash_111_n686) );
  AO22X1_LVT div_ash_111_U599 ( .A1(div_n170), .A2(div_ash_111_n748), .A3(
        div_ash_111_n680), .A4(div_ash_111_n686), .Y(div_n_T_442[67]) );
  AO22X1_LVT div_ash_111_U598 ( .A1(div_n170), .A2(div_ash_111_n746), .A3(
        div_ash_111_n680), .A4(div_ash_111_n747), .Y(div_n_T_442[68]) );
  AO22X1_LVT div_ash_111_U597 ( .A1(div_n170), .A2(div_ash_111_n744), .A3(
        div_ash_111_n680), .A4(div_ash_111_n745), .Y(div_n_T_442[69]) );
  AND2X1_LVT div_ash_111_U596 ( .A1(div_ash_111_n743), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[6]) );
  AO22X1_LVT div_ash_111_U595 ( .A1(div_n170), .A2(div_ash_111_n741), .A3(
        div_ash_111_n680), .A4(div_ash_111_n742), .Y(div_n_T_442[70]) );
  AO22X1_LVT div_ash_111_U594 ( .A1(div_n170), .A2(div_ash_111_n739), .A3(
        div_ash_111_n680), .A4(div_ash_111_n740), .Y(div_n_T_442[71]) );
  AO22X1_LVT div_ash_111_U593 ( .A1(div_n170), .A2(div_ash_111_n737), .A3(
        div_ash_111_n680), .A4(div_ash_111_n738), .Y(div_n_T_442[72]) );
  AO22X1_LVT div_ash_111_U592 ( .A1(div_n170), .A2(div_ash_111_n735), .A3(
        div_ash_111_n680), .A4(div_ash_111_n736), .Y(div_n_T_442[73]) );
  AO22X1_LVT div_ash_111_U591 ( .A1(div_n170), .A2(div_ash_111_n733), .A3(
        div_ash_111_n680), .A4(div_ash_111_n734), .Y(div_n_T_442[74]) );
  AO22X1_LVT div_ash_111_U590 ( .A1(div_n170), .A2(div_ash_111_n731), .A3(
        div_ash_111_n680), .A4(div_ash_111_n732), .Y(div_n_T_442[75]) );
  AO22X1_LVT div_ash_111_U589 ( .A1(div_n170), .A2(div_ash_111_n729), .A3(
        div_ash_111_n680), .A4(div_ash_111_n730), .Y(div_n_T_442[76]) );
  AO22X1_LVT div_ash_111_U588 ( .A1(div_n170), .A2(div_ash_111_n727), .A3(
        div_ash_111_n680), .A4(div_ash_111_n728), .Y(div_n_T_442[77]) );
  AO22X1_LVT div_ash_111_U587 ( .A1(div_n170), .A2(div_ash_111_n725), .A3(
        div_ash_111_n680), .A4(div_ash_111_n726), .Y(div_n_T_442[78]) );
  OA222X1_LVT div_ash_111_U586 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n723), .A5(div_ash_111_n680), .A6(div_ash_111_n724), 
        .Y(div_n_T_442[79]) );
  AND2X1_LVT div_ash_111_U585 ( .A1(div_ash_111_n722), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[7]) );
  OA222X1_LVT div_ash_111_U584 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n720), .A5(div_ash_111_n680), .A6(div_ash_111_n721), 
        .Y(div_n_T_442[80]) );
  OA222X1_LVT div_ash_111_U583 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n718), .A5(div_ash_111_n680), .A6(div_ash_111_n719), 
        .Y(div_n_T_442[81]) );
  OA222X1_LVT div_ash_111_U582 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n716), .A5(div_ash_111_n680), .A6(div_ash_111_n717), 
        .Y(div_n_T_442[82]) );
  OA222X1_LVT div_ash_111_U581 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n714), .A5(div_ash_111_n680), .A6(div_ash_111_n715), 
        .Y(div_n_T_442[83]) );
  OA222X1_LVT div_ash_111_U580 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n712), .A5(div_ash_111_n680), .A6(div_ash_111_n713), 
        .Y(div_n_T_442[84]) );
  OA222X1_LVT div_ash_111_U579 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n710), .A5(div_ash_111_n680), .A6(div_ash_111_n711), 
        .Y(div_n_T_442[85]) );
  OA222X1_LVT div_ash_111_U578 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n708), .A5(div_ash_111_n680), .A6(div_ash_111_n709), 
        .Y(div_n_T_442[86]) );
  AO22X1_LVT div_ash_111_U577 ( .A1(div_n170), .A2(div_ash_111_n706), .A3(
        div_ash_111_n680), .A4(div_ash_111_n707), .Y(div_n_T_442[87]) );
  AO22X1_LVT div_ash_111_U576 ( .A1(div_n170), .A2(div_ash_111_n704), .A3(
        div_ash_111_n680), .A4(div_ash_111_n705), .Y(div_n_T_442[88]) );
  AO22X1_LVT div_ash_111_U575 ( .A1(div_n170), .A2(div_ash_111_n702), .A3(
        div_ash_111_n680), .A4(div_ash_111_n703), .Y(div_n_T_442[89]) );
  AND2X1_LVT div_ash_111_U574 ( .A1(div_ash_111_n701), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[8]) );
  AO22X1_LVT div_ash_111_U573 ( .A1(div_n170), .A2(div_ash_111_n699), .A3(
        div_ash_111_n680), .A4(div_ash_111_n700), .Y(div_n_T_442[90]) );
  OA222X1_LVT div_ash_111_U572 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n697), .A5(div_ash_111_n680), .A6(div_ash_111_n698), 
        .Y(div_n_T_442[91]) );
  OA222X1_LVT div_ash_111_U571 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n695), .A5(div_ash_111_n680), .A6(div_ash_111_n696), 
        .Y(div_n_T_442[92]) );
  AO22X1_LVT div_ash_111_U570 ( .A1(div_n170), .A2(div_ash_111_n693), .A3(
        div_ash_111_n680), .A4(div_ash_111_n694), .Y(div_n_T_442[93]) );
  OA222X1_LVT div_ash_111_U569 ( .A1(div_n170), .A2(div_n169), .A3(div_n170), 
        .A4(div_ash_111_n691), .A5(div_ash_111_n680), .A6(div_ash_111_n692), 
        .Y(div_n_T_442[94]) );
  AND2X1_LVT div_ash_111_U568 ( .A1(div_n170), .A2(div_ash_111_n690), .Y(
        div_n_T_442[95]) );
  AND2X1_LVT div_ash_111_U567 ( .A1(div_n170), .A2(div_ash_111_n689), .Y(
        div_n_T_442[96]) );
  AND2X1_LVT div_ash_111_U566 ( .A1(div_n170), .A2(div_ash_111_n688), .Y(
        div_n_T_442[97]) );
  AND2X1_LVT div_ash_111_U565 ( .A1(div_n170), .A2(div_ash_111_n687), .Y(
        div_n_T_442[98]) );
  AND2X1_LVT div_ash_111_U564 ( .A1(div_n170), .A2(div_ash_111_n686), .Y(
        div_n_T_442[99]) );
  AND2X1_LVT div_ash_111_U563 ( .A1(div_ash_111_n685), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[9]) );
  INVX1_LVT div_ash_111_U562 ( .A(div_n166), .Y(div_ash_111_n684) );
  INVX1_LVT div_ash_111_U561 ( .A(div_n171), .Y(div_ash_111_n679) );
  INVX1_LVT div_ash_111_U560 ( .A(div_n170), .Y(div_ash_111_n680) );
  INVX1_LVT div_ash_111_U559 ( .A(div_n169), .Y(div_ash_111_n681) );
  INVX1_LVT div_ash_111_U558 ( .A(div_n168), .Y(div_ash_111_n682) );
  INVX1_LVT div_ash_111_U557 ( .A(div_n167), .Y(div_ash_111_n683) );
  AO22X1_LVT div_ash_111_U556 ( .A1(div_n170), .A2(div_ash_111_n789), .A3(
        div_ash_111_n713), .A4(div_ash_111_n680), .Y(div_n_T_442[52]) );
  AO22X1_LVT div_ash_111_U555 ( .A1(div_n170), .A2(div_ash_111_n885), .A3(
        div_ash_111_n754), .A4(div_ash_111_n680), .Y(div_n_T_442[32]) );
  AND2X1_LVT div_ash_111_U554 ( .A1(div_ash_111_n680), .A2(div_ash_111_n880), 
        .Y(div_n_T_442[1]) );
  AND2X1_LVT div_ash_111_U553 ( .A1(div_ash_111_n885), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[0]) );
  AND2X1_LVT div_ash_111_U552 ( .A1(div_ash_111_n680), .A2(div_ash_111_n800), 
        .Y(div_n_T_442[4]) );
  AND2X1_LVT div_ash_111_U551 ( .A1(div_ash_111_n805), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[16]) );
  AND2X1_LVT div_ash_111_U550 ( .A1(div_ash_111_n680), .A2(div_ash_111_n875), 
        .Y(div_n_T_442[2]) );
  AND2X1_LVT div_ash_111_U549 ( .A1(div_ash_111_n777), .A2(div_ash_111_n680), 
        .Y(div_n_T_442[24]) );
  AO22X1_LVT div_ash_111_U548 ( .A1(div_n170), .A2(div_ash_111_n701), .A3(
        div_ash_111_n737), .A4(div_ash_111_n680), .Y(div_n_T_442[40]) );
  AO22X1_LVT div_ash_111_U547 ( .A1(div_n170), .A2(div_ash_111_n754), .A3(
        div_ash_111_n680), .A4(div_ash_111_n689), .Y(div_n_T_442[64]) );
  AND2X1_LVT div_ash_111_U546 ( .A1(div_ash_111_n680), .A2(div_ash_111_n821), 
        .Y(div_n_T_442[12]) );
  AO22X1_LVT div_ash_111_U545 ( .A1(div_n170), .A2(div_ash_111_n805), .A3(
        div_ash_111_n721), .A4(div_ash_111_n680), .Y(div_n_T_442[48]) );
  AO22X1_LVT div_ash_111_U544 ( .A1(div_n170), .A2(div_ash_111_n777), .A3(
        div_ash_111_n704), .A4(div_ash_111_n680), .Y(div_n_T_442[56]) );
  AO22X1_LVT div_sub_x_110_U76 ( .A1(div_n_T_429[0]), .A2(div_sub_x_110_n64), 
        .A3(div_sub_x_110_n66), .A4(div_n_T_272[0]), .Y(div_n_T_434_0_) );
  NAND2X0_LVT div_sub_x_110_U75 ( .A1(div_n_T_272[0]), .A2(div_sub_x_110_n66), 
        .Y(div_sub_x_110_n83) );
  FADDX1_LVT div_sub_x_110_U74 ( .A(div_n_T_272[1]), .B(div_sub_x_110_n67), 
        .CI(div_sub_x_110_n83), .S(div_n_T_434_1_) );
  NAND2X0_LVT div_sub_x_110_U73 ( .A1(div_n_T_272[1]), .A2(div_sub_x_110_n67), 
        .Y(div_sub_x_110_n81) );
  AO22X1_LVT div_sub_x_110_U72 ( .A1(div_n_T_429[1]), .A2(div_sub_x_110_n65), 
        .A3(div_sub_x_110_n83), .A4(div_sub_x_110_n81), .Y(div_sub_x_110_n85)
         );
  FADDX1_LVT div_sub_x_110_U71 ( .A(div_n_T_272[2]), .B(div_sub_x_110_n69), 
        .CI(div_sub_x_110_n85), .S(div_n_T_434_2_) );
  NAND2X0_LVT div_sub_x_110_U70 ( .A1(div_n_T_429[1]), .A2(div_sub_x_110_n65), 
        .Y(div_sub_x_110_n84) );
  AO222X1_LVT div_sub_x_110_U69 ( .A1(div_n_T_272[2]), .A2(div_sub_x_110_n69), 
        .A3(div_n_T_272[2]), .A4(div_sub_x_110_n84), .A5(div_sub_x_110_n69), 
        .A6(div_sub_x_110_n84), .Y(div_sub_x_110_n79) );
  NAND2X0_LVT div_sub_x_110_U68 ( .A1(div_n_T_272[2]), .A2(div_sub_x_110_n69), 
        .Y(div_sub_x_110_n82) );
  NAND3X0_LVT div_sub_x_110_U67 ( .A1(div_sub_x_110_n81), .A2(
        div_sub_x_110_n82), .A3(div_sub_x_110_n83), .Y(div_sub_x_110_n80) );
  AND2X1_LVT div_sub_x_110_U66 ( .A1(div_sub_x_110_n79), .A2(div_sub_x_110_n80), .Y(div_sub_x_110_n76) );
  FADDX1_LVT div_sub_x_110_U65 ( .A(div_n_T_429[3]), .B(div_n_T_272[3]), .CI(
        div_sub_x_110_n76), .S(div_n_T_434_3_) );
  AO22X1_LVT div_sub_x_110_U64 ( .A1(div_n_T_272[3]), .A2(div_sub_x_110_n68), 
        .A3(div_sub_x_110_n77), .A4(div_sub_x_110_n76), .Y(div_sub_x_110_n78)
         );
  FADDX1_LVT div_sub_x_110_U63 ( .A(div_n_T_429[4]), .B(div_n_T_272[4]), .CI(
        div_sub_x_110_n78), .S(div_n_T_434_4_) );
  AO222X1_LVT div_sub_x_110_U62 ( .A1(div_n_T_272[4]), .A2(div_sub_x_110_n77), 
        .A3(div_n_T_272[4]), .A4(div_sub_x_110_n70), .A5(div_sub_x_110_n77), 
        .A6(div_sub_x_110_n70), .Y(div_sub_x_110_n75) );
  NAND3X0_LVT div_sub_x_110_U61 ( .A1(div_n_T_272[4]), .A2(div_sub_x_110_n70), 
        .A3(div_sub_x_110_n75), .Y(div_sub_x_110_n72) );
  NAND2X0_LVT div_sub_x_110_U60 ( .A1(div_sub_x_110_n75), .A2(
        div_sub_x_110_n76), .Y(div_sub_x_110_n73) );
  NAND3X0_LVT div_sub_x_110_U59 ( .A1(div_n_T_272[3]), .A2(div_sub_x_110_n68), 
        .A3(div_sub_x_110_n75), .Y(div_sub_x_110_n74) );
  NAND3X0_LVT div_sub_x_110_U58 ( .A1(div_sub_x_110_n72), .A2(
        div_sub_x_110_n73), .A3(div_sub_x_110_n74), .Y(div_sub_x_110_n71) );
  INVX1_LVT div_sub_x_110_U57 ( .A(div_n_T_429[4]), .Y(div_sub_x_110_n70) );
  INVX1_LVT div_sub_x_110_U56 ( .A(div_n_T_272[1]), .Y(div_sub_x_110_n65) );
  INVX1_LVT div_sub_x_110_U55 ( .A(div_n_T_272[0]), .Y(div_sub_x_110_n64) );
  FADDX1_LVT div_sub_x_110_U54 ( .A(div_n_T_273_5_), .B(div_n_T_430_5_), .CI(
        div_sub_x_110_n71), .S(div_n_T_434_5_) );
  OR2X1_LVT div_sub_x_110_U53 ( .A1(div_sub_x_110_n68), .A2(div_n_T_272[3]), 
        .Y(div_sub_x_110_n77) );
  INVX0_LVT div_sub_x_110_U52 ( .A(div_n_T_429[3]), .Y(div_sub_x_110_n68) );
  INVX0_LVT div_sub_x_110_U51 ( .A(div_n_T_429[0]), .Y(div_sub_x_110_n66) );
  INVX0_LVT div_sub_x_110_U50 ( .A(div_n_T_429[1]), .Y(div_sub_x_110_n67) );
  INVX0_LVT div_sub_x_110_U49 ( .A(div_n_T_429[2]), .Y(div_sub_x_110_n69) );
  AO22X1_LVT div_ashr_12_U971 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_56_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_48_), .Y(div_ashr_12_n1033) );
  AO22X1_LVT div_ashr_12_U970 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_40_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_32_), .Y(div_ashr_12_n1031) );
  AO22X1_LVT div_ashr_12_U969 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1033), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1031), .Y(div_ashr_12_n991) );
  AO22X1_LVT div_ashr_12_U968 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_24_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_16_), .Y(div_ashr_12_n1032) );
  AO22X1_LVT div_ashr_12_U967 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_66_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_58_), .Y(div_ashr_12_n1019) );
  AO22X1_LVT div_ashr_12_U966 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_50_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_42_), .Y(div_ashr_12_n1017) );
  AO22X1_LVT div_ashr_12_U965 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1019), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1017), .Y(div_ashr_12_n952) );
  AO22X1_LVT div_ashr_12_U964 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_34_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_26_), .Y(div_ashr_12_n1018) );
  AO22X1_LVT div_ashr_12_U963 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_18_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_10_), .Y(div_ashr_12_n1043) );
  AO22X1_LVT div_ashr_12_U962 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1018), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1043), .Y(div_ashr_12_n1042)
         );
  AO22X1_LVT div_ashr_12_U961 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n952), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1042), .Y(div_n_T_87[10]) );
  AO22X1_LVT div_ashr_12_U960 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_67_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_59_), .Y(div_ashr_12_n1015) );
  AO22X1_LVT div_ashr_12_U959 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_51_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_43_), .Y(div_ashr_12_n1013) );
  AO22X1_LVT div_ashr_12_U958 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1015), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1013), .Y(div_ashr_12_n949) );
  AO22X1_LVT div_ashr_12_U957 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_35_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_27_), .Y(div_ashr_12_n1014) );
  AO22X1_LVT div_ashr_12_U956 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_19_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_11_), .Y(div_ashr_12_n1041) );
  AO22X1_LVT div_ashr_12_U955 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1014), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1041), .Y(div_ashr_12_n1040)
         );
  AO22X1_LVT div_ashr_12_U954 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n949), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1040), .Y(div_n_T_87[11]) );
  AO22X1_LVT div_ashr_12_U953 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_68_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_60_), .Y(div_ashr_12_n1011) );
  AO22X1_LVT div_ashr_12_U952 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_52_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_44_), .Y(div_ashr_12_n1009) );
  AO22X1_LVT div_ashr_12_U951 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1011), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1009), .Y(div_ashr_12_n946) );
  AO22X1_LVT div_ashr_12_U950 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_36_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_28_), .Y(div_ashr_12_n1010) );
  AO22X1_LVT div_ashr_12_U949 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_69_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_61_), .Y(div_ashr_12_n1007) );
  AO22X1_LVT div_ashr_12_U948 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_53_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_45_), .Y(div_ashr_12_n1005) );
  AO22X1_LVT div_ashr_12_U947 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1007), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1005), .Y(div_ashr_12_n943) );
  AO22X1_LVT div_ashr_12_U946 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_37_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_29_), .Y(div_ashr_12_n1006) );
  AO22X1_LVT div_ashr_12_U945 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_21_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_13_), .Y(div_ashr_12_n1039) );
  AO22X1_LVT div_ashr_12_U944 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1006), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1039), .Y(div_ashr_12_n1038)
         );
  AO22X1_LVT div_ashr_12_U943 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n943), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1038), .Y(div_n_T_87[13]) );
  AO22X1_LVT div_ashr_12_U942 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_70_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_62_), .Y(div_ashr_12_n1000) );
  AO22X1_LVT div_ashr_12_U941 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_54_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_46_), .Y(div_ashr_12_n998) );
  AO22X1_LVT div_ashr_12_U940 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1000), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n998), .Y(div_ashr_12_n940) );
  AO22X1_LVT div_ashr_12_U939 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_38_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_30_), .Y(div_ashr_12_n999) );
  AO22X1_LVT div_ashr_12_U938 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_22_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_14_), .Y(div_ashr_12_n1037) );
  AO22X1_LVT div_ashr_12_U937 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n999), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1037), .Y(div_ashr_12_n1036)
         );
  AO22X1_LVT div_ashr_12_U936 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n940), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1036), .Y(div_n_T_87[14]) );
  AO22X1_LVT div_ashr_12_U935 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_71_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_63_), .Y(div_ashr_12_n996) );
  AO22X1_LVT div_ashr_12_U934 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_55_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_47_), .Y(div_ashr_12_n994) );
  AO22X1_LVT div_ashr_12_U933 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n996), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n994), .Y(div_ashr_12_n937) );
  AO22X1_LVT div_ashr_12_U932 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_39_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_31_), .Y(div_ashr_12_n995) );
  AO22X1_LVT div_ashr_12_U931 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_23_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_15_), .Y(div_ashr_12_n1035) );
  AO22X1_LVT div_ashr_12_U930 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n995), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1035), .Y(div_ashr_12_n1034)
         );
  AO22X1_LVT div_ashr_12_U929 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n937), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1034), .Y(div_n_T_87[15]) );
  AO22X1_LVT div_ashr_12_U928 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_72_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_64_), .Y(div_ashr_12_n992) );
  AO22X1_LVT div_ashr_12_U927 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n992), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1033), .Y(div_ashr_12_n934) );
  AO22X1_LVT div_ashr_12_U926 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_73_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_65_), .Y(div_ashr_12_n990) );
  AO22X1_LVT div_ashr_12_U925 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_57_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_49_), .Y(div_ashr_12_n1026) );
  AO22X1_LVT div_ashr_12_U924 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n990), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1026), .Y(div_ashr_12_n931) );
  AO22X1_LVT div_ashr_12_U923 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_41_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_33_), .Y(div_ashr_12_n1027) );
  AO22X1_LVT div_ashr_12_U922 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_25_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_17_), .Y(div_ashr_12_n1025) );
  AO22X1_LVT div_ashr_12_U921 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1027), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1025), .Y(div_ashr_12_n1030)
         );
  AO22X1_LVT div_ashr_12_U920 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n931), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1030), .Y(div_n_T_87[17]) );
  AO22X1_LVT div_ashr_12_U919 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_74_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_66_), .Y(div_ashr_12_n987) );
  AO22X1_LVT div_ashr_12_U918 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_58_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_50_), .Y(div_ashr_12_n1002) );
  AO22X1_LVT div_ashr_12_U917 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n987), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1002), .Y(div_ashr_12_n925) );
  AO22X1_LVT div_ashr_12_U916 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_42_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_34_), .Y(div_ashr_12_n1003) );
  AO22X1_LVT div_ashr_12_U915 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_26_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_18_), .Y(div_ashr_12_n1001) );
  AO22X1_LVT div_ashr_12_U914 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1003), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1001), .Y(div_ashr_12_n1029)
         );
  AO22X1_LVT div_ashr_12_U913 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n925), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1029), .Y(div_n_T_87[18]) );
  AO22X1_LVT div_ashr_12_U912 ( .A1(div_n300), .A2(div_n_T_51_75_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_67_), .Y(div_ashr_12_n984) );
  AO22X1_LVT div_ashr_12_U911 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_59_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_51_), .Y(div_ashr_12_n982) );
  AO22X1_LVT div_ashr_12_U910 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n984), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n982), .Y(div_ashr_12_n921) );
  AO22X1_LVT div_ashr_12_U909 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_43_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_35_), .Y(div_ashr_12_n983) );
  AO22X1_LVT div_ashr_12_U908 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_27_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_19_), .Y(div_ashr_12_n963) );
  AO22X1_LVT div_ashr_12_U907 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n983), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n963), .Y(div_ashr_12_n1028) );
  AO22X1_LVT div_ashr_12_U906 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n921), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1028), .Y(div_n_T_87[19]) );
  AO22X1_LVT div_ashr_12_U905 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1026), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1027), .Y(div_ashr_12_n989) );
  AO22X1_LVT div_ashr_12_U904 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_76_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_68_), .Y(div_ashr_12_n980) );
  AO22X1_LVT div_ashr_12_U903 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_60_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_52_), .Y(div_ashr_12_n978) );
  AO22X1_LVT div_ashr_12_U902 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n980), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n978), .Y(div_ashr_12_n918) );
  AO22X1_LVT div_ashr_12_U901 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_44_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_36_), .Y(div_ashr_12_n979) );
  AO22X1_LVT div_ashr_12_U900 ( .A1(div_n300), .A2(div_n_T_51_28_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_20_), .Y(div_ashr_12_n929) );
  AO22X1_LVT div_ashr_12_U899 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n979), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n929), .Y(div_ashr_12_n1024) );
  AO22X1_LVT div_ashr_12_U898 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n918), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1024), .Y(div_n_T_87[20]) );
  AO22X1_LVT div_ashr_12_U897 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_77_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_69_), .Y(div_ashr_12_n976) );
  AO22X1_LVT div_ashr_12_U896 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_61_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_53_), .Y(div_ashr_12_n974) );
  AO22X1_LVT div_ashr_12_U895 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n976), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n974), .Y(div_ashr_12_n915) );
  AO22X1_LVT div_ashr_12_U894 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_45_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_37_), .Y(div_ashr_12_n975) );
  AO22X1_LVT div_ashr_12_U893 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_29_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_21_), .Y(div_ashr_12_n890) );
  AO22X1_LVT div_ashr_12_U892 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n975), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n890), .Y(div_ashr_12_n1023) );
  AO22X1_LVT div_ashr_12_U891 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n915), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1023), .Y(div_n_T_87[21]) );
  AO22X1_LVT div_ashr_12_U890 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_78_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_70_), .Y(div_ashr_12_n972) );
  AO22X1_LVT div_ashr_12_U889 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_62_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_54_), .Y(div_ashr_12_n970) );
  AO22X1_LVT div_ashr_12_U888 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n972), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n970), .Y(div_ashr_12_n911) );
  AO22X1_LVT div_ashr_12_U887 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_46_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_38_), .Y(div_ashr_12_n971) );
  AO22X1_LVT div_ashr_12_U886 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_30_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_22_), .Y(div_ashr_12_n870) );
  AO22X1_LVT div_ashr_12_U885 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n971), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n870), .Y(div_ashr_12_n1022) );
  AO22X1_LVT div_ashr_12_U884 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n911), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1022), .Y(div_n_T_87[22]) );
  AO22X1_LVT div_ashr_12_U883 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_79_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_71_), .Y(div_ashr_12_n968) );
  AO22X1_LVT div_ashr_12_U882 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_63_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_55_), .Y(div_ashr_12_n966) );
  AO22X1_LVT div_ashr_12_U881 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n968), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n966), .Y(div_ashr_12_n907) );
  AO22X1_LVT div_ashr_12_U880 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_47_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_39_), .Y(div_ashr_12_n967) );
  AO22X1_LVT div_ashr_12_U879 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_31_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_23_), .Y(div_ashr_12_n866) );
  AO22X1_LVT div_ashr_12_U878 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n967), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n866), .Y(div_ashr_12_n1021) );
  AO22X1_LVT div_ashr_12_U877 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n907), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1021), .Y(div_n_T_87[23]) );
  AO22X1_LVT div_ashr_12_U876 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_80_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_72_), .Y(div_ashr_12_n960) );
  AO22X1_LVT div_ashr_12_U875 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_64_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_56_), .Y(div_ashr_12_n958) );
  AO22X1_LVT div_ashr_12_U874 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n960), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n958), .Y(div_ashr_12_n904) );
  AO22X1_LVT div_ashr_12_U873 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_48_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_40_), .Y(div_ashr_12_n959) );
  AO22X1_LVT div_ashr_12_U872 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_32_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_24_), .Y(div_ashr_12_n862) );
  AO22X1_LVT div_ashr_12_U871 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_81_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_73_), .Y(div_ashr_12_n957) );
  AO22X1_LVT div_ashr_12_U870 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_65_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_57_), .Y(div_ashr_12_n955) );
  AO22X1_LVT div_ashr_12_U869 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n957), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n955), .Y(div_ashr_12_n901) );
  AO22X1_LVT div_ashr_12_U868 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_49_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_41_), .Y(div_ashr_12_n956) );
  AO22X1_LVT div_ashr_12_U867 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_33_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_25_), .Y(div_ashr_12_n858) );
  AO22X1_LVT div_ashr_12_U866 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n956), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n858), .Y(div_ashr_12_n1020) );
  AO22X1_LVT div_ashr_12_U865 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n901), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1020), .Y(div_n_T_87[25]) );
  AO22X1_LVT div_ashr_12_U864 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_82_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_74_), .Y(div_ashr_12_n953) );
  AO22X1_LVT div_ashr_12_U863 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n953), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1019), .Y(div_ashr_12_n897) );
  AO22X1_LVT div_ashr_12_U862 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1017), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1018), .Y(div_ashr_12_n1016)
         );
  AO22X1_LVT div_ashr_12_U861 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n897), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1016), .Y(div_n_T_87[26]) );
  AO22X1_LVT div_ashr_12_U860 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_83_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_75_), .Y(div_ashr_12_n950) );
  AO22X1_LVT div_ashr_12_U859 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n950), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1015), .Y(div_ashr_12_n893) );
  AO22X1_LVT div_ashr_12_U858 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1013), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1014), .Y(div_ashr_12_n1012)
         );
  AO22X1_LVT div_ashr_12_U857 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n893), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1012), .Y(div_n_T_87[27]) );
  AO22X1_LVT div_ashr_12_U856 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_84_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_76_), .Y(div_ashr_12_n947) );
  AO22X1_LVT div_ashr_12_U855 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n947), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1011), .Y(div_ashr_12_n885) );
  AO22X1_LVT div_ashr_12_U854 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1009), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1010), .Y(div_ashr_12_n1008)
         );
  AO22X1_LVT div_ashr_12_U853 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n885), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1008), .Y(div_n_T_87[28]) );
  AO22X1_LVT div_ashr_12_U852 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_85_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_77_), .Y(div_ashr_12_n944) );
  AO22X1_LVT div_ashr_12_U851 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n944), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1007), .Y(div_ashr_12_n881) );
  AO22X1_LVT div_ashr_12_U850 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1005), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1006), .Y(div_ashr_12_n1004)
         );
  AO22X1_LVT div_ashr_12_U849 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n881), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n1004), .Y(div_n_T_87[29]) );
  AO22X1_LVT div_ashr_12_U848 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1002), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1003), .Y(div_ashr_12_n986) );
  AO22X1_LVT div_ashr_12_U847 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_86_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_78_), .Y(div_ashr_12_n941) );
  AO22X1_LVT div_ashr_12_U846 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n941), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1000), .Y(div_ashr_12_n877) );
  AO22X1_LVT div_ashr_12_U845 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n998), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n999), .Y(div_ashr_12_n997) );
  AO22X1_LVT div_ashr_12_U844 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n877), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n997), .Y(div_n_T_87[30]) );
  AO22X1_LVT div_ashr_12_U843 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_87_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_79_), .Y(div_ashr_12_n938) );
  AO22X1_LVT div_ashr_12_U842 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n938), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n996), .Y(div_ashr_12_n873) );
  AO22X1_LVT div_ashr_12_U841 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n994), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n995), .Y(div_ashr_12_n993) );
  AO22X1_LVT div_ashr_12_U840 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n873), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n993), .Y(div_n_T_87[31]) );
  AO22X1_LVT div_ashr_12_U839 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_88_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_80_), .Y(div_ashr_12_n935) );
  AO22X1_LVT div_ashr_12_U838 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_89_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_81_), .Y(div_ashr_12_n933) );
  AO22X1_LVT div_ashr_12_U837 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n933), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n990), .Y(div_ashr_12_n988) );
  AO22X1_LVT div_ashr_12_U836 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n988), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n989), .Y(div_n_T_87[33]) );
  AO22X1_LVT div_ashr_12_U835 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_90_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_82_), .Y(div_ashr_12_n927) );
  AO22X1_LVT div_ashr_12_U834 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n927), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n987), .Y(div_ashr_12_n985) );
  AO22X1_LVT div_ashr_12_U833 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n985), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n986), .Y(div_n_T_87[34]) );
  AO22X1_LVT div_ashr_12_U832 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_91_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_83_), .Y(div_ashr_12_n923) );
  AO22X1_LVT div_ashr_12_U831 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n923), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n984), .Y(div_ashr_12_n981) );
  AO22X1_LVT div_ashr_12_U830 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n982), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n983), .Y(div_ashr_12_n961) );
  AO22X1_LVT div_ashr_12_U829 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n981), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n961), .Y(div_n_T_87[35]) );
  AO22X1_LVT div_ashr_12_U828 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_92_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_84_), .Y(div_ashr_12_n919) );
  AO22X1_LVT div_ashr_12_U827 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n919), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n980), .Y(div_ashr_12_n977) );
  AO22X1_LVT div_ashr_12_U826 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n978), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n979), .Y(div_ashr_12_n928) );
  AO22X1_LVT div_ashr_12_U825 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n977), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n928), .Y(div_n_T_87[36]) );
  AO22X1_LVT div_ashr_12_U824 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_93_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_85_), .Y(div_ashr_12_n917) );
  AO22X1_LVT div_ashr_12_U823 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n917), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n976), .Y(div_ashr_12_n973) );
  AO22X1_LVT div_ashr_12_U822 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n974), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n975), .Y(div_ashr_12_n888) );
  AO22X1_LVT div_ashr_12_U821 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n973), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n888), .Y(div_n_T_87[37]) );
  AO22X1_LVT div_ashr_12_U820 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_94_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_86_), .Y(div_ashr_12_n913) );
  AO22X1_LVT div_ashr_12_U819 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n913), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n972), .Y(div_ashr_12_n969) );
  AO22X1_LVT div_ashr_12_U818 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n970), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n971), .Y(div_ashr_12_n868) );
  AO22X1_LVT div_ashr_12_U817 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n969), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n868), .Y(div_n_T_87[38]) );
  AO22X1_LVT div_ashr_12_U816 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_95_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_87_), .Y(div_ashr_12_n909) );
  AO22X1_LVT div_ashr_12_U815 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n909), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n968), .Y(div_ashr_12_n965) );
  AO22X1_LVT div_ashr_12_U814 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n966), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n967), .Y(div_ashr_12_n864) );
  AO22X1_LVT div_ashr_12_U813 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n965), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n864), .Y(div_n_T_87[39]) );
  AO22X1_LVT div_ashr_12_U812 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_11_), 
        .A3(div_ashr_12_n852), .A4(div_n305), .Y(div_ashr_12_n964) );
  AO22X1_LVT div_ashr_12_U811 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n963), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n964), .Y(div_ashr_12_n962) );
  AO22X1_LVT div_ashr_12_U810 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n961), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n962), .Y(div_n_T_87[3]) );
  AO22X1_LVT div_ashr_12_U809 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_96_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_88_), .Y(div_ashr_12_n905) );
  AO22X1_LVT div_ashr_12_U808 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n958), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n959), .Y(div_ashr_12_n860) );
  AO22X1_LVT div_ashr_12_U807 ( .A1(div_n300), .A2(div_n_T_51_97_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_89_), .Y(div_ashr_12_n903) );
  AO22X1_LVT div_ashr_12_U806 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n903), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n957), .Y(div_ashr_12_n954) );
  AO22X1_LVT div_ashr_12_U805 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n955), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n956), .Y(div_ashr_12_n856) );
  AO22X1_LVT div_ashr_12_U804 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n954), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n856), .Y(div_n_T_87[41]) );
  AO22X1_LVT div_ashr_12_U803 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_98_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_90_), .Y(div_ashr_12_n899) );
  AO22X1_LVT div_ashr_12_U802 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n899), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n953), .Y(div_ashr_12_n951) );
  AO22X1_LVT div_ashr_12_U801 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n951), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n952), .Y(div_n_T_87[42]) );
  AO22X1_LVT div_ashr_12_U800 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_99_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_91_), .Y(div_ashr_12_n895) );
  AO22X1_LVT div_ashr_12_U799 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n895), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n950), .Y(div_ashr_12_n948) );
  AO22X1_LVT div_ashr_12_U798 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n948), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n949), .Y(div_n_T_87[43]) );
  AO22X1_LVT div_ashr_12_U797 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_100_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_92_), .Y(div_ashr_12_n887) );
  AO22X1_LVT div_ashr_12_U796 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n887), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n947), .Y(div_ashr_12_n945) );
  AO22X1_LVT div_ashr_12_U795 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n945), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n946), .Y(div_n_T_87[44]) );
  AO22X1_LVT div_ashr_12_U794 ( .A1(div_n300), .A2(div_n_T_51_101_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_93_), .Y(div_ashr_12_n883) );
  AO22X1_LVT div_ashr_12_U793 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n883), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n944), .Y(div_ashr_12_n942) );
  AO22X1_LVT div_ashr_12_U792 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n942), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n943), .Y(div_n_T_87[45]) );
  AO22X1_LVT div_ashr_12_U791 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_102_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_94_), .Y(div_ashr_12_n879) );
  AO22X1_LVT div_ashr_12_U790 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n879), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n941), .Y(div_ashr_12_n939) );
  AO22X1_LVT div_ashr_12_U789 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n939), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n940), .Y(div_n_T_87[46]) );
  AO22X1_LVT div_ashr_12_U788 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_103_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_95_), .Y(div_ashr_12_n875) );
  AO22X1_LVT div_ashr_12_U787 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n875), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n938), .Y(div_ashr_12_n936) );
  AO22X1_LVT div_ashr_12_U786 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n936), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n937), .Y(div_n_T_87[47]) );
  AO22X1_LVT div_ashr_12_U785 ( .A1(div_n300), .A2(div_n_T_51_105_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_97_), .Y(div_ashr_12_n932) );
  AO22X1_LVT div_ashr_12_U784 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n932), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n933), .Y(div_ashr_12_n930) );
  AO22X1_LVT div_ashr_12_U783 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n930), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n931), .Y(div_n_T_87[49]) );
  AO22X1_LVT div_ashr_12_U782 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_106_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_98_), .Y(div_ashr_12_n926) );
  AO22X1_LVT div_ashr_12_U781 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n926), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n927), .Y(div_ashr_12_n924) );
  AO22X1_LVT div_ashr_12_U780 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n924), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n925), .Y(div_n_T_87[50]) );
  AO22X1_LVT div_ashr_12_U779 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_107_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_99_), .Y(div_ashr_12_n922) );
  AO22X1_LVT div_ashr_12_U778 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n922), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n923), .Y(div_ashr_12_n920) );
  AO22X1_LVT div_ashr_12_U777 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n920), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n921), .Y(div_n_T_87[51]) );
  AO22X1_LVT div_ashr_12_U776 ( .A1(div_n300), .A2(div_n_T_51_109_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_101_), .Y(div_ashr_12_n916) );
  AO22X1_LVT div_ashr_12_U775 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n916), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n917), .Y(div_ashr_12_n914) );
  AO22X1_LVT div_ashr_12_U774 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n914), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n915), .Y(div_n_T_87[53]) );
  AO22X1_LVT div_ashr_12_U773 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_110_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_102_), .Y(div_ashr_12_n912) );
  AO22X1_LVT div_ashr_12_U772 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n912), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n913), .Y(div_ashr_12_n910) );
  AO22X1_LVT div_ashr_12_U771 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n910), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n911), .Y(div_n_T_87[54]) );
  AO22X1_LVT div_ashr_12_U770 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_111_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_103_), .Y(div_ashr_12_n908) );
  AO22X1_LVT div_ashr_12_U769 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n908), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n909), .Y(div_ashr_12_n906) );
  AO22X1_LVT div_ashr_12_U768 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n906), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n907), .Y(div_n_T_87[55]) );
  AO22X1_LVT div_ashr_12_U767 ( .A1(div_n300), .A2(div_n_T_51_113_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_105_), .Y(div_ashr_12_n902) );
  AO22X1_LVT div_ashr_12_U766 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n902), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n903), .Y(div_ashr_12_n900) );
  AO22X1_LVT div_ashr_12_U765 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n900), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n901), .Y(div_n_T_87[57]) );
  AO22X1_LVT div_ashr_12_U764 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_114_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_106_), .Y(div_ashr_12_n898) );
  AO22X1_LVT div_ashr_12_U763 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n898), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n899), .Y(div_ashr_12_n896) );
  AO22X1_LVT div_ashr_12_U762 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n896), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n897), .Y(div_n_T_87[58]) );
  AO22X1_LVT div_ashr_12_U761 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_115_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_107_), .Y(div_ashr_12_n894) );
  AO22X1_LVT div_ashr_12_U760 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n894), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n895), .Y(div_ashr_12_n892) );
  AO22X1_LVT div_ashr_12_U759 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n892), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n893), .Y(div_n_T_87[59]) );
  AO22X1_LVT div_ashr_12_U758 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_13_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_5_), .Y(div_ashr_12_n891) );
  AO22X1_LVT div_ashr_12_U757 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n890), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n891), .Y(div_ashr_12_n889) );
  AO22X1_LVT div_ashr_12_U756 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n888), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n889), .Y(div_n_T_87[5]) );
  AO22X1_LVT div_ashr_12_U755 ( .A1(div_n300), .A2(div_n_T_51_116_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_108_), .Y(div_ashr_12_n886) );
  AO22X1_LVT div_ashr_12_U754 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n886), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n887), .Y(div_ashr_12_n884) );
  AO22X1_LVT div_ashr_12_U753 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n884), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n885), .Y(div_n_T_87[60]) );
  AO22X1_LVT div_ashr_12_U752 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_117_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_109_), .Y(div_ashr_12_n882) );
  AO22X1_LVT div_ashr_12_U751 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n882), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n883), .Y(div_ashr_12_n880) );
  AO22X1_LVT div_ashr_12_U750 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n880), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n881), .Y(div_n_T_87[61]) );
  AO22X1_LVT div_ashr_12_U749 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_118_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_110_), .Y(div_ashr_12_n878) );
  AO22X1_LVT div_ashr_12_U748 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n878), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n879), .Y(div_ashr_12_n876) );
  AO22X1_LVT div_ashr_12_U747 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n876), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n877), .Y(div_n_T_87[62]) );
  AO22X1_LVT div_ashr_12_U746 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_119_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_111_), .Y(div_ashr_12_n874) );
  AO22X1_LVT div_ashr_12_U745 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n874), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n875), .Y(div_ashr_12_n872) );
  AO22X1_LVT div_ashr_12_U744 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n872), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n873), .Y(div_n_T_87[63]) );
  AO22X1_LVT div_ashr_12_U743 ( .A1(div_n300), .A2(div_n_T_51_14_), .A3(
        div_ashr_12_n852), .A4(div_n307), .Y(div_ashr_12_n871) );
  AO22X1_LVT div_ashr_12_U742 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n870), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n871), .Y(div_ashr_12_n869) );
  AO22X1_LVT div_ashr_12_U741 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n868), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n869), .Y(div_n_T_87[6]) );
  AO22X1_LVT div_ashr_12_U740 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_15_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_7_), .Y(div_ashr_12_n867) );
  AO22X1_LVT div_ashr_12_U739 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n866), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n867), .Y(div_ashr_12_n865) );
  AO22X1_LVT div_ashr_12_U738 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n864), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n865), .Y(div_n_T_87[7]) );
  AO22X1_LVT div_ashr_12_U737 ( .A1(div_n300), .A2(div_n_T_51_16_), .A3(
        div_ashr_12_n852), .A4(div_n_T_51_8_), .Y(div_ashr_12_n863) );
  AO22X1_LVT div_ashr_12_U736 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n862), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n863), .Y(div_ashr_12_n861) );
  AO22X1_LVT div_ashr_12_U735 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n860), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n861), .Y(div_n_T_87[8]) );
  AO22X1_LVT div_ashr_12_U734 ( .A1(div_ashr_12_n853), .A2(div_n_T_51_17_), 
        .A3(div_ashr_12_n852), .A4(div_n_T_51_9_), .Y(div_ashr_12_n859) );
  AO22X1_LVT div_ashr_12_U733 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n858), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n859), .Y(div_ashr_12_n857) );
  AO22X1_LVT div_ashr_12_U732 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n856), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n857), .Y(div_n_T_87[9]) );
  INVX1_LVT div_ashr_12_U731 ( .A(div_n_T_85_4_), .Y(div_ashr_12_n854) );
  INVX1_LVT div_ashr_12_U730 ( .A(div_n_T_85_5_), .Y(div_ashr_12_n855) );
  INVX1_LVT div_ashr_12_U729 ( .A(div_ashr_12_n852), .Y(div_ashr_12_n853) );
  INVX1_LVT div_ashr_12_U728 ( .A(div_n300), .Y(div_ashr_12_n852) );
  AO22X1_LVT div_ashr_12_U727 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n851), 
        .A3(div_ashr_12_n918), .A4(div_ashr_12_n855), .Y(div_n_T_87[52]) );
  AO22X1_LVT div_ashr_12_U726 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n850), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n919), .Y(div_ashr_12_n851) );
  AO22X1_LVT div_ashr_12_U725 ( .A1(div_ashr_12_n852), .A2(div_n_T_51_100_), 
        .A3(div_ashr_12_n853), .A4(div_n_T_51_108_), .Y(div_ashr_12_n850) );
  AO22X1_LVT div_ashr_12_U724 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n849), 
        .A3(div_ashr_12_n991), .A4(div_ashr_12_n855), .Y(div_n_T_87[32]) );
  AO22X1_LVT div_ashr_12_U723 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n935), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n992), .Y(div_ashr_12_n849) );
  AO22X1_LVT div_ashr_12_U722 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n989), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n848), .Y(div_n_T_87[1]) );
  AO22X1_LVT div_ashr_12_U721 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1025), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n847), .Y(div_ashr_12_n848) );
  AO22X1_LVT div_ashr_12_U720 ( .A1(div_n300), .A2(div_n_T_51_9_), .A3(
        div_ashr_12_n852), .A4(div_n303), .Y(div_ashr_12_n847) );
  AO22X1_LVT div_ashr_12_U719 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n991), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n846), .Y(div_n_T_87[0]) );
  AO22X1_LVT div_ashr_12_U718 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1032), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n845), .Y(div_ashr_12_n846) );
  AO22X1_LVT div_ashr_12_U717 ( .A1(div_ashr_12_n852), .A2(div_n302), .A3(
        div_ashr_12_n853), .A4(div_n_T_51_8_), .Y(div_ashr_12_n845) );
  AO22X1_LVT div_ashr_12_U716 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n928), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n844), .Y(div_n_T_87[4]) );
  AO22X1_LVT div_ashr_12_U715 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n929), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n843), .Y(div_ashr_12_n844) );
  AO22X1_LVT div_ashr_12_U714 ( .A1(div_ashr_12_n852), .A2(div_n306), .A3(
        div_n_T_51_12_), .A4(div_ashr_12_n853), .Y(div_ashr_12_n843) );
  AO22X1_LVT div_ashr_12_U713 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n934), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n842), .Y(div_n_T_87[16]) );
  AO22X1_LVT div_ashr_12_U712 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1031), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n1032), .Y(div_ashr_12_n842) );
  AO22X1_LVT div_ashr_12_U711 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n986), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n841), .Y(div_n_T_87[2]) );
  AO22X1_LVT div_ashr_12_U710 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1001), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n840), .Y(div_ashr_12_n841) );
  AO22X1_LVT div_ashr_12_U709 ( .A1(div_ashr_12_n852), .A2(div_n304), .A3(
        div_ashr_12_n853), .A4(div_n_T_51_10_), .Y(div_ashr_12_n840) );
  AO22X1_LVT div_ashr_12_U708 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n904), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n839), .Y(div_n_T_87[24]) );
  AO22X1_LVT div_ashr_12_U707 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n959), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n862), .Y(div_ashr_12_n839) );
  AO22X1_LVT div_ashr_12_U706 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n838), 
        .A3(div_ashr_12_n860), .A4(div_ashr_12_n855), .Y(div_n_T_87[40]) );
  AO22X1_LVT div_ashr_12_U705 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n905), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n960), .Y(div_ashr_12_n838) );
  AO22X1_LVT div_ashr_12_U704 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n946), 
        .A3(div_ashr_12_n855), .A4(div_ashr_12_n837), .Y(div_n_T_87[12]) );
  AO22X1_LVT div_ashr_12_U703 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n1010), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n836), .Y(div_ashr_12_n837) );
  AO22X1_LVT div_ashr_12_U702 ( .A1(div_n_T_51_12_), .A2(div_ashr_12_n852), 
        .A3(div_n_T_51_20_), .A4(div_ashr_12_n853), .Y(div_ashr_12_n836) );
  AO22X1_LVT div_ashr_12_U701 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n835), 
        .A3(div_ashr_12_n934), .A4(div_ashr_12_n855), .Y(div_n_T_87[48]) );
  AO22X1_LVT div_ashr_12_U700 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n834), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n935), .Y(div_ashr_12_n835) );
  AO22X1_LVT div_ashr_12_U699 ( .A1(div_ashr_12_n852), .A2(div_n_T_51_96_), 
        .A3(div_ashr_12_n853), .A4(div_n_T_51_104_), .Y(div_ashr_12_n834) );
  AO22X1_LVT div_ashr_12_U698 ( .A1(div_n_T_85_5_), .A2(div_ashr_12_n833), 
        .A3(div_ashr_12_n904), .A4(div_ashr_12_n855), .Y(div_n_T_87[56]) );
  AO22X1_LVT div_ashr_12_U697 ( .A1(div_n_T_85_4_), .A2(div_ashr_12_n832), 
        .A3(div_ashr_12_n854), .A4(div_ashr_12_n905), .Y(div_ashr_12_n833) );
  AO22X1_LVT div_ashr_12_U696 ( .A1(div_ashr_12_n852), .A2(div_n_T_51_104_), 
        .A3(div_ashr_12_n853), .A4(div_n_T_51_112_), .Y(div_ashr_12_n832) );
  OR3X1_LVT div_sub_x_9_U395 ( .A1(div_result_3_), .A2(div_result_2_), .A3(
        div_sub_x_9_n388), .Y(div_sub_x_9_n412) );
  OR3X1_LVT div_sub_x_9_U394 ( .A1(div_result_5_), .A2(div_result_4_), .A3(
        div_sub_x_9_n412), .Y(div_sub_x_9_n394) );
  OR3X1_LVT div_sub_x_9_U393 ( .A1(div_result_7_), .A2(div_result_6_), .A3(
        div_sub_x_9_n394), .Y(div_sub_x_9_n392) );
  OR3X1_LVT div_sub_x_9_U392 ( .A1(div_result_9_), .A2(div_result_8_), .A3(
        div_sub_x_9_n392), .Y(div_sub_x_9_n465) );
  HADDX1_LVT div_sub_x_9_U391 ( .A0(div_result_10_), .B0(div_sub_x_9_n465), 
        .SO(div_negated_remainder[10]) );
  OR2X1_LVT div_sub_x_9_U390 ( .A1(div_result_10_), .A2(div_sub_x_9_n465), .Y(
        div_sub_x_9_n464) );
  HADDX1_LVT div_sub_x_9_U389 ( .A0(div_sub_x_9_n464), .B0(div_result_11_), 
        .SO(div_negated_remainder[11]) );
  NAND2X0_LVT div_sub_x_9_U388 ( .A1(div_sub_x_9_n384), .A2(div_sub_x_9_n463), 
        .Y(div_sub_x_9_n461) );
  NAND2X0_LVT div_sub_x_9_U387 ( .A1(div_sub_x_9_n381), .A2(div_sub_x_9_n382), 
        .Y(div_sub_x_9_n462) );
  HADDX1_LVT div_sub_x_9_U386 ( .A0(div_sub_x_9_n462), .B0(div_result_13_), 
        .SO(div_negated_remainder[13]) );
  OR3X1_LVT div_sub_x_9_U385 ( .A1(div_result_13_), .A2(div_result_12_), .A3(
        div_sub_x_9_n461), .Y(div_sub_x_9_n459) );
  HADDX1_LVT div_sub_x_9_U384 ( .A0(div_result_14_), .B0(div_sub_x_9_n459), 
        .SO(div_negated_remainder[14]) );
  OR2X1_LVT div_sub_x_9_U383 ( .A1(div_result_14_), .A2(div_sub_x_9_n459), .Y(
        div_sub_x_9_n460) );
  HADDX1_LVT div_sub_x_9_U382 ( .A0(div_sub_x_9_n460), .B0(div_result_15_), 
        .SO(div_negated_remainder[15]) );
  OR3X1_LVT div_sub_x_9_U381 ( .A1(div_result_15_), .A2(div_result_14_), .A3(
        div_sub_x_9_n459), .Y(div_sub_x_9_n453) );
  NAND2X0_LVT div_sub_x_9_U380 ( .A1(div_sub_x_9_n380), .A2(div_sub_x_9_n379), 
        .Y(div_sub_x_9_n458) );
  HADDX1_LVT div_sub_x_9_U379 ( .A0(div_result_17_), .B0(div_sub_x_9_n458), 
        .SO(div_negated_remainder[17]) );
  OR2X1_LVT div_sub_x_9_U378 ( .A1(div_result_17_), .A2(div_result_16_), .Y(
        div_sub_x_9_n455) );
  OR2X1_LVT div_sub_x_9_U377 ( .A1(div_sub_x_9_n453), .A2(div_sub_x_9_n455), 
        .Y(div_sub_x_9_n457) );
  HADDX1_LVT div_sub_x_9_U376 ( .A0(div_result_18_), .B0(div_sub_x_9_n457), 
        .SO(div_negated_remainder[18]) );
  OR3X1_LVT div_sub_x_9_U375 ( .A1(div_result_18_), .A2(div_sub_x_9_n455), 
        .A3(div_sub_x_9_n453), .Y(div_sub_x_9_n456) );
  HADDX1_LVT div_sub_x_9_U374 ( .A0(div_result_19_), .B0(div_sub_x_9_n456), 
        .SO(div_negated_remainder[19]) );
  OR3X1_LVT div_sub_x_9_U373 ( .A1(div_result_19_), .A2(div_result_18_), .A3(
        div_sub_x_9_n455), .Y(div_sub_x_9_n448) );
  OR2X1_LVT div_sub_x_9_U372 ( .A1(div_sub_x_9_n453), .A2(div_sub_x_9_n448), 
        .Y(div_sub_x_9_n451) );
  HADDX1_LVT div_sub_x_9_U371 ( .A0(div_result_20_), .B0(div_sub_x_9_n451), 
        .SO(div_negated_remainder[20]) );
  OR2X1_LVT div_sub_x_9_U370 ( .A1(div_result_20_), .A2(div_sub_x_9_n451), .Y(
        div_sub_x_9_n454) );
  HADDX1_LVT div_sub_x_9_U369 ( .A0(div_sub_x_9_n454), .B0(div_result_21_), 
        .SO(div_negated_remainder[21]) );
  OR2X1_LVT div_sub_x_9_U368 ( .A1(div_result_21_), .A2(div_result_20_), .Y(
        div_sub_x_9_n449) );
  OR3X1_LVT div_sub_x_9_U367 ( .A1(div_sub_x_9_n453), .A2(div_sub_x_9_n448), 
        .A3(div_sub_x_9_n449), .Y(div_sub_x_9_n452) );
  HADDX1_LVT div_sub_x_9_U366 ( .A0(div_result_22_), .B0(div_sub_x_9_n452), 
        .SO(div_negated_remainder[22]) );
  OR3X1_LVT div_sub_x_9_U365 ( .A1(div_result_22_), .A2(div_sub_x_9_n449), 
        .A3(div_sub_x_9_n451), .Y(div_sub_x_9_n450) );
  HADDX1_LVT div_sub_x_9_U364 ( .A0(div_result_23_), .B0(div_sub_x_9_n450), 
        .SO(div_negated_remainder[23]) );
  NAND2X0_LVT div_sub_x_9_U363 ( .A1(div_sub_x_9_n380), .A2(div_sub_x_9_n447), 
        .Y(div_sub_x_9_n445) );
  NAND2X0_LVT div_sub_x_9_U362 ( .A1(div_sub_x_9_n378), .A2(div_sub_x_9_n377), 
        .Y(div_sub_x_9_n446) );
  HADDX1_LVT div_sub_x_9_U361 ( .A0(div_result_25_), .B0(div_sub_x_9_n446), 
        .SO(div_negated_remainder[25]) );
  OR3X1_LVT div_sub_x_9_U360 ( .A1(div_result_25_), .A2(div_result_24_), .A3(
        div_sub_x_9_n445), .Y(div_sub_x_9_n444) );
  HADDX1_LVT div_sub_x_9_U359 ( .A0(div_result_26_), .B0(div_sub_x_9_n444), 
        .SO(div_negated_remainder[26]) );
  OR2X1_LVT div_sub_x_9_U358 ( .A1(div_result_26_), .A2(div_sub_x_9_n444), .Y(
        div_sub_x_9_n443) );
  HADDX1_LVT div_sub_x_9_U357 ( .A0(div_sub_x_9_n443), .B0(div_result_27_), 
        .SO(div_negated_remainder[27]) );
  NAND2X0_LVT div_sub_x_9_U356 ( .A1(div_sub_x_9_n440), .A2(div_sub_x_9_n378), 
        .Y(div_sub_x_9_n438) );
  HADDX1_LVT div_sub_x_9_U355 ( .A0(div_result_28_), .B0(div_sub_x_9_n438), 
        .SO(div_negated_remainder[28]) );
  NAND3X0_LVT div_sub_x_9_U354 ( .A1(div_sub_x_9_n440), .A2(div_sub_x_9_n378), 
        .A3(div_sub_x_9_n376), .Y(div_sub_x_9_n442) );
  HADDX1_LVT div_sub_x_9_U353 ( .A0(div_result_29_), .B0(div_sub_x_9_n442), 
        .SO(div_negated_remainder[29]) );
  OR2X1_LVT div_sub_x_9_U352 ( .A1(div_result_29_), .A2(div_result_28_), .Y(
        div_sub_x_9_n437) );
  NAND3X0_LVT div_sub_x_9_U351 ( .A1(div_sub_x_9_n440), .A2(div_sub_x_9_n375), 
        .A3(div_sub_x_9_n378), .Y(div_sub_x_9_n441) );
  HADDX1_LVT div_sub_x_9_U350 ( .A0(div_result_30_), .B0(div_sub_x_9_n441), 
        .SO(div_negated_remainder[30]) );
  NAND4X0_LVT div_sub_x_9_U349 ( .A1(div_sub_x_9_n375), .A2(div_sub_x_9_n440), 
        .A3(div_sub_x_9_n378), .A4(div_sub_x_9_n374), .Y(div_sub_x_9_n439) );
  HADDX1_LVT div_sub_x_9_U348 ( .A0(div_result_31_), .B0(div_sub_x_9_n439), 
        .SO(div_negated_remainder[31]) );
  NAND2X0_LVT div_sub_x_9_U347 ( .A1(div_sub_x_9_n424), .A2(div_sub_x_9_n372), 
        .Y(div_sub_x_9_n436) );
  HADDX1_LVT div_sub_x_9_U346 ( .A0(div_result_33_), .B0(div_sub_x_9_n436), 
        .SO(div_negated_remainder[33]) );
  OR2X1_LVT div_sub_x_9_U345 ( .A1(div_result_33_), .A2(div_result_32_), .Y(
        div_sub_x_9_n433) );
  OR2X1_LVT div_sub_x_9_U344 ( .A1(div_sub_x_9_n373), .A2(div_sub_x_9_n433), 
        .Y(div_sub_x_9_n435) );
  HADDX1_LVT div_sub_x_9_U343 ( .A0(div_result_34_), .B0(div_sub_x_9_n435), 
        .SO(div_negated_remainder[34]) );
  OR3X1_LVT div_sub_x_9_U342 ( .A1(div_result_34_), .A2(div_sub_x_9_n433), 
        .A3(div_sub_x_9_n373), .Y(div_sub_x_9_n434) );
  HADDX1_LVT div_sub_x_9_U341 ( .A0(div_result_35_), .B0(div_sub_x_9_n434), 
        .SO(div_negated_remainder[35]) );
  OR3X1_LVT div_sub_x_9_U340 ( .A1(div_result_35_), .A2(div_result_34_), .A3(
        div_sub_x_9_n433), .Y(div_sub_x_9_n426) );
  OR2X1_LVT div_sub_x_9_U339 ( .A1(div_sub_x_9_n373), .A2(div_sub_x_9_n426), 
        .Y(div_sub_x_9_n430) );
  HADDX1_LVT div_sub_x_9_U338 ( .A0(div_result_36_), .B0(div_sub_x_9_n430), 
        .SO(div_negated_remainder[36]) );
  OR2X1_LVT div_sub_x_9_U337 ( .A1(div_result_36_), .A2(div_sub_x_9_n430), .Y(
        div_sub_x_9_n432) );
  HADDX1_LVT div_sub_x_9_U336 ( .A0(div_sub_x_9_n432), .B0(div_result_37_), 
        .SO(div_negated_remainder[37]) );
  OR2X1_LVT div_sub_x_9_U335 ( .A1(div_result_37_), .A2(div_result_36_), .Y(
        div_sub_x_9_n427) );
  OR3X1_LVT div_sub_x_9_U334 ( .A1(div_sub_x_9_n373), .A2(div_sub_x_9_n426), 
        .A3(div_sub_x_9_n427), .Y(div_sub_x_9_n431) );
  HADDX1_LVT div_sub_x_9_U333 ( .A0(div_result_38_), .B0(div_sub_x_9_n431), 
        .SO(div_negated_remainder[38]) );
  OR3X1_LVT div_sub_x_9_U332 ( .A1(div_result_38_), .A2(div_sub_x_9_n427), 
        .A3(div_sub_x_9_n430), .Y(div_sub_x_9_n429) );
  HADDX1_LVT div_sub_x_9_U331 ( .A0(div_result_39_), .B0(div_sub_x_9_n429), 
        .SO(div_negated_remainder[39]) );
  NAND2X0_LVT div_sub_x_9_U330 ( .A1(div_sub_x_9_n161), .A2(div_sub_x_9_n387), 
        .Y(div_sub_x_9_n428) );
  HADDX1_LVT div_sub_x_9_U329 ( .A0(div_result_3_), .B0(div_sub_x_9_n428), 
        .SO(div_negated_remainder[3]) );
  NAND2X0_LVT div_sub_x_9_U328 ( .A1(div_sub_x_9_n424), .A2(div_sub_x_9_n425), 
        .Y(div_sub_x_9_n422) );
  NAND2X0_LVT div_sub_x_9_U327 ( .A1(div_sub_x_9_n371), .A2(div_sub_x_9_n370), 
        .Y(div_sub_x_9_n423) );
  HADDX1_LVT div_sub_x_9_U326 ( .A0(div_result_41_), .B0(div_sub_x_9_n423), 
        .SO(div_negated_remainder[41]) );
  OR3X1_LVT div_sub_x_9_U325 ( .A1(div_result_41_), .A2(div_result_40_), .A3(
        div_sub_x_9_n422), .Y(div_sub_x_9_n421) );
  HADDX1_LVT div_sub_x_9_U324 ( .A0(div_result_42_), .B0(div_sub_x_9_n421), 
        .SO(div_negated_remainder[42]) );
  OR2X1_LVT div_sub_x_9_U323 ( .A1(div_result_42_), .A2(div_sub_x_9_n421), .Y(
        div_sub_x_9_n420) );
  HADDX1_LVT div_sub_x_9_U322 ( .A0(div_sub_x_9_n420), .B0(div_result_43_), 
        .SO(div_negated_remainder[43]) );
  NAND2X0_LVT div_sub_x_9_U321 ( .A1(div_sub_x_9_n417), .A2(div_sub_x_9_n371), 
        .Y(div_sub_x_9_n415) );
  HADDX1_LVT div_sub_x_9_U320 ( .A0(div_result_44_), .B0(div_sub_x_9_n415), 
        .SO(div_negated_remainder[44]) );
  NAND3X0_LVT div_sub_x_9_U319 ( .A1(div_sub_x_9_n417), .A2(div_sub_x_9_n371), 
        .A3(div_sub_x_9_n369), .Y(div_sub_x_9_n419) );
  HADDX1_LVT div_sub_x_9_U318 ( .A0(div_result_45_), .B0(div_sub_x_9_n419), 
        .SO(div_negated_remainder[45]) );
  OR2X1_LVT div_sub_x_9_U317 ( .A1(div_result_45_), .A2(div_result_44_), .Y(
        div_sub_x_9_n414) );
  NAND3X0_LVT div_sub_x_9_U316 ( .A1(div_sub_x_9_n417), .A2(div_sub_x_9_n368), 
        .A3(div_sub_x_9_n371), .Y(div_sub_x_9_n418) );
  HADDX1_LVT div_sub_x_9_U315 ( .A0(div_result_46_), .B0(div_sub_x_9_n418), 
        .SO(div_negated_remainder[46]) );
  NAND4X0_LVT div_sub_x_9_U314 ( .A1(div_sub_x_9_n368), .A2(div_sub_x_9_n417), 
        .A3(div_sub_x_9_n371), .A4(div_sub_x_9_n367), .Y(div_sub_x_9_n416) );
  HADDX1_LVT div_sub_x_9_U313 ( .A0(div_result_47_), .B0(div_sub_x_9_n416), 
        .SO(div_negated_remainder[47]) );
  NAND2X0_LVT div_sub_x_9_U312 ( .A1(div_sub_x_9_n408), .A2(div_sub_x_9_n365), 
        .Y(div_sub_x_9_n413) );
  HADDX1_LVT div_sub_x_9_U311 ( .A0(div_result_49_), .B0(div_sub_x_9_n413), 
        .SO(div_negated_remainder[49]) );
  OR3X1_LVT div_sub_x_9_U310 ( .A1(div_result_49_), .A2(div_result_48_), .A3(
        div_sub_x_9_n366), .Y(div_sub_x_9_n411) );
  HADDX1_LVT div_sub_x_9_U309 ( .A0(div_result_50_), .B0(div_sub_x_9_n411), 
        .SO(div_negated_remainder[50]) );
  OR2X1_LVT div_sub_x_9_U308 ( .A1(div_result_50_), .A2(div_sub_x_9_n411), .Y(
        div_sub_x_9_n410) );
  HADDX1_LVT div_sub_x_9_U307 ( .A0(div_sub_x_9_n410), .B0(div_result_51_), 
        .SO(div_negated_remainder[51]) );
  NAND2X0_LVT div_sub_x_9_U306 ( .A1(div_sub_x_9_n408), .A2(div_sub_x_9_n409), 
        .Y(div_sub_x_9_n406) );
  NAND2X0_LVT div_sub_x_9_U305 ( .A1(div_sub_x_9_n363), .A2(div_sub_x_9_n364), 
        .Y(div_sub_x_9_n407) );
  HADDX1_LVT div_sub_x_9_U304 ( .A0(div_sub_x_9_n407), .B0(div_result_53_), 
        .SO(div_negated_remainder[53]) );
  OR3X1_LVT div_sub_x_9_U303 ( .A1(div_result_53_), .A2(div_result_52_), .A3(
        div_sub_x_9_n406), .Y(div_sub_x_9_n404) );
  HADDX1_LVT div_sub_x_9_U302 ( .A0(div_result_54_), .B0(div_sub_x_9_n404), 
        .SO(div_negated_remainder[54]) );
  OR2X1_LVT div_sub_x_9_U301 ( .A1(div_result_54_), .A2(div_sub_x_9_n404), .Y(
        div_sub_x_9_n405) );
  HADDX1_LVT div_sub_x_9_U300 ( .A0(div_sub_x_9_n405), .B0(div_result_55_), 
        .SO(div_negated_remainder[55]) );
  OR3X1_LVT div_sub_x_9_U299 ( .A1(div_result_55_), .A2(div_result_54_), .A3(
        div_sub_x_9_n404), .Y(div_sub_x_9_n402) );
  NAND2X0_LVT div_sub_x_9_U298 ( .A1(div_sub_x_9_n361), .A2(div_sub_x_9_n362), 
        .Y(div_sub_x_9_n403) );
  HADDX1_LVT div_sub_x_9_U297 ( .A0(div_sub_x_9_n403), .B0(div_result_57_), 
        .SO(div_negated_remainder[57]) );
  OR3X1_LVT div_sub_x_9_U296 ( .A1(div_result_57_), .A2(div_result_56_), .A3(
        div_sub_x_9_n402), .Y(div_sub_x_9_n399) );
  HADDX1_LVT div_sub_x_9_U295 ( .A0(div_result_58_), .B0(div_sub_x_9_n399), 
        .SO(div_negated_remainder[58]) );
  OR2X1_LVT div_sub_x_9_U294 ( .A1(div_result_58_), .A2(div_sub_x_9_n399), .Y(
        div_sub_x_9_n401) );
  HADDX1_LVT div_sub_x_9_U293 ( .A0(div_result_59_), .B0(div_sub_x_9_n401), 
        .SO(div_negated_remainder[59]) );
  NAND2X0_LVT div_sub_x_9_U292 ( .A1(div_sub_x_9_n385), .A2(div_sub_x_9_n386), 
        .Y(div_sub_x_9_n400) );
  HADDX1_LVT div_sub_x_9_U291 ( .A0(div_sub_x_9_n400), .B0(div_result_5_), 
        .SO(div_negated_remainder[5]) );
  OR3X1_LVT div_sub_x_9_U290 ( .A1(div_result_59_), .A2(div_result_58_), .A3(
        div_sub_x_9_n399), .Y(div_sub_x_9_n397) );
  HADDX1_LVT div_sub_x_9_U289 ( .A0(div_result_60_), .B0(div_sub_x_9_n397), 
        .SO(div_negated_remainder[60]) );
  OR2X1_LVT div_sub_x_9_U288 ( .A1(div_result_60_), .A2(div_sub_x_9_n397), .Y(
        div_sub_x_9_n398) );
  HADDX1_LVT div_sub_x_9_U287 ( .A0(div_result_61_), .B0(div_sub_x_9_n398), 
        .SO(div_negated_remainder[61]) );
  OR3X1_LVT div_sub_x_9_U286 ( .A1(div_result_61_), .A2(div_result_60_), .A3(
        div_sub_x_9_n397), .Y(div_sub_x_9_n396) );
  HADDX1_LVT div_sub_x_9_U285 ( .A0(div_result_62_), .B0(div_sub_x_9_n396), 
        .SO(div_negated_remainder[62]) );
  OR2X1_LVT div_sub_x_9_U284 ( .A1(div_result_62_), .A2(div_sub_x_9_n396), .Y(
        div_sub_x_9_n395) );
  HADDX1_LVT div_sub_x_9_U283 ( .A0(div_sub_x_9_n395), .B0(div_result_63_), 
        .SO(div_negated_remainder[63]) );
  HADDX1_LVT div_sub_x_9_U282 ( .A0(div_result_6_), .B0(div_sub_x_9_n394), 
        .SO(div_negated_remainder[6]) );
  OR2X1_LVT div_sub_x_9_U281 ( .A1(div_result_6_), .A2(div_sub_x_9_n394), .Y(
        div_sub_x_9_n393) );
  HADDX1_LVT div_sub_x_9_U280 ( .A0(div_result_7_), .B0(div_sub_x_9_n393), 
        .SO(div_negated_remainder[7]) );
  AO22X1_LVT div_sub_x_9_U279 ( .A1(div_sub_x_9_n384), .A2(div_result_8_), 
        .A3(div_sub_x_9_n392), .A4(div_sub_x_9_n383), .Y(
        div_negated_remainder[8]) );
  NAND2X0_LVT div_sub_x_9_U278 ( .A1(div_sub_x_9_n384), .A2(div_sub_x_9_n383), 
        .Y(div_sub_x_9_n391) );
  HADDX1_LVT div_sub_x_9_U277 ( .A0(div_result_9_), .B0(div_sub_x_9_n391), 
        .SO(div_negated_remainder[9]) );
  INVX1_LVT div_sub_x_9_U276 ( .A(div_sub_x_9_n161), .Y(div_sub_x_9_n388) );
  INVX1_LVT div_sub_x_9_U275 ( .A(div_sub_x_9_n412), .Y(div_sub_x_9_n386) );
  INVX1_LVT div_sub_x_9_U274 ( .A(div_sub_x_9_n392), .Y(div_sub_x_9_n384) );
  INVX1_LVT div_sub_x_9_U273 ( .A(div_sub_x_9_n453), .Y(div_sub_x_9_n380) );
  INVX1_LVT div_sub_x_9_U272 ( .A(div_sub_x_9_n445), .Y(div_sub_x_9_n378) );
  INVX1_LVT div_sub_x_9_U271 ( .A(div_sub_x_9_n437), .Y(div_sub_x_9_n375) );
  INVX1_LVT div_sub_x_9_U270 ( .A(div_sub_x_9_n424), .Y(div_sub_x_9_n373) );
  INVX1_LVT div_sub_x_9_U269 ( .A(div_sub_x_9_n422), .Y(div_sub_x_9_n371) );
  INVX1_LVT div_sub_x_9_U268 ( .A(div_sub_x_9_n414), .Y(div_sub_x_9_n368) );
  INVX1_LVT div_sub_x_9_U267 ( .A(div_sub_x_9_n408), .Y(div_sub_x_9_n366) );
  INVX1_LVT div_sub_x_9_U266 ( .A(div_sub_x_9_n402), .Y(div_sub_x_9_n362) );
  NOR4X1_LVT div_sub_x_9_U265 ( .A1(div_result_41_), .A2(div_result_40_), .A3(
        div_result_43_), .A4(div_result_42_), .Y(div_sub_x_9_n417) );
  NOR4X1_LVT div_sub_x_9_U264 ( .A1(div_result_25_), .A2(div_result_24_), .A3(
        div_result_27_), .A4(div_result_26_), .Y(div_sub_x_9_n440) );
  NOR4X1_LVT div_sub_x_9_U263 ( .A1(div_result_22_), .A2(div_result_23_), .A3(
        div_sub_x_9_n448), .A4(div_sub_x_9_n449), .Y(div_sub_x_9_n447) );
  NOR4X1_LVT div_sub_x_9_U262 ( .A1(div_result_30_), .A2(div_result_31_), .A3(
        div_sub_x_9_n437), .A4(div_sub_x_9_n438), .Y(div_sub_x_9_n424) );
  NOR4X1_LVT div_sub_x_9_U261 ( .A1(div_result_38_), .A2(div_result_39_), .A3(
        div_sub_x_9_n426), .A4(div_sub_x_9_n427), .Y(div_sub_x_9_n425) );
  NOR4X1_LVT div_sub_x_9_U260 ( .A1(div_result_46_), .A2(div_result_47_), .A3(
        div_sub_x_9_n414), .A4(div_sub_x_9_n415), .Y(div_sub_x_9_n408) );
  NOR4X1_LVT div_sub_x_9_U259 ( .A1(div_result_49_), .A2(div_result_48_), .A3(
        div_result_51_), .A4(div_result_50_), .Y(div_sub_x_9_n409) );
  INVX0_LVT div_sub_x_9_U258 ( .A(div_result_30_), .Y(div_sub_x_9_n374) );
  INVX0_LVT div_sub_x_9_U257 ( .A(div_result_32_), .Y(div_sub_x_9_n372) );
  INVX0_LVT div_sub_x_9_U256 ( .A(div_result_24_), .Y(div_sub_x_9_n377) );
  INVX0_LVT div_sub_x_9_U255 ( .A(div_result_28_), .Y(div_sub_x_9_n376) );
  INVX0_LVT div_sub_x_9_U254 ( .A(div_result_4_), .Y(div_sub_x_9_n385) );
  INVX0_LVT div_sub_x_9_U253 ( .A(div_result_48_), .Y(div_sub_x_9_n365) );
  INVX0_LVT div_sub_x_9_U252 ( .A(div_result_46_), .Y(div_sub_x_9_n367) );
  INVX0_LVT div_sub_x_9_U251 ( .A(div_result_44_), .Y(div_sub_x_9_n369) );
  INVX0_LVT div_sub_x_9_U250 ( .A(div_result_12_), .Y(div_sub_x_9_n381) );
  INVX0_LVT div_sub_x_9_U249 ( .A(div_result_52_), .Y(div_sub_x_9_n363) );
  INVX0_LVT div_sub_x_9_U248 ( .A(div_result_56_), .Y(div_sub_x_9_n361) );
  INVX0_LVT div_sub_x_9_U247 ( .A(div_result_8_), .Y(div_sub_x_9_n383) );
  INVX0_LVT div_sub_x_9_U246 ( .A(div_result_40_), .Y(div_sub_x_9_n370) );
  INVX0_LVT div_sub_x_9_U245 ( .A(div_result_16_), .Y(div_sub_x_9_n379) );
  INVX0_LVT div_sub_x_9_U244 ( .A(div_result_1_), .Y(div_sub_x_9_n389) );
  INVX0_LVT div_sub_x_9_U243 ( .A(div_result_0_), .Y(div_sub_x_9_n390) );
  INVX0_LVT div_sub_x_9_U242 ( .A(div_result_2_), .Y(div_sub_x_9_n387) );
  INVX0_LVT div_sub_x_9_U241 ( .A(div_sub_x_9_n461), .Y(div_sub_x_9_n382) );
  INVX0_LVT div_sub_x_9_U240 ( .A(div_sub_x_9_n406), .Y(div_sub_x_9_n364) );
  NOR4X1_LVT div_sub_x_9_U239 ( .A1(div_result_9_), .A2(div_result_8_), .A3(
        div_result_11_), .A4(div_result_10_), .Y(div_sub_x_9_n463) );
  AO22X1_LVT div_sub_x_9_U238 ( .A1(div_result_52_), .A2(div_sub_x_9_n364), 
        .A3(div_sub_x_9_n406), .A4(div_sub_x_9_n363), .Y(
        div_negated_remainder[52]) );
  AO22X1_LVT div_sub_x_9_U237 ( .A1(div_result_32_), .A2(div_sub_x_9_n424), 
        .A3(div_sub_x_9_n372), .A4(div_sub_x_9_n373), .Y(
        div_negated_remainder[32]) );
  AO22X1_LVT div_sub_x_9_U236 ( .A1(div_result_4_), .A2(div_sub_x_9_n386), 
        .A3(div_sub_x_9_n412), .A4(div_sub_x_9_n385), .Y(
        div_negated_remainder[4]) );
  AO22X1_LVT div_sub_x_9_U235 ( .A1(div_result_16_), .A2(div_sub_x_9_n380), 
        .A3(div_sub_x_9_n453), .A4(div_sub_x_9_n379), .Y(
        div_negated_remainder[16]) );
  AO22X1_LVT div_sub_x_9_U234 ( .A1(div_result_2_), .A2(div_sub_x_9_n161), 
        .A3(div_sub_x_9_n387), .A4(div_sub_x_9_n388), .Y(
        div_negated_remainder[2]) );
  AO22X1_LVT div_sub_x_9_U233 ( .A1(div_result_24_), .A2(div_sub_x_9_n378), 
        .A3(div_sub_x_9_n445), .A4(div_sub_x_9_n377), .Y(
        div_negated_remainder[24]) );
  AO22X1_LVT div_sub_x_9_U232 ( .A1(div_result_40_), .A2(div_sub_x_9_n371), 
        .A3(div_sub_x_9_n422), .A4(div_sub_x_9_n370), .Y(
        div_negated_remainder[40]) );
  AO22X1_LVT div_sub_x_9_U231 ( .A1(div_sub_x_9_n461), .A2(div_sub_x_9_n381), 
        .A3(div_sub_x_9_n382), .A4(div_result_12_), .Y(
        div_negated_remainder[12]) );
  AO22X1_LVT div_sub_x_9_U230 ( .A1(div_result_48_), .A2(div_sub_x_9_n408), 
        .A3(div_sub_x_9_n365), .A4(div_sub_x_9_n366), .Y(
        div_negated_remainder[48]) );
  AO22X1_LVT div_sub_x_9_U229 ( .A1(div_result_56_), .A2(div_sub_x_9_n362), 
        .A3(div_sub_x_9_n402), .A4(div_sub_x_9_n361), .Y(
        div_negated_remainder[56]) );
  HADDX1_LVT div_sub_x_9_U223 ( .A0(div_sub_x_9_n389), .B0(div_sub_x_9_n390), 
        .C1(div_sub_x_9_n161), .SO(div_negated_remainder[1]) );
  AO22X1_LVT div_sub_x_7_U1048 ( .A1(div_n301), .A2(div_sub_x_7_n877), .A3(
        div_sub_x_7_n833), .A4(div_divisor_0_), .Y(div_subtractor_0_) );
  NOR2X0_LVT div_sub_x_7_U1047 ( .A1(div_sub_x_7_n901), .A2(div_divisor_9_), 
        .Y(div_sub_x_7_n1104) );
  OR2X1_LVT div_sub_x_7_U1046 ( .A1(div_sub_x_7_n871), .A2(div_n_T_51_71_), 
        .Y(div_sub_x_7_n1109) );
  AO22X1_LVT div_sub_x_7_U1045 ( .A1(div_n_T_51_71_), .A2(div_sub_x_7_n871), 
        .A3(div_sub_x_7_n911), .A4(div_sub_x_7_n1109), .Y(div_sub_x_7_n1107)
         );
  NAND2X0_LVT div_sub_x_7_U1044 ( .A1(div_divisor_7_), .A2(div_sub_x_7_n902), 
        .Y(div_sub_x_7_n910) );
  NAND2X0_LVT div_sub_x_7_U1043 ( .A1(div_divisor_6_), .A2(div_sub_x_7_n903), 
        .Y(div_sub_x_7_n1116) );
  OR2X1_LVT div_sub_x_7_U1042 ( .A1(div_sub_x_7_n873), .A2(div_n_T_51_68_), 
        .Y(div_sub_x_7_n915) );
  NAND2X0_LVT div_sub_x_7_U1041 ( .A1(div_sub_x_7_n1116), .A2(div_sub_x_7_n915), .Y(div_sub_x_7_n1111) );
  NAND2X0_LVT div_sub_x_7_U1040 ( .A1(div_n_T_51_66_), .A2(div_sub_x_7_n874), 
        .Y(div_sub_x_7_n976) );
  AO222X1_LVT div_sub_x_7_U1039 ( .A1(div_divisor_4_), .A2(div_sub_x_7_n904), 
        .A3(div_divisor_4_), .A4(div_sub_x_7_n976), .A5(div_sub_x_7_n904), 
        .A6(div_sub_x_7_n976), .Y(div_sub_x_7_n934) );
  NAND2X0_LVT div_sub_x_7_U1038 ( .A1(div_divisor_4_), .A2(div_sub_x_7_n904), 
        .Y(div_sub_x_7_n1114) );
  NAND2X0_LVT div_sub_x_7_U1037 ( .A1(div_divisor_1_), .A2(div_sub_x_7_n907), 
        .Y(div_sub_x_7_n1050) );
  NAND2X0_LVT div_sub_x_7_U1036 ( .A1(div_divisor_0_), .A2(div_sub_x_7_n833), 
        .Y(div_sub_x_7_n1049) );
  NAND2X0_LVT div_sub_x_7_U1035 ( .A1(div_divisor_3_), .A2(div_sub_x_7_n905), 
        .Y(div_sub_x_7_n1115) );
  NAND3X0_LVT div_sub_x_7_U1034 ( .A1(div_sub_x_7_n1114), .A2(div_sub_x_7_n977), .A3(div_sub_x_7_n1115), .Y(div_sub_x_7_n935) );
  NAND2X0_LVT div_sub_x_7_U1033 ( .A1(div_n_T_51_68_), .A2(div_sub_x_7_n873), 
        .Y(div_sub_x_7_n1113) );
  AO222X1_LVT div_sub_x_7_U1032 ( .A1(div_divisor_6_), .A2(div_sub_x_7_n903), 
        .A3(div_divisor_6_), .A4(div_sub_x_7_n1113), .A5(div_sub_x_7_n903), 
        .A6(div_sub_x_7_n1113), .Y(div_sub_x_7_n1112) );
  OA221X1_LVT div_sub_x_7_U1031 ( .A1(div_sub_x_7_n1111), .A2(div_sub_x_7_n934), .A3(div_sub_x_7_n1111), .A4(div_sub_x_7_n935), .A5(div_sub_x_7_n1112), .Y(
        div_sub_x_7_n912) );
  OA222X1_LVT div_sub_x_7_U1030 ( .A1(div_sub_x_7_n1107), .A2(
        div_sub_x_7_n1109), .A3(div_sub_x_7_n1107), .A4(div_sub_x_7_n910), 
        .A5(div_sub_x_7_n1107), .A6(div_sub_x_7_n872), .Y(div_sub_x_7_n908) );
  NAND2X0_LVT div_sub_x_7_U1029 ( .A1(div_divisor_9_), .A2(div_sub_x_7_n901), 
        .Y(div_sub_x_7_n1108) );
  OA21X1_LVT div_sub_x_7_U1028 ( .A1(div_sub_x_7_n1104), .A2(div_sub_x_7_n908), 
        .A3(div_sub_x_7_n1108), .Y(div_sub_x_7_n1110) );
  FADDX1_LVT div_sub_x_7_U1027 ( .A(div_n_T_51_73_), .B(div_sub_x_7_n1110), 
        .CI(div_sub_x_7_n870), .S(div_subtractor_10_) );
  OR2X1_LVT div_sub_x_7_U1026 ( .A1(div_sub_x_7_n870), .A2(div_n_T_51_73_), 
        .Y(div_sub_x_7_n1105) );
  AND4X1_LVT div_sub_x_7_U1025 ( .A1(div_sub_x_7_n1109), .A2(div_sub_x_7_n910), 
        .A3(div_sub_x_7_n1108), .A4(div_sub_x_7_n1105), .Y(div_sub_x_7_n1092)
         );
  AND2X1_LVT div_sub_x_7_U1024 ( .A1(div_sub_x_7_n1108), .A2(div_sub_x_7_n1105), .Y(div_sub_x_7_n1106) );
  AO222X1_LVT div_sub_x_7_U1023 ( .A1(div_n_T_51_73_), .A2(div_sub_x_7_n870), 
        .A3(div_sub_x_7_n1104), .A4(div_sub_x_7_n1105), .A5(div_sub_x_7_n1106), 
        .A6(div_sub_x_7_n1107), .Y(div_sub_x_7_n1094) );
  AO21X1_LVT div_sub_x_7_U1022 ( .A1(div_sub_x_7_n1092), .A2(div_sub_x_7_n872), 
        .A3(div_sub_x_7_n1094), .Y(div_sub_x_7_n1101) );
  FADDX1_LVT div_sub_x_7_U1021 ( .A(div_n_T_51_74_), .B(div_sub_x_7_n869), 
        .CI(div_sub_x_7_n1101), .S(div_subtractor_11_) );
  NAND2X0_LVT div_sub_x_7_U1020 ( .A1(div_n_T_51_74_), .A2(div_sub_x_7_n869), 
        .Y(div_sub_x_7_n1102) );
  OR2X1_LVT div_sub_x_7_U1019 ( .A1(div_sub_x_7_n869), .A2(div_n_T_51_74_), 
        .Y(div_sub_x_7_n1096) );
  OA21X1_LVT div_sub_x_7_U1018 ( .A1(div_sub_x_7_n868), .A2(div_sub_x_7_n1101), 
        .A3(div_sub_x_7_n1096), .Y(div_sub_x_7_n1103) );
  FADDX1_LVT div_sub_x_7_U1017 ( .A(div_divisor_12_), .B(div_sub_x_7_n1103), 
        .CI(div_sub_x_7_n900), .S(div_subtractor_12_) );
  AO222X1_LVT div_sub_x_7_U1016 ( .A1(div_divisor_12_), .A2(div_sub_x_7_n900), 
        .A3(div_divisor_12_), .A4(div_sub_x_7_n1102), .A5(div_sub_x_7_n900), 
        .A6(div_sub_x_7_n1102), .Y(div_sub_x_7_n1093) );
  NAND2X0_LVT div_sub_x_7_U1015 ( .A1(div_divisor_12_), .A2(div_sub_x_7_n900), 
        .Y(div_sub_x_7_n1095) );
  NAND3X0_LVT div_sub_x_7_U1014 ( .A1(div_sub_x_7_n1101), .A2(
        div_sub_x_7_n1095), .A3(div_sub_x_7_n1096), .Y(div_sub_x_7_n1100) );
  AND2X1_LVT div_sub_x_7_U1013 ( .A1(div_sub_x_7_n1093), .A2(div_sub_x_7_n1100), .Y(div_sub_x_7_n1099) );
  FADDX1_LVT div_sub_x_7_U1012 ( .A(div_n_T_51_76_), .B(div_divisor_13_), .CI(
        div_sub_x_7_n1099), .S(div_subtractor_13_) );
  OR2X1_LVT div_sub_x_7_U1011 ( .A1(div_sub_x_7_n899), .A2(div_divisor_13_), 
        .Y(div_sub_x_7_n1097) );
  AO22X1_LVT div_sub_x_7_U1010 ( .A1(div_sub_x_7_n1099), .A2(div_sub_x_7_n1097), .A3(div_divisor_13_), .A4(div_sub_x_7_n899), .Y(div_sub_x_7_n1098) );
  FADDX1_LVT div_sub_x_7_U1009 ( .A(div_n_T_51_77_), .B(div_divisor_14_), .CI(
        div_sub_x_7_n1098), .S(div_subtractor_14_) );
  FADDX1_LVT div_sub_x_7_U1008 ( .A(div_sub_x_7_n1041), .B(div_n_T_51_78_), 
        .CI(div_sub_x_7_n867), .S(div_subtractor_15_) );
  AND2X1_LVT div_sub_x_7_U1007 ( .A1(div_n_T_51_78_), .A2(div_sub_x_7_n867), 
        .Y(div_sub_x_7_n1090) );
  OR2X1_LVT div_sub_x_7_U1006 ( .A1(div_sub_x_7_n867), .A2(div_n_T_51_78_), 
        .Y(div_sub_x_7_n1087) );
  OA21X1_LVT div_sub_x_7_U1005 ( .A1(div_sub_x_7_n1041), .A2(div_sub_x_7_n1090), .A3(div_sub_x_7_n1087), .Y(div_sub_x_7_n1091) );
  FADDX1_LVT div_sub_x_7_U1004 ( .A(div_n_T_51_79_), .B(div_sub_x_7_n1091), 
        .CI(div_sub_x_7_n866), .S(div_subtractor_16_) );
  OR2X1_LVT div_sub_x_7_U1003 ( .A1(div_sub_x_7_n866), .A2(div_n_T_51_79_), 
        .Y(div_sub_x_7_n1086) );
  AO22X1_LVT div_sub_x_7_U1002 ( .A1(div_n_T_51_79_), .A2(div_sub_x_7_n866), 
        .A3(div_sub_x_7_n1090), .A4(div_sub_x_7_n1086), .Y(div_sub_x_7_n1084)
         );
  OA222X1_LVT div_sub_x_7_U1001 ( .A1(div_sub_x_7_n1084), .A2(
        div_sub_x_7_n1041), .A3(div_sub_x_7_n1084), .A4(div_sub_x_7_n1086), 
        .A5(div_sub_x_7_n1084), .A6(div_sub_x_7_n1087), .Y(div_sub_x_7_n1089)
         );
  FADDX1_LVT div_sub_x_7_U1000 ( .A(div_n_T_51_80_), .B(div_sub_x_7_n1089), 
        .CI(div_sub_x_7_n865), .S(div_subtractor_17_) );
  OR2X1_LVT div_sub_x_7_U999 ( .A1(div_sub_x_7_n865), .A2(div_n_T_51_80_), .Y(
        div_sub_x_7_n1085) );
  AND2X1_LVT div_sub_x_7_U998 ( .A1(div_n_T_51_80_), .A2(div_sub_x_7_n865), 
        .Y(div_sub_x_7_n1081) );
  AO21X1_LVT div_sub_x_7_U997 ( .A1(div_sub_x_7_n1089), .A2(div_sub_x_7_n1085), 
        .A3(div_sub_x_7_n1081), .Y(div_sub_x_7_n1088) );
  FADDX1_LVT div_sub_x_7_U996 ( .A(div_n_T_51_81_), .B(div_sub_x_7_n864), .CI(
        div_sub_x_7_n1088), .S(div_subtractor_18_) );
  OR2X1_LVT div_sub_x_7_U995 ( .A1(div_sub_x_7_n864), .A2(div_n_T_51_81_), .Y(
        div_sub_x_7_n1082) );
  AND4X1_LVT div_sub_x_7_U994 ( .A1(div_sub_x_7_n1082), .A2(div_sub_x_7_n1085), 
        .A3(div_sub_x_7_n1086), .A4(div_sub_x_7_n1087), .Y(div_sub_x_7_n1072)
         );
  AND2X1_LVT div_sub_x_7_U993 ( .A1(div_sub_x_7_n1082), .A2(div_sub_x_7_n1085), 
        .Y(div_sub_x_7_n1083) );
  AO222X1_LVT div_sub_x_7_U992 ( .A1(div_n_T_51_81_), .A2(div_sub_x_7_n864), 
        .A3(div_sub_x_7_n1081), .A4(div_sub_x_7_n1082), .A5(div_sub_x_7_n1083), 
        .A6(div_sub_x_7_n1084), .Y(div_sub_x_7_n1069) );
  AO21X1_LVT div_sub_x_7_U991 ( .A1(div_sub_x_7_n1041), .A2(div_sub_x_7_n1072), 
        .A3(div_sub_x_7_n1069), .Y(div_sub_x_7_n1078) );
  FADDX1_LVT div_sub_x_7_U990 ( .A(div_n_T_51_82_), .B(div_sub_x_7_n1078), 
        .CI(div_sub_x_7_n863), .S(div_subtractor_19_) );
  FADDX1_LVT div_sub_x_7_U989 ( .A(div_divisor_1_), .B(div_sub_x_7_n907), .CI(
        div_sub_x_7_n1049), .S(div_subtractor_1_) );
  OR2X1_LVT div_sub_x_7_U988 ( .A1(div_sub_x_7_n863), .A2(div_n_T_51_82_), .Y(
        div_sub_x_7_n1074) );
  AO22X1_LVT div_sub_x_7_U987 ( .A1(div_n_T_51_82_), .A2(div_sub_x_7_n863), 
        .A3(div_sub_x_7_n1078), .A4(div_sub_x_7_n1074), .Y(div_sub_x_7_n1080)
         );
  FADDX1_LVT div_sub_x_7_U986 ( .A(div_divisor_20_), .B(div_sub_x_7_n898), 
        .CI(div_sub_x_7_n1080), .S(div_subtractor_20_) );
  NAND2X0_LVT div_sub_x_7_U985 ( .A1(div_n_T_51_82_), .A2(div_sub_x_7_n863), 
        .Y(div_sub_x_7_n1079) );
  AO222X1_LVT div_sub_x_7_U984 ( .A1(div_divisor_20_), .A2(div_sub_x_7_n898), 
        .A3(div_divisor_20_), .A4(div_sub_x_7_n1079), .A5(div_sub_x_7_n898), 
        .A6(div_sub_x_7_n1079), .Y(div_sub_x_7_n1067) );
  NAND2X0_LVT div_sub_x_7_U983 ( .A1(div_divisor_20_), .A2(div_sub_x_7_n898), 
        .Y(div_sub_x_7_n1073) );
  NAND3X0_LVT div_sub_x_7_U982 ( .A1(div_sub_x_7_n1073), .A2(div_sub_x_7_n1078), .A3(div_sub_x_7_n1074), .Y(div_sub_x_7_n1077) );
  NAND2X0_LVT div_sub_x_7_U981 ( .A1(div_sub_x_7_n1067), .A2(div_sub_x_7_n1077), .Y(div_sub_x_7_n1076) );
  FADDX1_LVT div_sub_x_7_U980 ( .A(div_n_T_51_84_), .B(div_sub_x_7_n1076), 
        .CI(div_sub_x_7_n862), .S(div_subtractor_21_) );
  OR2X1_LVT div_sub_x_7_U979 ( .A1(div_sub_x_7_n862), .A2(div_n_T_51_84_), .Y(
        div_sub_x_7_n1071) );
  AO22X1_LVT div_sub_x_7_U978 ( .A1(div_n_T_51_84_), .A2(div_sub_x_7_n862), 
        .A3(div_sub_x_7_n1076), .A4(div_sub_x_7_n1071), .Y(div_sub_x_7_n1075)
         );
  FADDX1_LVT div_sub_x_7_U977 ( .A(div_divisor_22_), .B(div_sub_x_7_n897), 
        .CI(div_sub_x_7_n1075), .S(div_subtractor_22_) );
  NAND2X0_LVT div_sub_x_7_U976 ( .A1(div_divisor_22_), .A2(div_sub_x_7_n897), 
        .Y(div_sub_x_7_n1070) );
  AND4X1_LVT div_sub_x_7_U975 ( .A1(div_sub_x_7_n1070), .A2(div_sub_x_7_n1071), 
        .A3(div_sub_x_7_n1073), .A4(div_sub_x_7_n1074), .Y(div_sub_x_7_n1068)
         );
  AND2X1_LVT div_sub_x_7_U974 ( .A1(div_sub_x_7_n1072), .A2(div_sub_x_7_n1068), 
        .Y(div_sub_x_7_n1042) );
  FADDX1_LVT div_sub_x_7_U973 ( .A(div_n_T_51_86_), .B(div_sub_x_7_n1055), 
        .CI(div_sub_x_7_n861), .S(div_subtractor_23_) );
  OR2X1_LVT div_sub_x_7_U972 ( .A1(div_sub_x_7_n861), .A2(div_n_T_51_86_), .Y(
        div_sub_x_7_n1062) );
  AND2X1_LVT div_sub_x_7_U971 ( .A1(div_n_T_51_86_), .A2(div_sub_x_7_n861), 
        .Y(div_sub_x_7_n1065) );
  AO21X1_LVT div_sub_x_7_U970 ( .A1(div_sub_x_7_n1055), .A2(div_sub_x_7_n1062), 
        .A3(div_sub_x_7_n1065), .Y(div_sub_x_7_n1066) );
  FADDX1_LVT div_sub_x_7_U969 ( .A(div_n_T_51_87_), .B(div_sub_x_7_n860), .CI(
        div_sub_x_7_n1066), .S(div_subtractor_24_) );
  OR2X1_LVT div_sub_x_7_U968 ( .A1(div_sub_x_7_n860), .A2(div_n_T_51_87_), .Y(
        div_sub_x_7_n1061) );
  AO22X1_LVT div_sub_x_7_U967 ( .A1(div_n_T_51_87_), .A2(div_sub_x_7_n860), 
        .A3(div_sub_x_7_n1065), .A4(div_sub_x_7_n1061), .Y(div_sub_x_7_n1059)
         );
  OA222X1_LVT div_sub_x_7_U966 ( .A1(div_sub_x_7_n1059), .A2(div_sub_x_7_n1055), .A3(div_sub_x_7_n1059), .A4(div_sub_x_7_n1061), .A5(div_sub_x_7_n1059), .A6(
        div_sub_x_7_n1062), .Y(div_sub_x_7_n1064) );
  FADDX1_LVT div_sub_x_7_U965 ( .A(div_n_T_51_88_), .B(div_sub_x_7_n1064), 
        .CI(div_sub_x_7_n859), .S(div_subtractor_25_) );
  OR2X1_LVT div_sub_x_7_U964 ( .A1(div_sub_x_7_n859), .A2(div_n_T_51_88_), .Y(
        div_sub_x_7_n1060) );
  AND2X1_LVT div_sub_x_7_U963 ( .A1(div_n_T_51_88_), .A2(div_sub_x_7_n859), 
        .Y(div_sub_x_7_n1056) );
  AO21X1_LVT div_sub_x_7_U962 ( .A1(div_sub_x_7_n1064), .A2(div_sub_x_7_n1060), 
        .A3(div_sub_x_7_n1056), .Y(div_sub_x_7_n1063) );
  FADDX1_LVT div_sub_x_7_U961 ( .A(div_n_T_51_89_), .B(div_sub_x_7_n858), .CI(
        div_sub_x_7_n1063), .S(div_subtractor_26_) );
  OR2X1_LVT div_sub_x_7_U960 ( .A1(div_sub_x_7_n858), .A2(div_n_T_51_89_), .Y(
        div_sub_x_7_n1057) );
  AND4X1_LVT div_sub_x_7_U959 ( .A1(div_sub_x_7_n1057), .A2(div_sub_x_7_n1060), 
        .A3(div_sub_x_7_n1061), .A4(div_sub_x_7_n1062), .Y(div_sub_x_7_n1043)
         );
  AND2X1_LVT div_sub_x_7_U958 ( .A1(div_sub_x_7_n1057), .A2(div_sub_x_7_n1060), 
        .Y(div_sub_x_7_n1058) );
  AO222X1_LVT div_sub_x_7_U957 ( .A1(div_n_T_51_89_), .A2(div_sub_x_7_n858), 
        .A3(div_sub_x_7_n1056), .A4(div_sub_x_7_n1057), .A5(div_sub_x_7_n1058), 
        .A6(div_sub_x_7_n1059), .Y(div_sub_x_7_n1039) );
  AO21X1_LVT div_sub_x_7_U956 ( .A1(div_sub_x_7_n1043), .A2(div_sub_x_7_n1055), 
        .A3(div_sub_x_7_n1039), .Y(div_sub_x_7_n1052) );
  FADDX1_LVT div_sub_x_7_U955 ( .A(div_n_T_51_90_), .B(div_sub_x_7_n1052), 
        .CI(div_sub_x_7_n857), .S(div_subtractor_27_) );
  OR2X1_LVT div_sub_x_7_U954 ( .A1(div_sub_x_7_n857), .A2(div_n_T_51_90_), .Y(
        div_sub_x_7_n1045) );
  AO22X1_LVT div_sub_x_7_U953 ( .A1(div_n_T_51_90_), .A2(div_sub_x_7_n857), 
        .A3(div_sub_x_7_n1052), .A4(div_sub_x_7_n1045), .Y(div_sub_x_7_n1054)
         );
  FADDX1_LVT div_sub_x_7_U952 ( .A(div_divisor_28_), .B(div_sub_x_7_n896), 
        .CI(div_sub_x_7_n1054), .S(div_subtractor_28_) );
  NAND2X0_LVT div_sub_x_7_U951 ( .A1(div_n_T_51_90_), .A2(div_sub_x_7_n857), 
        .Y(div_sub_x_7_n1053) );
  AO222X1_LVT div_sub_x_7_U950 ( .A1(div_divisor_28_), .A2(div_sub_x_7_n896), 
        .A3(div_divisor_28_), .A4(div_sub_x_7_n1053), .A5(div_sub_x_7_n896), 
        .A6(div_sub_x_7_n1053), .Y(div_sub_x_7_n1038) );
  NAND2X0_LVT div_sub_x_7_U949 ( .A1(div_divisor_28_), .A2(div_sub_x_7_n896), 
        .Y(div_sub_x_7_n1044) );
  NAND3X0_LVT div_sub_x_7_U948 ( .A1(div_sub_x_7_n1044), .A2(div_sub_x_7_n1052), .A3(div_sub_x_7_n1045), .Y(div_sub_x_7_n1051) );
  NAND2X0_LVT div_sub_x_7_U947 ( .A1(div_sub_x_7_n1038), .A2(div_sub_x_7_n1051), .Y(div_sub_x_7_n1047) );
  FADDX1_LVT div_sub_x_7_U946 ( .A(div_n_T_51_92_), .B(div_sub_x_7_n1047), 
        .CI(div_sub_x_7_n856), .S(div_subtractor_29_) );
  AO22X1_LVT div_sub_x_7_U945 ( .A1(div_n_T_51_64_), .A2(div_sub_x_7_n876), 
        .A3(div_sub_x_7_n1049), .A4(div_sub_x_7_n1050), .Y(div_sub_x_7_n1048)
         );
  FADDX1_LVT div_sub_x_7_U944 ( .A(div_divisor_2_), .B(div_sub_x_7_n906), .CI(
        div_sub_x_7_n1048), .S(div_subtractor_2_) );
  OR2X1_LVT div_sub_x_7_U943 ( .A1(div_sub_x_7_n856), .A2(div_n_T_51_92_), .Y(
        div_sub_x_7_n1040) );
  AO22X1_LVT div_sub_x_7_U942 ( .A1(div_n_T_51_92_), .A2(div_sub_x_7_n856), 
        .A3(div_sub_x_7_n1047), .A4(div_sub_x_7_n1040), .Y(div_sub_x_7_n1046)
         );
  FADDX1_LVT div_sub_x_7_U941 ( .A(div_divisor_30_), .B(div_sub_x_7_n895), 
        .CI(div_sub_x_7_n1046), .S(div_subtractor_30_) );
  FADDX1_LVT div_sub_x_7_U940 ( .A(div_n_T_51_94_), .B(div_divisor_31_), .CI(
        div_sub_x_7_n918), .S(div_subtractor_31_) );
  NAND2X0_LVT div_sub_x_7_U939 ( .A1(div_divisor_31_), .A2(div_sub_x_7_n894), 
        .Y(div_sub_x_7_n1032) );
  AO21X1_LVT div_sub_x_7_U938 ( .A1(div_sub_x_7_n1032), .A2(div_sub_x_7_n834), 
        .A3(div_sub_x_7_n1035), .Y(div_sub_x_7_n1036) );
  FADDX1_LVT div_sub_x_7_U937 ( .A(div_n_T_51_95_), .B(div_sub_x_7_n855), .CI(
        div_sub_x_7_n1036), .S(div_subtractor_32_) );
  OR2X1_LVT div_sub_x_7_U936 ( .A1(div_sub_x_7_n855), .A2(div_n_T_51_95_), .Y(
        div_sub_x_7_n1031) );
  AO22X1_LVT div_sub_x_7_U935 ( .A1(div_n_T_51_95_), .A2(div_sub_x_7_n855), 
        .A3(div_sub_x_7_n1035), .A4(div_sub_x_7_n1031), .Y(div_sub_x_7_n1029)
         );
  OA222X1_LVT div_sub_x_7_U934 ( .A1(div_sub_x_7_n1029), .A2(div_sub_x_7_n1031), .A3(div_sub_x_7_n1029), .A4(div_sub_x_7_n1032), .A5(div_sub_x_7_n1029), .A6(
        div_sub_x_7_n834), .Y(div_sub_x_7_n1034) );
  FADDX1_LVT div_sub_x_7_U933 ( .A(div_n_T_51_96_), .B(div_sub_x_7_n854), .CI(
        div_sub_x_7_n1034), .S(div_subtractor_33_) );
  AND2X1_LVT div_sub_x_7_U932 ( .A1(div_n_T_51_96_), .A2(div_sub_x_7_n854), 
        .Y(div_sub_x_7_n1026) );
  OR2X1_LVT div_sub_x_7_U931 ( .A1(div_sub_x_7_n854), .A2(div_n_T_51_96_), .Y(
        div_sub_x_7_n1030) );
  OA21X1_LVT div_sub_x_7_U930 ( .A1(div_sub_x_7_n1026), .A2(div_sub_x_7_n1034), 
        .A3(div_sub_x_7_n1030), .Y(div_sub_x_7_n1033) );
  FADDX1_LVT div_sub_x_7_U929 ( .A(div_n_T_51_97_), .B(div_sub_x_7_n1033), 
        .CI(div_sub_x_7_n853), .S(div_subtractor_34_) );
  OR2X1_LVT div_sub_x_7_U928 ( .A1(div_sub_x_7_n853), .A2(div_n_T_51_97_), .Y(
        div_sub_x_7_n1027) );
  AND4X1_LVT div_sub_x_7_U927 ( .A1(div_sub_x_7_n1027), .A2(div_sub_x_7_n1030), 
        .A3(div_sub_x_7_n1031), .A4(div_sub_x_7_n1032), .Y(div_sub_x_7_n1012)
         );
  AND2X1_LVT div_sub_x_7_U926 ( .A1(div_sub_x_7_n1027), .A2(div_sub_x_7_n1030), 
        .Y(div_sub_x_7_n1028) );
  AO222X1_LVT div_sub_x_7_U925 ( .A1(div_n_T_51_97_), .A2(div_sub_x_7_n853), 
        .A3(div_sub_x_7_n1026), .A4(div_sub_x_7_n1027), .A5(div_sub_x_7_n1028), 
        .A6(div_sub_x_7_n1029), .Y(div_sub_x_7_n1014) );
  AO21X1_LVT div_sub_x_7_U924 ( .A1(div_sub_x_7_n1012), .A2(div_sub_x_7_n834), 
        .A3(div_sub_x_7_n1014), .Y(div_sub_x_7_n1023) );
  FADDX1_LVT div_sub_x_7_U923 ( .A(div_n_T_51_98_), .B(div_sub_x_7_n852), .CI(
        div_sub_x_7_n1023), .S(div_subtractor_35_) );
  NAND2X0_LVT div_sub_x_7_U922 ( .A1(div_n_T_51_98_), .A2(div_sub_x_7_n852), 
        .Y(div_sub_x_7_n1024) );
  OR2X1_LVT div_sub_x_7_U921 ( .A1(div_sub_x_7_n852), .A2(div_n_T_51_98_), .Y(
        div_sub_x_7_n1018) );
  OA21X1_LVT div_sub_x_7_U920 ( .A1(div_sub_x_7_n851), .A2(div_sub_x_7_n1023), 
        .A3(div_sub_x_7_n1018), .Y(div_sub_x_7_n1025) );
  FADDX1_LVT div_sub_x_7_U919 ( .A(div_divisor_36_), .B(div_sub_x_7_n1025), 
        .CI(div_sub_x_7_n893), .S(div_subtractor_36_) );
  AO222X1_LVT div_sub_x_7_U918 ( .A1(div_divisor_36_), .A2(div_sub_x_7_n893), 
        .A3(div_divisor_36_), .A4(div_sub_x_7_n1024), .A5(div_sub_x_7_n893), 
        .A6(div_sub_x_7_n1024), .Y(div_sub_x_7_n1013) );
  NAND2X0_LVT div_sub_x_7_U917 ( .A1(div_divisor_36_), .A2(div_sub_x_7_n893), 
        .Y(div_sub_x_7_n1017) );
  NAND3X0_LVT div_sub_x_7_U916 ( .A1(div_sub_x_7_n1023), .A2(div_sub_x_7_n1017), .A3(div_sub_x_7_n1018), .Y(div_sub_x_7_n1022) );
  AND2X1_LVT div_sub_x_7_U915 ( .A1(div_sub_x_7_n1013), .A2(div_sub_x_7_n1022), 
        .Y(div_sub_x_7_n1021) );
  FADDX1_LVT div_sub_x_7_U914 ( .A(div_n_T_51_100_), .B(div_divisor_37_), .CI(
        div_sub_x_7_n1021), .S(div_subtractor_37_) );
  OR2X1_LVT div_sub_x_7_U913 ( .A1(div_sub_x_7_n892), .A2(div_divisor_37_), 
        .Y(div_sub_x_7_n1019) );
  AO22X1_LVT div_sub_x_7_U912 ( .A1(div_sub_x_7_n1021), .A2(div_sub_x_7_n1019), 
        .A3(div_divisor_37_), .A4(div_sub_x_7_n892), .Y(div_sub_x_7_n1020) );
  FADDX1_LVT div_sub_x_7_U911 ( .A(div_n_T_51_101_), .B(div_divisor_38_), .CI(
        div_sub_x_7_n1020), .S(div_subtractor_38_) );
  NAND2X0_LVT div_sub_x_7_U910 ( .A1(div_divisor_38_), .A2(div_sub_x_7_n891), 
        .Y(div_sub_x_7_n1015) );
  NAND2X0_LVT div_sub_x_7_U909 ( .A1(div_divisor_37_), .A2(div_sub_x_7_n892), 
        .Y(div_sub_x_7_n1016) );
  AND4X1_LVT div_sub_x_7_U908 ( .A1(div_sub_x_7_n1015), .A2(div_sub_x_7_n1016), 
        .A3(div_sub_x_7_n1017), .A4(div_sub_x_7_n1018), .Y(div_sub_x_7_n1011)
         );
  AND2X1_LVT div_sub_x_7_U907 ( .A1(div_sub_x_7_n1011), .A2(div_sub_x_7_n1012), 
        .Y(div_sub_x_7_n988) );
  NAND2X0_LVT div_sub_x_7_U906 ( .A1(div_sub_x_7_n988), .A2(div_sub_x_7_n834), 
        .Y(div_sub_x_7_n1010) );
  NAND2X0_LVT div_sub_x_7_U905 ( .A1(div_sub_x_7_n980), .A2(div_sub_x_7_n1010), 
        .Y(div_sub_x_7_n998) );
  FADDX1_LVT div_sub_x_7_U904 ( .A(div_n_T_51_102_), .B(div_sub_x_7_n850), 
        .CI(div_sub_x_7_n998), .S(div_subtractor_39_) );
  FADDX1_LVT div_sub_x_7_U903 ( .A(div_sub_x_7_n977), .B(div_n_T_51_66_), .CI(
        div_sub_x_7_n874), .S(div_subtractor_3_) );
  AND2X1_LVT div_sub_x_7_U902 ( .A1(div_n_T_51_102_), .A2(div_sub_x_7_n850), 
        .Y(div_sub_x_7_n1008) );
  OR2X1_LVT div_sub_x_7_U901 ( .A1(div_sub_x_7_n850), .A2(div_n_T_51_102_), 
        .Y(div_sub_x_7_n1005) );
  OA21X1_LVT div_sub_x_7_U900 ( .A1(div_sub_x_7_n1008), .A2(div_sub_x_7_n998), 
        .A3(div_sub_x_7_n1005), .Y(div_sub_x_7_n1009) );
  FADDX1_LVT div_sub_x_7_U899 ( .A(div_n_T_51_103_), .B(div_sub_x_7_n1009), 
        .CI(div_sub_x_7_n849), .S(div_subtractor_40_) );
  OR2X1_LVT div_sub_x_7_U898 ( .A1(div_sub_x_7_n849), .A2(div_n_T_51_103_), 
        .Y(div_sub_x_7_n1004) );
  AO22X1_LVT div_sub_x_7_U897 ( .A1(div_n_T_51_103_), .A2(div_sub_x_7_n849), 
        .A3(div_sub_x_7_n1008), .A4(div_sub_x_7_n1004), .Y(div_sub_x_7_n1002)
         );
  OA222X1_LVT div_sub_x_7_U896 ( .A1(div_sub_x_7_n1002), .A2(div_sub_x_7_n1004), .A3(div_sub_x_7_n1002), .A4(div_sub_x_7_n1005), .A5(div_sub_x_7_n1002), .A6(
        div_sub_x_7_n998), .Y(div_sub_x_7_n1007) );
  FADDX1_LVT div_sub_x_7_U895 ( .A(div_n_T_51_104_), .B(div_sub_x_7_n848), 
        .CI(div_sub_x_7_n1007), .S(div_subtractor_41_) );
  AND2X1_LVT div_sub_x_7_U894 ( .A1(div_n_T_51_104_), .A2(div_sub_x_7_n848), 
        .Y(div_sub_x_7_n999) );
  OR2X1_LVT div_sub_x_7_U893 ( .A1(div_sub_x_7_n848), .A2(div_n_T_51_104_), 
        .Y(div_sub_x_7_n1003) );
  OA21X1_LVT div_sub_x_7_U892 ( .A1(div_sub_x_7_n999), .A2(div_sub_x_7_n1007), 
        .A3(div_sub_x_7_n1003), .Y(div_sub_x_7_n1006) );
  FADDX1_LVT div_sub_x_7_U891 ( .A(div_n_T_51_105_), .B(div_sub_x_7_n1006), 
        .CI(div_sub_x_7_n847), .S(div_subtractor_42_) );
  OR2X1_LVT div_sub_x_7_U890 ( .A1(div_sub_x_7_n847), .A2(div_n_T_51_105_), 
        .Y(div_sub_x_7_n1000) );
  AND4X1_LVT div_sub_x_7_U889 ( .A1(div_sub_x_7_n1000), .A2(div_sub_x_7_n1003), 
        .A3(div_sub_x_7_n1004), .A4(div_sub_x_7_n1005), .Y(div_sub_x_7_n989)
         );
  AND2X1_LVT div_sub_x_7_U888 ( .A1(div_sub_x_7_n1000), .A2(div_sub_x_7_n1003), 
        .Y(div_sub_x_7_n1001) );
  AO222X1_LVT div_sub_x_7_U887 ( .A1(div_n_T_51_105_), .A2(div_sub_x_7_n847), 
        .A3(div_sub_x_7_n999), .A4(div_sub_x_7_n1000), .A5(div_sub_x_7_n1001), 
        .A6(div_sub_x_7_n1002), .Y(div_sub_x_7_n984) );
  AO21X1_LVT div_sub_x_7_U886 ( .A1(div_sub_x_7_n989), .A2(div_sub_x_7_n998), 
        .A3(div_sub_x_7_n984), .Y(div_sub_x_7_n995) );
  FADDX1_LVT div_sub_x_7_U885 ( .A(div_n_T_51_106_), .B(div_sub_x_7_n846), 
        .CI(div_sub_x_7_n995), .S(div_subtractor_43_) );
  NAND2X0_LVT div_sub_x_7_U884 ( .A1(div_n_T_51_106_), .A2(div_sub_x_7_n846), 
        .Y(div_sub_x_7_n996) );
  OR2X1_LVT div_sub_x_7_U883 ( .A1(div_sub_x_7_n846), .A2(div_n_T_51_106_), 
        .Y(div_sub_x_7_n991) );
  OA21X1_LVT div_sub_x_7_U882 ( .A1(div_sub_x_7_n845), .A2(div_sub_x_7_n995), 
        .A3(div_sub_x_7_n991), .Y(div_sub_x_7_n997) );
  FADDX1_LVT div_sub_x_7_U881 ( .A(div_divisor_44_), .B(div_sub_x_7_n997), 
        .CI(div_sub_x_7_n890), .S(div_subtractor_44_) );
  AO222X1_LVT div_sub_x_7_U880 ( .A1(div_divisor_44_), .A2(div_sub_x_7_n890), 
        .A3(div_divisor_44_), .A4(div_sub_x_7_n996), .A5(div_sub_x_7_n890), 
        .A6(div_sub_x_7_n996), .Y(div_sub_x_7_n982) );
  NAND2X0_LVT div_sub_x_7_U879 ( .A1(div_divisor_44_), .A2(div_sub_x_7_n890), 
        .Y(div_sub_x_7_n990) );
  NAND3X0_LVT div_sub_x_7_U878 ( .A1(div_sub_x_7_n995), .A2(div_sub_x_7_n990), 
        .A3(div_sub_x_7_n991), .Y(div_sub_x_7_n994) );
  AND2X1_LVT div_sub_x_7_U877 ( .A1(div_sub_x_7_n982), .A2(div_sub_x_7_n994), 
        .Y(div_sub_x_7_n993) );
  FADDX1_LVT div_sub_x_7_U876 ( .A(div_n_T_51_108_), .B(div_divisor_45_), .CI(
        div_sub_x_7_n993), .S(div_subtractor_45_) );
  OR2X1_LVT div_sub_x_7_U875 ( .A1(div_sub_x_7_n889), .A2(div_divisor_45_), 
        .Y(div_sub_x_7_n987) );
  AO22X1_LVT div_sub_x_7_U874 ( .A1(div_sub_x_7_n993), .A2(div_sub_x_7_n987), 
        .A3(div_divisor_45_), .A4(div_sub_x_7_n889), .Y(div_sub_x_7_n992) );
  FADDX1_LVT div_sub_x_7_U873 ( .A(div_n_T_51_109_), .B(div_divisor_46_), .CI(
        div_sub_x_7_n992), .S(div_subtractor_46_) );
  NAND2X0_LVT div_sub_x_7_U872 ( .A1(div_divisor_46_), .A2(div_sub_x_7_n888), 
        .Y(div_sub_x_7_n985) );
  NAND2X0_LVT div_sub_x_7_U871 ( .A1(div_divisor_45_), .A2(div_sub_x_7_n889), 
        .Y(div_sub_x_7_n986) );
  AND4X1_LVT div_sub_x_7_U870 ( .A1(div_sub_x_7_n985), .A2(div_sub_x_7_n986), 
        .A3(div_sub_x_7_n990), .A4(div_sub_x_7_n991), .Y(div_sub_x_7_n983) );
  NAND2X0_LVT div_sub_x_7_U869 ( .A1(div_sub_x_7_n989), .A2(div_sub_x_7_n983), 
        .Y(div_sub_x_7_n981) );
  NAND2X0_LVT div_sub_x_7_U868 ( .A1(div_sub_x_7_n844), .A2(div_sub_x_7_n988), 
        .Y(div_sub_x_7_n919) );
  OA21X1_LVT div_sub_x_7_U867 ( .A1(div_sub_x_7_n918), .A2(div_sub_x_7_n919), 
        .A3(div_sub_x_7_n920), .Y(div_sub_x_7_n950) );
  FADDX1_LVT div_sub_x_7_U866 ( .A(div_n_T_51_110_), .B(div_divisor_47_), .CI(
        div_sub_x_7_n950), .S(div_subtractor_47_) );
  AND2X1_LVT div_sub_x_7_U865 ( .A1(div_n_T_51_110_), .A2(div_sub_x_7_n843), 
        .Y(div_sub_x_7_n978) );
  OR2X1_LVT div_sub_x_7_U864 ( .A1(div_sub_x_7_n843), .A2(div_n_T_51_110_), 
        .Y(div_sub_x_7_n972) );
  OA21X1_LVT div_sub_x_7_U863 ( .A1(div_sub_x_7_n978), .A2(div_sub_x_7_n835), 
        .A3(div_sub_x_7_n972), .Y(div_sub_x_7_n979) );
  FADDX1_LVT div_sub_x_7_U862 ( .A(div_n_T_51_111_), .B(div_sub_x_7_n979), 
        .CI(div_sub_x_7_n842), .S(div_subtractor_48_) );
  OR2X1_LVT div_sub_x_7_U861 ( .A1(div_sub_x_7_n842), .A2(div_n_T_51_111_), 
        .Y(div_sub_x_7_n971) );
  AO22X1_LVT div_sub_x_7_U860 ( .A1(div_n_T_51_111_), .A2(div_sub_x_7_n842), 
        .A3(div_sub_x_7_n978), .A4(div_sub_x_7_n971), .Y(div_sub_x_7_n969) );
  OA222X1_LVT div_sub_x_7_U859 ( .A1(div_sub_x_7_n969), .A2(div_sub_x_7_n971), 
        .A3(div_sub_x_7_n969), .A4(div_sub_x_7_n972), .A5(div_sub_x_7_n969), 
        .A6(div_sub_x_7_n835), .Y(div_sub_x_7_n974) );
  FADDX1_LVT div_sub_x_7_U858 ( .A(div_n_T_51_112_), .B(div_sub_x_7_n841), 
        .CI(div_sub_x_7_n974), .S(div_subtractor_49_) );
  AO22X1_LVT div_sub_x_7_U857 ( .A1(div_divisor_3_), .A2(div_sub_x_7_n905), 
        .A3(div_sub_x_7_n875), .A4(div_sub_x_7_n976), .Y(div_sub_x_7_n975) );
  FADDX1_LVT div_sub_x_7_U856 ( .A(div_n_T_51_67_), .B(div_divisor_4_), .CI(
        div_sub_x_7_n975), .S(div_subtractor_4_) );
  AND2X1_LVT div_sub_x_7_U855 ( .A1(div_n_T_51_112_), .A2(div_sub_x_7_n841), 
        .Y(div_sub_x_7_n966) );
  OR2X1_LVT div_sub_x_7_U854 ( .A1(div_sub_x_7_n841), .A2(div_n_T_51_112_), 
        .Y(div_sub_x_7_n970) );
  OA21X1_LVT div_sub_x_7_U853 ( .A1(div_sub_x_7_n966), .A2(div_sub_x_7_n974), 
        .A3(div_sub_x_7_n970), .Y(div_sub_x_7_n973) );
  FADDX1_LVT div_sub_x_7_U852 ( .A(div_n_T_51_113_), .B(div_sub_x_7_n973), 
        .CI(div_sub_x_7_n840), .S(div_subtractor_50_) );
  OR2X1_LVT div_sub_x_7_U851 ( .A1(div_sub_x_7_n840), .A2(div_n_T_51_113_), 
        .Y(div_sub_x_7_n967) );
  AND4X1_LVT div_sub_x_7_U850 ( .A1(div_sub_x_7_n967), .A2(div_sub_x_7_n970), 
        .A3(div_sub_x_7_n971), .A4(div_sub_x_7_n972), .Y(div_sub_x_7_n957) );
  AND2X1_LVT div_sub_x_7_U849 ( .A1(div_sub_x_7_n967), .A2(div_sub_x_7_n970), 
        .Y(div_sub_x_7_n968) );
  AO222X1_LVT div_sub_x_7_U848 ( .A1(div_n_T_51_113_), .A2(div_sub_x_7_n840), 
        .A3(div_sub_x_7_n966), .A4(div_sub_x_7_n967), .A5(div_sub_x_7_n968), 
        .A6(div_sub_x_7_n969), .Y(div_sub_x_7_n953) );
  AO21X1_LVT div_sub_x_7_U847 ( .A1(div_sub_x_7_n957), .A2(div_sub_x_7_n835), 
        .A3(div_sub_x_7_n953), .Y(div_sub_x_7_n963) );
  FADDX1_LVT div_sub_x_7_U846 ( .A(div_n_T_51_114_), .B(div_sub_x_7_n839), 
        .CI(div_sub_x_7_n963), .S(div_subtractor_51_) );
  NAND2X0_LVT div_sub_x_7_U845 ( .A1(div_n_T_51_114_), .A2(div_sub_x_7_n839), 
        .Y(div_sub_x_7_n964) );
  OR2X1_LVT div_sub_x_7_U844 ( .A1(div_sub_x_7_n839), .A2(div_n_T_51_114_), 
        .Y(div_sub_x_7_n959) );
  OA21X1_LVT div_sub_x_7_U843 ( .A1(div_sub_x_7_n838), .A2(div_sub_x_7_n963), 
        .A3(div_sub_x_7_n959), .Y(div_sub_x_7_n965) );
  FADDX1_LVT div_sub_x_7_U842 ( .A(div_divisor_52_), .B(div_sub_x_7_n965), 
        .CI(div_sub_x_7_n887), .S(div_subtractor_52_) );
  AO222X1_LVT div_sub_x_7_U841 ( .A1(div_divisor_52_), .A2(div_sub_x_7_n887), 
        .A3(div_divisor_52_), .A4(div_sub_x_7_n964), .A5(div_sub_x_7_n887), 
        .A6(div_sub_x_7_n964), .Y(div_sub_x_7_n951) );
  NAND2X0_LVT div_sub_x_7_U840 ( .A1(div_divisor_52_), .A2(div_sub_x_7_n887), 
        .Y(div_sub_x_7_n958) );
  NAND3X0_LVT div_sub_x_7_U839 ( .A1(div_sub_x_7_n963), .A2(div_sub_x_7_n958), 
        .A3(div_sub_x_7_n959), .Y(div_sub_x_7_n962) );
  AND2X1_LVT div_sub_x_7_U838 ( .A1(div_sub_x_7_n951), .A2(div_sub_x_7_n962), 
        .Y(div_sub_x_7_n961) );
  FADDX1_LVT div_sub_x_7_U837 ( .A(div_n_T_51_116_), .B(div_divisor_53_), .CI(
        div_sub_x_7_n961), .S(div_subtractor_53_) );
  OR2X1_LVT div_sub_x_7_U836 ( .A1(div_sub_x_7_n886), .A2(div_divisor_53_), 
        .Y(div_sub_x_7_n956) );
  AO22X1_LVT div_sub_x_7_U835 ( .A1(div_sub_x_7_n961), .A2(div_sub_x_7_n956), 
        .A3(div_divisor_53_), .A4(div_sub_x_7_n886), .Y(div_sub_x_7_n960) );
  FADDX1_LVT div_sub_x_7_U834 ( .A(div_n_T_51_117_), .B(div_divisor_54_), .CI(
        div_sub_x_7_n960), .S(div_subtractor_54_) );
  NAND2X0_LVT div_sub_x_7_U833 ( .A1(div_divisor_54_), .A2(div_sub_x_7_n885), 
        .Y(div_sub_x_7_n954) );
  NAND2X0_LVT div_sub_x_7_U832 ( .A1(div_divisor_53_), .A2(div_sub_x_7_n886), 
        .Y(div_sub_x_7_n955) );
  AND4X1_LVT div_sub_x_7_U831 ( .A1(div_sub_x_7_n954), .A2(div_sub_x_7_n955), 
        .A3(div_sub_x_7_n958), .A4(div_sub_x_7_n959), .Y(div_sub_x_7_n952) );
  NAND2X0_LVT div_sub_x_7_U830 ( .A1(div_sub_x_7_n952), .A2(div_sub_x_7_n957), 
        .Y(div_sub_x_7_n924) );
  OA21X1_LVT div_sub_x_7_U829 ( .A1(div_sub_x_7_n950), .A2(div_sub_x_7_n924), 
        .A3(div_sub_x_7_n921), .Y(div_sub_x_7_n936) );
  FADDX1_LVT div_sub_x_7_U828 ( .A(div_n_T_51_118_), .B(div_divisor_55_), .CI(
        div_sub_x_7_n936), .S(div_subtractor_55_) );
  OR2X1_LVT div_sub_x_7_U827 ( .A1(div_sub_x_7_n884), .A2(div_divisor_55_), 
        .Y(div_sub_x_7_n948) );
  AO22X1_LVT div_sub_x_7_U826 ( .A1(div_sub_x_7_n936), .A2(div_sub_x_7_n948), 
        .A3(div_divisor_55_), .A4(div_sub_x_7_n884), .Y(div_sub_x_7_n949) );
  FADDX1_LVT div_sub_x_7_U825 ( .A(div_n_T_51_119_), .B(div_divisor_56_), .CI(
        div_sub_x_7_n949), .S(div_subtractor_56_) );
  NAND2X0_LVT div_sub_x_7_U824 ( .A1(div_divisor_56_), .A2(div_sub_x_7_n883), 
        .Y(div_sub_x_7_n943) );
  NAND2X0_LVT div_sub_x_7_U823 ( .A1(div_divisor_55_), .A2(div_sub_x_7_n884), 
        .Y(div_sub_x_7_n944) );
  NAND2X0_LVT div_sub_x_7_U822 ( .A1(div_sub_x_7_n943), .A2(div_sub_x_7_n944), 
        .Y(div_sub_x_7_n947) );
  AO222X1_LVT div_sub_x_7_U821 ( .A1(div_divisor_56_), .A2(div_sub_x_7_n883), 
        .A3(div_divisor_56_), .A4(div_sub_x_7_n948), .A5(div_sub_x_7_n883), 
        .A6(div_sub_x_7_n948), .Y(div_sub_x_7_n937) );
  OA21X1_LVT div_sub_x_7_U820 ( .A1(div_sub_x_7_n936), .A2(div_sub_x_7_n947), 
        .A3(div_sub_x_7_n937), .Y(div_sub_x_7_n946) );
  FADDX1_LVT div_sub_x_7_U819 ( .A(div_n_T_51_120_), .B(div_divisor_57_), .CI(
        div_sub_x_7_n946), .S(div_subtractor_57_) );
  OR2X1_LVT div_sub_x_7_U818 ( .A1(div_sub_x_7_n882), .A2(div_divisor_57_), 
        .Y(div_sub_x_7_n940) );
  AO22X1_LVT div_sub_x_7_U817 ( .A1(div_sub_x_7_n946), .A2(div_sub_x_7_n940), 
        .A3(div_divisor_57_), .A4(div_sub_x_7_n882), .Y(div_sub_x_7_n945) );
  FADDX1_LVT div_sub_x_7_U816 ( .A(div_n_T_51_121_), .B(div_divisor_58_), .CI(
        div_sub_x_7_n945), .S(div_subtractor_58_) );
  NAND2X0_LVT div_sub_x_7_U815 ( .A1(div_divisor_58_), .A2(div_sub_x_7_n881), 
        .Y(div_sub_x_7_n941) );
  NAND2X0_LVT div_sub_x_7_U814 ( .A1(div_divisor_57_), .A2(div_sub_x_7_n882), 
        .Y(div_sub_x_7_n942) );
  NAND4X0_LVT div_sub_x_7_U813 ( .A1(div_sub_x_7_n941), .A2(div_sub_x_7_n942), 
        .A3(div_sub_x_7_n943), .A4(div_sub_x_7_n944), .Y(div_sub_x_7_n925) );
  NAND2X0_LVT div_sub_x_7_U812 ( .A1(div_sub_x_7_n941), .A2(div_sub_x_7_n942), 
        .Y(div_sub_x_7_n938) );
  AO222X1_LVT div_sub_x_7_U811 ( .A1(div_divisor_58_), .A2(div_sub_x_7_n881), 
        .A3(div_divisor_58_), .A4(div_sub_x_7_n940), .A5(div_sub_x_7_n881), 
        .A6(div_sub_x_7_n940), .Y(div_sub_x_7_n939) );
  OA21X1_LVT div_sub_x_7_U810 ( .A1(div_sub_x_7_n937), .A2(div_sub_x_7_n938), 
        .A3(div_sub_x_7_n939), .Y(div_sub_x_7_n922) );
  OA21X1_LVT div_sub_x_7_U809 ( .A1(div_sub_x_7_n936), .A2(div_sub_x_7_n925), 
        .A3(div_sub_x_7_n922), .Y(div_sub_x_7_n930) );
  FADDX1_LVT div_sub_x_7_U808 ( .A(div_n_T_51_122_), .B(div_divisor_59_), .CI(
        div_sub_x_7_n930), .S(div_subtractor_59_) );
  NAND2X0_LVT div_sub_x_7_U807 ( .A1(div_sub_x_7_n934), .A2(div_sub_x_7_n935), 
        .Y(div_sub_x_7_n914) );
  FADDX1_LVT div_sub_x_7_U806 ( .A(div_n_T_51_68_), .B(div_sub_x_7_n914), .CI(
        div_sub_x_7_n873), .S(div_subtractor_5_) );
  OR2X1_LVT div_sub_x_7_U805 ( .A1(div_sub_x_7_n837), .A2(div_n_T_51_122_), 
        .Y(div_sub_x_7_n927) );
  NAND2X0_LVT div_sub_x_7_U804 ( .A1(div_n_T_51_122_), .A2(div_sub_x_7_n837), 
        .Y(div_sub_x_7_n932) );
  OA21X1_LVT div_sub_x_7_U803 ( .A1(div_sub_x_7_n836), .A2(div_sub_x_7_n930), 
        .A3(div_sub_x_7_n932), .Y(div_sub_x_7_n933) );
  FADDX1_LVT div_sub_x_7_U802 ( .A(div_n_T_51_123_), .B(div_divisor_60_), .CI(
        div_sub_x_7_n933), .S(div_subtractor_60_) );
  NAND2X0_LVT div_sub_x_7_U801 ( .A1(div_divisor_60_), .A2(div_sub_x_7_n880), 
        .Y(div_sub_x_7_n926) );
  NAND2X0_LVT div_sub_x_7_U800 ( .A1(div_sub_x_7_n926), .A2(div_sub_x_7_n927), 
        .Y(div_sub_x_7_n931) );
  AO222X1_LVT div_sub_x_7_U799 ( .A1(div_divisor_60_), .A2(div_sub_x_7_n880), 
        .A3(div_divisor_60_), .A4(div_sub_x_7_n932), .A5(div_sub_x_7_n880), 
        .A6(div_sub_x_7_n932), .Y(div_sub_x_7_n923) );
  OA21X1_LVT div_sub_x_7_U798 ( .A1(div_sub_x_7_n930), .A2(div_sub_x_7_n931), 
        .A3(div_sub_x_7_n923), .Y(div_sub_x_7_n929) );
  FADDX1_LVT div_sub_x_7_U797 ( .A(div_n_T_51_124_), .B(div_divisor_61_), .CI(
        div_sub_x_7_n929), .S(div_subtractor_61_) );
  AO222X1_LVT div_sub_x_7_U796 ( .A1(div_divisor_61_), .A2(div_sub_x_7_n879), 
        .A3(div_divisor_61_), .A4(div_sub_x_7_n929), .A5(div_sub_x_7_n879), 
        .A6(div_sub_x_7_n929), .Y(div_sub_x_7_n928) );
  FADDX1_LVT div_sub_x_7_U795 ( .A(div_sub_x_7_n928), .B(div_n_T_51_125_), 
        .CI(div_divisor_62_), .S(div_subtractor_62_) );
  FADDX1_LVT div_sub_x_7_U794 ( .A(div_n_T_51_126_), .B(div_divisor_63_), .CI(
        div_sub_x_7_n917), .S(div_subtractor_63_) );
  AO222X1_LVT div_sub_x_7_U793 ( .A1(div_divisor_63_), .A2(div_sub_x_7_n878), 
        .A3(div_divisor_63_), .A4(div_sub_x_7_n917), .A5(div_sub_x_7_n878), 
        .A6(div_sub_x_7_n917), .Y(div_sub_x_7_n916) );
  FADDX1_LVT div_sub_x_7_U792 ( .A(div_divisor_64_), .B(div_n_T_51_127_), .CI(
        div_sub_x_7_n916), .S(div_subtractor_64_) );
  AO22X1_LVT div_sub_x_7_U791 ( .A1(div_n_T_51_68_), .A2(div_sub_x_7_n873), 
        .A3(div_sub_x_7_n914), .A4(div_sub_x_7_n915), .Y(div_sub_x_7_n913) );
  FADDX1_LVT div_sub_x_7_U790 ( .A(div_divisor_6_), .B(div_sub_x_7_n903), .CI(
        div_sub_x_7_n913), .S(div_subtractor_6_) );
  FADDX1_LVT div_sub_x_7_U789 ( .A(div_n_T_51_70_), .B(div_divisor_7_), .CI(
        div_sub_x_7_n912), .S(div_subtractor_7_) );
  AO21X1_LVT div_sub_x_7_U788 ( .A1(div_sub_x_7_n910), .A2(div_sub_x_7_n872), 
        .A3(div_sub_x_7_n911), .Y(div_sub_x_7_n909) );
  FADDX1_LVT div_sub_x_7_U787 ( .A(div_n_T_51_71_), .B(div_sub_x_7_n871), .CI(
        div_sub_x_7_n909), .S(div_subtractor_8_) );
  FADDX1_LVT div_sub_x_7_U786 ( .A(div_divisor_9_), .B(div_sub_x_7_n901), .CI(
        div_sub_x_7_n908), .S(div_subtractor_9_) );
  INVX1_LVT div_sub_x_7_U785 ( .A(div_divisor_3_), .Y(div_sub_x_7_n874) );
  INVX1_LVT div_sub_x_7_U784 ( .A(div_divisor_16_), .Y(div_sub_x_7_n866) );
  INVX1_LVT div_sub_x_7_U783 ( .A(div_divisor_17_), .Y(div_sub_x_7_n865) );
  INVX1_LVT div_sub_x_7_U782 ( .A(div_divisor_18_), .Y(div_sub_x_7_n864) );
  INVX1_LVT div_sub_x_7_U781 ( .A(div_divisor_19_), .Y(div_sub_x_7_n863) );
  INVX1_LVT div_sub_x_7_U780 ( .A(div_divisor_23_), .Y(div_sub_x_7_n861) );
  INVX1_LVT div_sub_x_7_U779 ( .A(div_divisor_25_), .Y(div_sub_x_7_n859) );
  INVX1_LVT div_sub_x_7_U778 ( .A(div_divisor_32_), .Y(div_sub_x_7_n855) );
  INVX1_LVT div_sub_x_7_U777 ( .A(div_divisor_33_), .Y(div_sub_x_7_n854) );
  INVX1_LVT div_sub_x_7_U776 ( .A(div_divisor_34_), .Y(div_sub_x_7_n853) );
  INVX1_LVT div_sub_x_7_U775 ( .A(div_divisor_35_), .Y(div_sub_x_7_n852) );
  INVX1_LVT div_sub_x_7_U774 ( .A(div_divisor_39_), .Y(div_sub_x_7_n850) );
  INVX1_LVT div_sub_x_7_U773 ( .A(div_divisor_40_), .Y(div_sub_x_7_n849) );
  INVX1_LVT div_sub_x_7_U772 ( .A(div_divisor_41_), .Y(div_sub_x_7_n848) );
  INVX1_LVT div_sub_x_7_U771 ( .A(div_divisor_42_), .Y(div_sub_x_7_n847) );
  INVX1_LVT div_sub_x_7_U770 ( .A(div_divisor_43_), .Y(div_sub_x_7_n846) );
  INVX1_LVT div_sub_x_7_U769 ( .A(div_divisor_48_), .Y(div_sub_x_7_n842) );
  INVX1_LVT div_sub_x_7_U768 ( .A(div_divisor_49_), .Y(div_sub_x_7_n841) );
  INVX1_LVT div_sub_x_7_U767 ( .A(div_divisor_50_), .Y(div_sub_x_7_n840) );
  INVX1_LVT div_sub_x_7_U766 ( .A(div_divisor_51_), .Y(div_sub_x_7_n839) );
  INVX1_LVT div_sub_x_7_U765 ( .A(div_sub_x_7_n927), .Y(div_sub_x_7_n836) );
  INVX1_LVT div_sub_x_7_U764 ( .A(div_n301), .Y(div_sub_x_7_n833) );
  INVX1_LVT div_sub_x_7_U763 ( .A(div_divisor_26_), .Y(div_sub_x_7_n858) );
  INVX1_LVT div_sub_x_7_U762 ( .A(div_divisor_24_), .Y(div_sub_x_7_n860) );
  INVX1_LVT div_sub_x_7_U761 ( .A(div_divisor_29_), .Y(div_sub_x_7_n856) );
  INVX1_LVT div_sub_x_7_U760 ( .A(div_divisor_27_), .Y(div_sub_x_7_n857) );
  INVX1_LVT div_sub_x_7_U759 ( .A(div_divisor_21_), .Y(div_sub_x_7_n862) );
  INVX1_LVT div_sub_x_7_U758 ( .A(div_divisor_15_), .Y(div_sub_x_7_n867) );
  INVX1_LVT div_sub_x_7_U757 ( .A(div_divisor_11_), .Y(div_sub_x_7_n869) );
  INVX1_LVT div_sub_x_7_U756 ( .A(div_divisor_10_), .Y(div_sub_x_7_n870) );
  INVX1_LVT div_sub_x_7_U755 ( .A(div_divisor_8_), .Y(div_sub_x_7_n871) );
  INVX1_LVT div_sub_x_7_U754 ( .A(div_divisor_5_), .Y(div_sub_x_7_n873) );
  INVX0_LVT div_sub_x_7_U753 ( .A(div_n_T_51_108_), .Y(div_sub_x_7_n889) );
  INVX0_LVT div_sub_x_7_U752 ( .A(div_n_T_51_109_), .Y(div_sub_x_7_n888) );
  INVX0_LVT div_sub_x_7_U751 ( .A(div_n_T_51_107_), .Y(div_sub_x_7_n890) );
  INVX0_LVT div_sub_x_7_U750 ( .A(div_n_T_51_100_), .Y(div_sub_x_7_n892) );
  INVX0_LVT div_sub_x_7_U749 ( .A(div_n_T_51_101_), .Y(div_sub_x_7_n891) );
  INVX0_LVT div_sub_x_7_U748 ( .A(div_n_T_51_99_), .Y(div_sub_x_7_n893) );
  INVX0_LVT div_sub_x_7_U747 ( .A(div_divisor_59_), .Y(div_sub_x_7_n837) );
  INVX0_LVT div_sub_x_7_U746 ( .A(div_n_T_51_123_), .Y(div_sub_x_7_n880) );
  INVX0_LVT div_sub_x_7_U745 ( .A(div_n_T_51_124_), .Y(div_sub_x_7_n879) );
  INVX0_LVT div_sub_x_7_U744 ( .A(div_n_T_51_118_), .Y(div_sub_x_7_n884) );
  INVX0_LVT div_sub_x_7_U743 ( .A(div_n_T_51_119_), .Y(div_sub_x_7_n883) );
  INVX0_LVT div_sub_x_7_U742 ( .A(div_n_T_51_120_), .Y(div_sub_x_7_n882) );
  INVX0_LVT div_sub_x_7_U741 ( .A(div_n_T_51_121_), .Y(div_sub_x_7_n881) );
  INVX0_LVT div_sub_x_7_U740 ( .A(div_divisor_47_), .Y(div_sub_x_7_n843) );
  INVX0_LVT div_sub_x_7_U739 ( .A(div_n_T_51_115_), .Y(div_sub_x_7_n887) );
  INVX0_LVT div_sub_x_7_U738 ( .A(div_n_T_51_116_), .Y(div_sub_x_7_n886) );
  INVX0_LVT div_sub_x_7_U737 ( .A(div_n_T_51_117_), .Y(div_sub_x_7_n885) );
  INVX0_LVT div_sub_x_7_U736 ( .A(div_n_T_51_85_), .Y(div_sub_x_7_n897) );
  INVX0_LVT div_sub_x_7_U735 ( .A(div_n_T_51_126_), .Y(div_sub_x_7_n878) );
  INVX0_LVT div_sub_x_7_U734 ( .A(div_n_T_51_72_), .Y(div_sub_x_7_n901) );
  INVX0_LVT div_sub_x_7_U733 ( .A(div_n_T_51_70_), .Y(div_sub_x_7_n902) );
  INVX0_LVT div_sub_x_7_U732 ( .A(div_n_T_51_69_), .Y(div_sub_x_7_n903) );
  INVX0_LVT div_sub_x_7_U731 ( .A(div_n_T_51_66_), .Y(div_sub_x_7_n905) );
  INVX0_LVT div_sub_x_7_U730 ( .A(div_n_T_51_64_), .Y(div_sub_x_7_n907) );
  INVX0_LVT div_sub_x_7_U729 ( .A(div_n_T_51_65_), .Y(div_sub_x_7_n906) );
  INVX0_LVT div_sub_x_7_U728 ( .A(div_divisor_1_), .Y(div_sub_x_7_n876) );
  INVX0_LVT div_sub_x_7_U727 ( .A(div_n_T_51_67_), .Y(div_sub_x_7_n904) );
  INVX0_LVT div_sub_x_7_U726 ( .A(div_divisor_0_), .Y(div_sub_x_7_n877) );
  INVX0_LVT div_sub_x_7_U725 ( .A(div_n_T_51_75_), .Y(div_sub_x_7_n900) );
  INVX0_LVT div_sub_x_7_U724 ( .A(div_n_T_51_76_), .Y(div_sub_x_7_n899) );
  INVX0_LVT div_sub_x_7_U723 ( .A(div_n_T_51_94_), .Y(div_sub_x_7_n894) );
  INVX0_LVT div_sub_x_7_U722 ( .A(div_n_T_51_93_), .Y(div_sub_x_7_n895) );
  INVX0_LVT div_sub_x_7_U721 ( .A(div_n_T_51_91_), .Y(div_sub_x_7_n896) );
  INVX0_LVT div_sub_x_7_U720 ( .A(div_n_T_51_83_), .Y(div_sub_x_7_n898) );
  NOR2X1_LVT div_sub_x_7_U719 ( .A1(div_sub_x_7_n902), .A2(div_divisor_7_), 
        .Y(div_sub_x_7_n911) );
  NOR2X1_LVT div_sub_x_7_U718 ( .A1(div_sub_x_7_n894), .A2(div_divisor_31_), 
        .Y(div_sub_x_7_n1035) );
  INVX0_LVT div_sub_x_7_U717 ( .A(div_sub_x_7_n1024), .Y(div_sub_x_7_n851) );
  INVX0_LVT div_sub_x_7_U716 ( .A(div_sub_x_7_n1102), .Y(div_sub_x_7_n868) );
  INVX0_LVT div_sub_x_7_U715 ( .A(div_sub_x_7_n996), .Y(div_sub_x_7_n845) );
  INVX0_LVT div_sub_x_7_U714 ( .A(div_sub_x_7_n964), .Y(div_sub_x_7_n838) );
  INVX0_LVT div_sub_x_7_U713 ( .A(div_sub_x_7_n981), .Y(div_sub_x_7_n844) );
  INVX0_LVT div_sub_x_7_U712 ( .A(div_sub_x_7_n977), .Y(div_sub_x_7_n875) );
  INVX0_LVT div_sub_x_7_U711 ( .A(div_sub_x_7_n912), .Y(div_sub_x_7_n872) );
  INVX0_LVT div_sub_x_7_U710 ( .A(div_sub_x_7_n918), .Y(div_sub_x_7_n834) );
  INVX0_LVT div_sub_x_7_U709 ( .A(div_sub_x_7_n950), .Y(div_sub_x_7_n835) );
  NAND2X0_LVT div_sub_x_7_U708 ( .A1(div_sub_x_7_n1037), .A2(div_sub_x_7_n832), 
        .Y(div_sub_x_7_n1055) );
  NAND2X0_LVT div_sub_x_7_U707 ( .A1(div_sub_x_7_n1041), .A2(div_sub_x_7_n1042), .Y(div_sub_x_7_n832) );
  AND4X1_LVT div_sub_x_7_U706 ( .A1(div_sub_x_7_n827), .A2(div_sub_x_7_n829), 
        .A3(div_sub_x_7_n830), .A4(div_sub_x_7_n831), .Y(div_sub_x_7_n920) );
  AO222X1_LVT div_sub_x_7_U705 ( .A1(div_divisor_46_), .A2(div_sub_x_7_n888), 
        .A3(div_divisor_46_), .A4(div_sub_x_7_n987), .A5(div_sub_x_7_n888), 
        .A6(div_sub_x_7_n987), .Y(div_sub_x_7_n831) );
  NAND2X0_LVT div_sub_x_7_U704 ( .A1(div_sub_x_7_n983), .A2(div_sub_x_7_n984), 
        .Y(div_sub_x_7_n830) );
  NAND3X0_LVT div_sub_x_7_U703 ( .A1(div_sub_x_7_n986), .A2(div_sub_x_7_n985), 
        .A3(div_sub_x_7_n828), .Y(div_sub_x_7_n829) );
  INVX0_LVT div_sub_x_7_U702 ( .A(div_sub_x_7_n982), .Y(div_sub_x_7_n828) );
  OR2X1_LVT div_sub_x_7_U701 ( .A1(div_sub_x_7_n981), .A2(div_sub_x_7_n980), 
        .Y(div_sub_x_7_n827) );
  NAND2X0_LVT div_sub_x_7_U699 ( .A1(div_sub_x_7_n1069), .A2(div_sub_x_7_n1068), .Y(div_sub_x_7_n825) );
  NAND2X0_LVT div_sub_x_7_U698 ( .A1(div_sub_x_7_n1070), .A2(div_sub_x_7_n1071), .Y(div_sub_x_7_n824) );
  AO222X1_LVT div_sub_x_7_U697 ( .A1(div_divisor_22_), .A2(div_sub_x_7_n897), 
        .A3(div_divisor_22_), .A4(div_sub_x_7_n822), .A5(div_sub_x_7_n897), 
        .A6(div_sub_x_7_n822), .Y(div_sub_x_7_n823) );
  NAND2X0_LVT div_sub_x_7_U696 ( .A1(div_sub_x_7_n862), .A2(div_n_T_51_84_), 
        .Y(div_sub_x_7_n822) );
  OAI222X1_LVT div_sub_x_7_U694 ( .A1(div_sub_x_7_n816), .A2(div_divisor_14_), 
        .A3(div_sub_x_7_n816), .A4(div_sub_x_7_n1097), .A5(div_divisor_14_), 
        .A6(div_sub_x_7_n1097), .Y(div_sub_x_7_n820) );
  AND3X1_LVT div_sub_x_7_U693 ( .A1(div_sub_x_7_n1096), .A2(div_sub_x_7_n817), 
        .A3(div_sub_x_7_n1095), .Y(div_sub_x_7_n819) );
  AO21X1_LVT div_sub_x_7_U692 ( .A1(div_sub_x_7_n872), .A2(div_sub_x_7_n1092), 
        .A3(div_sub_x_7_n1094), .Y(div_sub_x_7_n818) );
  AOI22X1_LVT div_sub_x_7_U691 ( .A1(div_sub_x_7_n899), .A2(div_divisor_13_), 
        .A3(div_divisor_14_), .A4(div_sub_x_7_n816), .Y(div_sub_x_7_n817) );
  INVX0_LVT div_sub_x_7_U690 ( .A(div_n_T_51_77_), .Y(div_sub_x_7_n816) );
  INVX0_LVT div_sub_x_7_U689 ( .A(div_sub_x_7_n1093), .Y(div_sub_x_7_n815) );
  NAND2X0_LVT div_sub_x_7_U687 ( .A1(div_sub_x_7_n1014), .A2(div_sub_x_7_n1011), .Y(div_sub_x_7_n813) );
  NAND2X0_LVT div_sub_x_7_U686 ( .A1(div_sub_x_7_n1015), .A2(div_sub_x_7_n1016), .Y(div_sub_x_7_n812) );
  AO222X1_LVT div_sub_x_7_U685 ( .A1(div_divisor_38_), .A2(div_sub_x_7_n891), 
        .A3(div_divisor_38_), .A4(div_sub_x_7_n1019), .A5(div_sub_x_7_n891), 
        .A6(div_sub_x_7_n1019), .Y(div_sub_x_7_n811) );
  OA221X1_LVT div_sub_x_7_U684 ( .A1(div_sub_x_7_n803), .A2(div_sub_x_7_n1037), 
        .A3(div_sub_x_7_n803), .A4(div_sub_x_7_n804), .A5(div_sub_x_7_n810), 
        .Y(div_sub_x_7_n918) );
  AO222X1_LVT div_sub_x_7_U682 ( .A1(div_divisor_30_), .A2(div_sub_x_7_n895), 
        .A3(div_divisor_30_), .A4(div_sub_x_7_n807), .A5(div_sub_x_7_n895), 
        .A6(div_sub_x_7_n807), .Y(div_sub_x_7_n808) );
  NAND2X0_LVT div_sub_x_7_U681 ( .A1(div_sub_x_7_n856), .A2(div_n_T_51_92_), 
        .Y(div_sub_x_7_n807) );
  NAND2X0_LVT div_sub_x_7_U680 ( .A1(div_sub_x_7_n1040), .A2(div_sub_x_7_n801), 
        .Y(div_sub_x_7_n806) );
  NAND2X0_LVT div_sub_x_7_U679 ( .A1(div_sub_x_7_n802), .A2(div_sub_x_7_n1039), 
        .Y(div_sub_x_7_n805) );
  NAND2X0_LVT div_sub_x_7_U678 ( .A1(div_sub_x_7_n1041), .A2(div_sub_x_7_n1042), .Y(div_sub_x_7_n804) );
  NAND2X0_LVT div_sub_x_7_U677 ( .A1(div_sub_x_7_n802), .A2(div_sub_x_7_n1043), 
        .Y(div_sub_x_7_n803) );
  AND4X1_LVT div_sub_x_7_U676 ( .A1(div_sub_x_7_n1045), .A2(div_sub_x_7_n1044), 
        .A3(div_sub_x_7_n1040), .A4(div_sub_x_7_n801), .Y(div_sub_x_7_n802) );
  NAND2X0_LVT div_sub_x_7_U675 ( .A1(div_divisor_30_), .A2(div_sub_x_7_n895), 
        .Y(div_sub_x_7_n801) );
  OR3X1_LVT div_sub_x_7_U674 ( .A1(div_sub_x_7_n918), .A2(div_sub_x_7_n919), 
        .A3(div_sub_x_7_n799), .Y(div_sub_x_7_n800) );
  OR2X1_LVT div_sub_x_7_U673 ( .A1(div_sub_x_7_n924), .A2(div_sub_x_7_n794), 
        .Y(div_sub_x_7_n799) );
  AO222X1_LVT div_sub_x_7_U671 ( .A1(div_divisor_62_), .A2(div_sub_x_7_n789), 
        .A3(div_divisor_62_), .A4(div_sub_x_7_n795), .A5(div_sub_x_7_n789), 
        .A6(div_sub_x_7_n795), .Y(div_sub_x_7_n796) );
  OR2X1_LVT div_sub_x_7_U670 ( .A1(div_divisor_61_), .A2(div_sub_x_7_n879), 
        .Y(div_sub_x_7_n795) );
  OR2X1_LVT div_sub_x_7_U669 ( .A1(div_sub_x_7_n925), .A2(div_sub_x_7_n792), 
        .Y(div_sub_x_7_n794) );
  OA22X1_LVT div_sub_x_7_U668 ( .A1(div_sub_x_7_n923), .A2(div_sub_x_7_n790), 
        .A3(div_sub_x_7_n922), .A4(div_sub_x_7_n792), .Y(div_sub_x_7_n793) );
  NAND3X0_LVT div_sub_x_7_U667 ( .A1(div_sub_x_7_n927), .A2(div_sub_x_7_n926), 
        .A3(div_sub_x_7_n791), .Y(div_sub_x_7_n792) );
  INVX0_LVT div_sub_x_7_U666 ( .A(div_sub_x_7_n790), .Y(div_sub_x_7_n791) );
  AO22X1_LVT div_sub_x_7_U665 ( .A1(div_divisor_61_), .A2(div_sub_x_7_n879), 
        .A3(div_divisor_62_), .A4(div_sub_x_7_n789), .Y(div_sub_x_7_n790) );
  INVX0_LVT div_sub_x_7_U664 ( .A(div_n_T_51_125_), .Y(div_sub_x_7_n789) );
  NAND2X0_LVT div_sub_x_7_U663 ( .A1(div_sub_x_7_n953), .A2(div_sub_x_7_n952), 
        .Y(div_sub_x_7_n788) );
  NAND2X0_LVT div_sub_x_7_U662 ( .A1(div_sub_x_7_n954), .A2(div_sub_x_7_n955), 
        .Y(div_sub_x_7_n787) );
  AO222X1_LVT div_sub_x_7_U661 ( .A1(div_divisor_54_), .A2(div_sub_x_7_n885), 
        .A3(div_divisor_54_), .A4(div_sub_x_7_n956), .A5(div_sub_x_7_n885), 
        .A6(div_sub_x_7_n956), .Y(div_sub_x_7_n786) );
  OA21X1_LVT div_sub_x_7_U659 ( .A1(div_sub_x_7_n782), .A2(div_sub_x_7_n783), 
        .A3(div_sub_x_7_n784), .Y(div_sub_x_7_n977) );
  AO222X1_LVT div_sub_x_7_U658 ( .A1(div_sub_x_7_n783), .A2(div_sub_x_7_n782), 
        .A3(div_sub_x_7_n1050), .A4(div_sub_x_7_n1049), .A5(div_n_T_51_64_), 
        .A6(div_sub_x_7_n876), .Y(div_sub_x_7_n784) );
  INVX0_LVT div_sub_x_7_U657 ( .A(div_divisor_2_), .Y(div_sub_x_7_n783) );
  INVX0_LVT div_sub_x_7_U656 ( .A(div_sub_x_7_n906), .Y(div_sub_x_7_n782) );
  OA221X1_LVT div_sub_x_7_U655 ( .A1(1'b0), .A2(div_sub_x_7_n786), .A3(
        div_sub_x_7_n951), .A4(div_sub_x_7_n787), .A5(div_sub_x_7_n788), .Y(
        div_sub_x_7_n921) );
  OA221X1_LVT div_sub_x_7_U654 ( .A1(1'b0), .A2(div_sub_x_7_n798), .A3(
        div_sub_x_7_n920), .A4(div_sub_x_7_n799), .A5(div_sub_x_7_n800), .Y(
        div_sub_x_7_n917) );
  OA221X1_LVT div_sub_x_7_U653 ( .A1(1'b0), .A2(div_sub_x_7_n793), .A3(
        div_sub_x_7_n921), .A4(div_sub_x_7_n794), .A5(div_sub_x_7_n796), .Y(
        div_sub_x_7_n798) );
  OA221X1_LVT div_sub_x_7_U652 ( .A1(1'b0), .A2(div_sub_x_7_n805), .A3(
        div_sub_x_7_n1038), .A4(div_sub_x_7_n806), .A5(div_sub_x_7_n808), .Y(
        div_sub_x_7_n810) );
  OA221X1_LVT div_sub_x_7_U651 ( .A1(1'b0), .A2(div_sub_x_7_n811), .A3(
        div_sub_x_7_n1013), .A4(div_sub_x_7_n812), .A5(div_sub_x_7_n813), .Y(
        div_sub_x_7_n980) );
  OA221X1_LVT div_sub_x_7_U650 ( .A1(1'b0), .A2(div_sub_x_7_n823), .A3(
        div_sub_x_7_n1067), .A4(div_sub_x_7_n824), .A5(div_sub_x_7_n825), .Y(
        div_sub_x_7_n1037) );
  AO222X1_LVT div_sub_x_7_U649 ( .A1(div_sub_x_7_n815), .A2(div_sub_x_7_n817), 
        .A3(div_sub_x_7_n818), .A4(div_sub_x_7_n819), .A5(div_sub_x_7_n820), 
        .A6(1'b1), .Y(div_sub_x_7_n1041) );
  NAND3X0_LVT add_x_94_U264 ( .A1(add_x_94_n125), .A2(mem_reg_pc[3]), .A3(
        mem_reg_pc[4]), .Y(add_x_94_n272) );
  AND3X1_LVT add_x_94_U263 ( .A1(mem_reg_pc[5]), .A2(mem_reg_pc[6]), .A3(
        add_x_94_n258), .Y(add_x_94_n270) );
  NAND3X0_LVT add_x_94_U262 ( .A1(mem_reg_pc[7]), .A2(mem_reg_pc[8]), .A3(
        add_x_94_n270), .Y(add_x_94_n268) );
  AND2X1_LVT add_x_94_U261 ( .A1(mem_reg_pc[9]), .A2(add_x_94_n257), .Y(
        add_x_94_n309) );
  HADDX1_LVT add_x_94_U260 ( .A0(add_x_94_n309), .B0(mem_reg_pc[10]), .SO(
        io_imem_btb_update_bits_br_pc[10]) );
  AND3X1_LVT add_x_94_U259 ( .A1(add_x_94_n257), .A2(mem_reg_pc[9]), .A3(
        mem_reg_pc[10]), .Y(add_x_94_n308) );
  HADDX1_LVT add_x_94_U258 ( .A0(mem_reg_pc[11]), .B0(add_x_94_n308), .SO(
        io_imem_btb_update_bits_br_pc[11]) );
  AND4X1_LVT add_x_94_U257 ( .A1(add_x_94_n257), .A2(mem_reg_pc[9]), .A3(
        mem_reg_pc[10]), .A4(mem_reg_pc[11]), .Y(add_x_94_n307) );
  HADDX1_LVT add_x_94_U256 ( .A0(mem_reg_pc[12]), .B0(add_x_94_n307), .SO(
        io_imem_btb_update_bits_br_pc[12]) );
  AND4X1_LVT add_x_94_U255 ( .A1(mem_reg_pc[9]), .A2(mem_reg_pc[10]), .A3(
        mem_reg_pc[12]), .A4(mem_reg_pc[11]), .Y(add_x_94_n306) );
  NAND2X0_LVT add_x_94_U254 ( .A1(add_x_94_n257), .A2(add_x_94_n306), .Y(
        add_x_94_n305) );
  AO22X1_LVT add_x_94_U253 ( .A1(mem_reg_pc[13]), .A2(add_x_94_n305), .A3(
        add_x_94_n264), .A4(add_x_94_n256), .Y(
        io_imem_btb_update_bits_br_pc[13]) );
  AND2X1_LVT add_x_94_U252 ( .A1(add_x_94_n256), .A2(mem_reg_pc[13]), .Y(
        add_x_94_n304) );
  HADDX1_LVT add_x_94_U251 ( .A0(add_x_94_n304), .B0(mem_reg_pc[14]), .SO(
        io_imem_btb_update_bits_br_pc[14]) );
  AND3X1_LVT add_x_94_U250 ( .A1(mem_reg_pc[13]), .A2(mem_reg_pc[14]), .A3(
        add_x_94_n256), .Y(add_x_94_n302) );
  HADDX1_LVT add_x_94_U249 ( .A0(mem_reg_pc[15]), .B0(add_x_94_n302), .SO(
        io_imem_btb_update_bits_br_pc[15]) );
  AND4X1_LVT add_x_94_U248 ( .A1(mem_reg_pc[13]), .A2(mem_reg_pc[14]), .A3(
        mem_reg_pc[15]), .A4(add_x_94_n256), .Y(add_x_94_n303) );
  HADDX1_LVT add_x_94_U247 ( .A0(mem_reg_pc[16]), .B0(add_x_94_n303), .SO(
        io_imem_btb_update_bits_br_pc[16]) );
  NAND3X0_LVT add_x_94_U246 ( .A1(mem_reg_pc[15]), .A2(mem_reg_pc[16]), .A3(
        add_x_94_n302), .Y(add_x_94_n301) );
  AO22X1_LVT add_x_94_U245 ( .A1(mem_reg_pc[17]), .A2(add_x_94_n301), .A3(
        add_x_94_n263), .A4(add_x_94_n255), .Y(
        io_imem_btb_update_bits_br_pc[17]) );
  AND2X1_LVT add_x_94_U244 ( .A1(add_x_94_n255), .A2(mem_reg_pc[17]), .Y(
        add_x_94_n300) );
  HADDX1_LVT add_x_94_U243 ( .A0(add_x_94_n300), .B0(mem_reg_pc[18]), .SO(
        io_imem_btb_update_bits_br_pc[18]) );
  AND3X1_LVT add_x_94_U242 ( .A1(mem_reg_pc[17]), .A2(mem_reg_pc[18]), .A3(
        add_x_94_n255), .Y(add_x_94_n299) );
  HADDX1_LVT add_x_94_U241 ( .A0(mem_reg_pc[19]), .B0(add_x_94_n299), .SO(
        io_imem_btb_update_bits_br_pc[19]) );
  NAND2X0_LVT add_x_94_U240 ( .A1(mem_reg_pc[1]), .A2(n570), .Y(add_x_94_n267)
         );
  OA21X1_LVT add_x_94_U239 ( .A1(mem_reg_pc[1]), .A2(n570), .A3(add_x_94_n267), 
        .Y(io_imem_btb_update_bits_br_pc[1]) );
  AND4X1_LVT add_x_94_U238 ( .A1(mem_reg_pc[17]), .A2(mem_reg_pc[18]), .A3(
        mem_reg_pc[19]), .A4(add_x_94_n255), .Y(add_x_94_n298) );
  HADDX1_LVT add_x_94_U237 ( .A0(mem_reg_pc[20]), .B0(add_x_94_n298), .SO(
        io_imem_btb_update_bits_br_pc[20]) );
  AND4X1_LVT add_x_94_U236 ( .A1(mem_reg_pc[17]), .A2(mem_reg_pc[18]), .A3(
        mem_reg_pc[20]), .A4(mem_reg_pc[19]), .Y(add_x_94_n293) );
  AND2X1_LVT add_x_94_U235 ( .A1(add_x_94_n293), .A2(add_x_94_n255), .Y(
        add_x_94_n297) );
  HADDX1_LVT add_x_94_U234 ( .A0(mem_reg_pc[21]), .B0(add_x_94_n297), .SO(
        io_imem_btb_update_bits_br_pc[21]) );
  AND3X1_LVT add_x_94_U233 ( .A1(add_x_94_n293), .A2(mem_reg_pc[21]), .A3(
        add_x_94_n255), .Y(add_x_94_n296) );
  HADDX1_LVT add_x_94_U232 ( .A0(add_x_94_n296), .B0(mem_reg_pc[22]), .SO(
        io_imem_btb_update_bits_br_pc[22]) );
  AND2X1_LVT add_x_94_U231 ( .A1(mem_reg_pc[21]), .A2(mem_reg_pc[22]), .Y(
        add_x_94_n292) );
  AND3X1_LVT add_x_94_U230 ( .A1(add_x_94_n292), .A2(add_x_94_n293), .A3(
        add_x_94_n255), .Y(add_x_94_n295) );
  HADDX1_LVT add_x_94_U229 ( .A0(mem_reg_pc[23]), .B0(add_x_94_n295), .SO(
        io_imem_btb_update_bits_br_pc[23]) );
  AND4X1_LVT add_x_94_U228 ( .A1(mem_reg_pc[23]), .A2(add_x_94_n292), .A3(
        add_x_94_n293), .A4(add_x_94_n255), .Y(add_x_94_n294) );
  HADDX1_LVT add_x_94_U227 ( .A0(mem_reg_pc[24]), .B0(add_x_94_n294), .SO(
        io_imem_btb_update_bits_br_pc[24]) );
  AND4X1_LVT add_x_94_U226 ( .A1(mem_reg_pc[23]), .A2(mem_reg_pc[24]), .A3(
        add_x_94_n292), .A4(add_x_94_n293), .Y(add_x_94_n291) );
  NAND2X0_LVT add_x_94_U225 ( .A1(add_x_94_n291), .A2(add_x_94_n255), .Y(
        add_x_94_n290) );
  AO22X1_LVT add_x_94_U224 ( .A1(mem_reg_pc[25]), .A2(add_x_94_n290), .A3(
        add_x_94_n262), .A4(add_x_94_n254), .Y(
        io_imem_btb_update_bits_br_pc[25]) );
  AND2X1_LVT add_x_94_U223 ( .A1(add_x_94_n254), .A2(mem_reg_pc[25]), .Y(
        add_x_94_n289) );
  HADDX1_LVT add_x_94_U222 ( .A0(add_x_94_n289), .B0(mem_reg_pc[26]), .SO(
        io_imem_btb_update_bits_br_pc[26]) );
  AND3X1_LVT add_x_94_U221 ( .A1(mem_reg_pc[25]), .A2(mem_reg_pc[26]), .A3(
        add_x_94_n254), .Y(add_x_94_n288) );
  HADDX1_LVT add_x_94_U220 ( .A0(mem_reg_pc[27]), .B0(add_x_94_n288), .SO(
        io_imem_btb_update_bits_br_pc[27]) );
  AND4X1_LVT add_x_94_U219 ( .A1(mem_reg_pc[25]), .A2(mem_reg_pc[26]), .A3(
        mem_reg_pc[27]), .A4(add_x_94_n254), .Y(add_x_94_n287) );
  HADDX1_LVT add_x_94_U218 ( .A0(mem_reg_pc[28]), .B0(add_x_94_n287), .SO(
        io_imem_btb_update_bits_br_pc[28]) );
  AND4X1_LVT add_x_94_U217 ( .A1(mem_reg_pc[25]), .A2(mem_reg_pc[26]), .A3(
        mem_reg_pc[28]), .A4(mem_reg_pc[27]), .Y(add_x_94_n282) );
  NAND2X0_LVT add_x_94_U216 ( .A1(add_x_94_n282), .A2(add_x_94_n254), .Y(
        add_x_94_n286) );
  AO22X1_LVT add_x_94_U215 ( .A1(mem_reg_pc[29]), .A2(add_x_94_n286), .A3(
        add_x_94_n261), .A4(add_x_94_n252), .Y(
        io_imem_btb_update_bits_br_pc[29]) );
  AND2X1_LVT add_x_94_U214 ( .A1(add_x_94_n252), .A2(mem_reg_pc[29]), .Y(
        add_x_94_n285) );
  HADDX1_LVT add_x_94_U213 ( .A0(add_x_94_n285), .B0(mem_reg_pc[30]), .SO(
        io_imem_btb_update_bits_br_pc[30]) );
  AND3X1_LVT add_x_94_U212 ( .A1(mem_reg_pc[29]), .A2(mem_reg_pc[30]), .A3(
        add_x_94_n252), .Y(add_x_94_n284) );
  HADDX1_LVT add_x_94_U211 ( .A0(mem_reg_pc[31]), .B0(add_x_94_n284), .SO(
        io_imem_btb_update_bits_br_pc[31]) );
  AND4X1_LVT add_x_94_U210 ( .A1(mem_reg_pc[31]), .A2(mem_reg_pc[29]), .A3(
        mem_reg_pc[30]), .A4(add_x_94_n252), .Y(add_x_94_n283) );
  HADDX1_LVT add_x_94_U209 ( .A0(mem_reg_pc[32]), .B0(add_x_94_n283), .SO(
        io_imem_btb_update_bits_br_pc[32]) );
  AND4X1_LVT add_x_94_U208 ( .A1(mem_reg_pc[29]), .A2(mem_reg_pc[30]), .A3(
        add_x_94_n282), .A4(add_x_94_n254), .Y(add_x_94_n281) );
  NAND3X0_LVT add_x_94_U207 ( .A1(mem_reg_pc[32]), .A2(mem_reg_pc[31]), .A3(
        add_x_94_n281), .Y(add_x_94_n280) );
  AO22X1_LVT add_x_94_U206 ( .A1(add_x_94_n253), .A2(add_x_94_n260), .A3(
        add_x_94_n280), .A4(mem_reg_pc[33]), .Y(
        io_imem_btb_update_bits_br_pc[33]) );
  AND2X1_LVT add_x_94_U205 ( .A1(mem_reg_pc[33]), .A2(add_x_94_n253), .Y(
        add_x_94_n279) );
  HADDX1_LVT add_x_94_U204 ( .A0(add_x_94_n279), .B0(mem_reg_pc[34]), .SO(
        io_imem_btb_update_bits_br_pc[34]) );
  AND3X1_LVT add_x_94_U203 ( .A1(add_x_94_n253), .A2(mem_reg_pc[34]), .A3(
        mem_reg_pc[33]), .Y(add_x_94_n278) );
  HADDX1_LVT add_x_94_U202 ( .A0(add_x_94_n278), .B0(mem_reg_pc[35]), .SO(
        io_imem_btb_update_bits_br_pc[35]) );
  AND4X1_LVT add_x_94_U201 ( .A1(mem_reg_pc[34]), .A2(add_x_94_n253), .A3(
        mem_reg_pc[33]), .A4(mem_reg_pc[35]), .Y(add_x_94_n277) );
  HADDX1_LVT add_x_94_U200 ( .A0(mem_reg_pc[36]), .B0(add_x_94_n277), .SO(
        io_imem_btb_update_bits_br_pc[36]) );
  AND4X1_LVT add_x_94_U199 ( .A1(mem_reg_pc[34]), .A2(mem_reg_pc[33]), .A3(
        mem_reg_pc[35]), .A4(mem_reg_pc[36]), .Y(add_x_94_n276) );
  AND2X1_LVT add_x_94_U198 ( .A1(add_x_94_n253), .A2(add_x_94_n276), .Y(
        add_x_94_n275) );
  HADDX1_LVT add_x_94_U197 ( .A0(mem_reg_pc[37]), .B0(add_x_94_n275), .SO(
        io_imem_btb_update_bits_br_pc[37]) );
  AND2X1_LVT add_x_94_U196 ( .A1(add_x_94_n275), .A2(mem_reg_pc[37]), .Y(
        add_x_94_n274) );
  HADDX1_LVT add_x_94_U195 ( .A0(add_x_94_n274), .B0(mem_reg_pc[38]), .SO(
        io_imem_btb_update_bits_br_pc[38]) );
  HADDX1_LVT add_x_94_U194 ( .A0(add_x_94_n125), .B0(mem_reg_pc[3]), .SO(
        io_imem_btb_update_bits_br_pc[3]) );
  AND2X1_LVT add_x_94_U193 ( .A1(add_x_94_n125), .A2(mem_reg_pc[3]), .Y(
        add_x_94_n273) );
  HADDX1_LVT add_x_94_U192 ( .A0(mem_reg_pc[4]), .B0(add_x_94_n273), .SO(
        io_imem_btb_update_bits_br_pc[4]) );
  AO22X1_LVT add_x_94_U191 ( .A1(mem_reg_pc[5]), .A2(add_x_94_n272), .A3(
        add_x_94_n266), .A4(add_x_94_n258), .Y(
        io_imem_btb_update_bits_br_pc[5]) );
  AND2X1_LVT add_x_94_U190 ( .A1(add_x_94_n258), .A2(mem_reg_pc[5]), .Y(
        add_x_94_n271) );
  HADDX1_LVT add_x_94_U189 ( .A0(add_x_94_n271), .B0(mem_reg_pc[6]), .SO(
        io_imem_btb_update_bits_br_pc[6]) );
  HADDX1_LVT add_x_94_U188 ( .A0(mem_reg_pc[7]), .B0(add_x_94_n270), .SO(
        io_imem_btb_update_bits_br_pc[7]) );
  AND2X1_LVT add_x_94_U187 ( .A1(mem_reg_pc[7]), .A2(add_x_94_n270), .Y(
        add_x_94_n269) );
  HADDX1_LVT add_x_94_U186 ( .A0(mem_reg_pc[8]), .B0(add_x_94_n269), .SO(
        io_imem_btb_update_bits_br_pc[8]) );
  AO22X1_LVT add_x_94_U185 ( .A1(add_x_94_n257), .A2(add_x_94_n265), .A3(
        add_x_94_n268), .A4(mem_reg_pc[9]), .Y(
        io_imem_btb_update_bits_br_pc[9]) );
  INVX1_LVT add_x_94_U184 ( .A(mem_reg_pc[5]), .Y(add_x_94_n266) );
  INVX1_LVT add_x_94_U183 ( .A(mem_reg_pc[9]), .Y(add_x_94_n265) );
  INVX1_LVT add_x_94_U182 ( .A(mem_reg_pc[13]), .Y(add_x_94_n264) );
  INVX1_LVT add_x_94_U181 ( .A(mem_reg_pc[17]), .Y(add_x_94_n263) );
  INVX1_LVT add_x_94_U180 ( .A(mem_reg_pc[25]), .Y(add_x_94_n262) );
  INVX1_LVT add_x_94_U179 ( .A(mem_reg_pc[29]), .Y(add_x_94_n261) );
  INVX1_LVT add_x_94_U178 ( .A(mem_reg_pc[33]), .Y(add_x_94_n260) );
  INVX1_LVT add_x_94_U177 ( .A(add_x_94_n267), .Y(add_x_94_n259) );
  INVX1_LVT add_x_94_U176 ( .A(add_x_94_n272), .Y(add_x_94_n258) );
  INVX1_LVT add_x_94_U175 ( .A(add_x_94_n305), .Y(add_x_94_n256) );
  INVX1_LVT add_x_94_U174 ( .A(add_x_94_n290), .Y(add_x_94_n254) );
  INVX1_LVT add_x_94_U173 ( .A(add_x_94_n280), .Y(add_x_94_n253) );
  INVX1_LVT add_x_94_U172 ( .A(add_x_94_n286), .Y(add_x_94_n252) );
  INVX1_LVT add_x_94_U171 ( .A(add_x_94_n268), .Y(add_x_94_n257) );
  INVX1_LVT add_x_94_U170 ( .A(add_x_94_n301), .Y(add_x_94_n255) );
  HADDX1_LVT add_x_94_U160 ( .A0(mem_reg_pc[2]), .B0(add_x_94_n259), .C1(
        add_x_94_n125), .SO(io_imem_btb_update_bits_br_pc[2]) );
  AND2X1_LVT add_x_5_U477 ( .A1(mem_reg_pc[3]), .A2(n_T_914[3]), .Y(
        add_x_5_n421) );
  OR2X1_LVT add_x_5_U476 ( .A1(n_T_914[4]), .A2(mem_reg_pc[4]), .Y(
        add_x_5_n504) );
  AO22X1_LVT add_x_5_U475 ( .A1(n_T_914[4]), .A2(mem_reg_pc[4]), .A3(
        add_x_5_n421), .A4(add_x_5_n504), .Y(add_x_5_n503) );
  OR2X1_LVT add_x_5_U474 ( .A1(mem_reg_pc[3]), .A2(n_T_914[3]), .Y(
        add_x_5_n420) );
  OA222X1_LVT add_x_5_U473 ( .A1(add_x_5_n503), .A2(add_x_5_n246), .A3(
        add_x_5_n503), .A4(add_x_5_n504), .A5(add_x_5_n503), .A6(add_x_5_n420), 
        .Y(add_x_5_n415) );
  OA22X1_LVT add_x_5_U472 ( .A1(n_T_914[6]), .A2(mem_reg_pc[6]), .A3(
        n_T_914[5]), .A4(mem_reg_pc[5]), .Y(add_x_5_n414) );
  AND2X1_LVT add_x_5_U471 ( .A1(n_T_914[5]), .A2(mem_reg_pc[5]), .Y(
        add_x_5_n418) );
  AND2X1_LVT add_x_5_U470 ( .A1(n_T_914[7]), .A2(mem_reg_pc[7]), .Y(
        add_x_5_n413) );
  AND2X1_LVT add_x_5_U469 ( .A1(mem_reg_pc[9]), .A2(n_T_914[9]), .Y(
        add_x_5_n501) );
  AO221X1_LVT add_x_5_U468 ( .A1(add_x_5_n410), .A2(mem_reg_pc[9]), .A3(
        add_x_5_n410), .A4(n_T_914[9]), .A5(add_x_5_n501), .Y(add_x_5_n502) );
  FADDX1_LVT add_x_5_U467 ( .A(n_T_914[10]), .B(mem_reg_pc[10]), .CI(
        add_x_5_n502), .S(mem_br_target_10_) );
  OA22X1_LVT add_x_5_U466 ( .A1(mem_reg_pc[9]), .A2(n_T_914[9]), .A3(
        n_T_914[10]), .A4(mem_reg_pc[10]), .Y(add_x_5_n498) );
  AO21X1_LVT add_x_5_U465 ( .A1(add_x_5_n498), .A2(add_x_5_n410), .A3(
        add_x_5_n497), .Y(add_x_5_n500) );
  FADDX1_LVT add_x_5_U464 ( .A(n_T_914[11]), .B(mem_reg_pc[11]), .CI(
        add_x_5_n500), .S(mem_br_target_11_) );
  AND2X1_LVT add_x_5_U463 ( .A1(n_T_914[11]), .A2(mem_reg_pc[11]), .Y(
        add_x_5_n494) );
  OA22X1_LVT add_x_5_U462 ( .A1(add_x_5_n494), .A2(add_x_5_n500), .A3(
        n_T_914[11]), .A4(mem_reg_pc[11]), .Y(add_x_5_n499) );
  FADDX1_LVT add_x_5_U461 ( .A(n_T_914[12]), .B(mem_reg_pc[12]), .CI(
        add_x_5_n499), .S(mem_br_target_12_) );
  OA22X1_LVT add_x_5_U460 ( .A1(n_T_914[12]), .A2(mem_reg_pc[12]), .A3(
        n_T_914[11]), .A4(mem_reg_pc[11]), .Y(add_x_5_n496) );
  AND2X1_LVT add_x_5_U459 ( .A1(add_x_5_n496), .A2(add_x_5_n498), .Y(
        add_x_5_n484) );
  OR2X1_LVT add_x_5_U458 ( .A1(mem_reg_pc[12]), .A2(n_T_914[12]), .Y(
        add_x_5_n495) );
  AO222X1_LVT add_x_5_U457 ( .A1(n_T_914[12]), .A2(mem_reg_pc[12]), .A3(
        add_x_5_n494), .A4(add_x_5_n495), .A5(add_x_5_n496), .A6(add_x_5_n497), 
        .Y(add_x_5_n486) );
  AO21X1_LVT add_x_5_U456 ( .A1(add_x_5_n484), .A2(add_x_5_n410), .A3(
        add_x_5_n486), .Y(add_x_5_n491) );
  FADDX1_LVT add_x_5_U455 ( .A(n_T_914[13]), .B(mem_reg_pc[13]), .CI(
        add_x_5_n491), .S(mem_br_target_13_) );
  AND2X1_LVT add_x_5_U454 ( .A1(n_T_914[13]), .A2(mem_reg_pc[13]), .Y(
        add_x_5_n492) );
  OA22X1_LVT add_x_5_U453 ( .A1(add_x_5_n492), .A2(add_x_5_n491), .A3(
        n_T_914[13]), .A4(mem_reg_pc[13]), .Y(add_x_5_n493) );
  FADDX1_LVT add_x_5_U452 ( .A(n_T_914[14]), .B(mem_reg_pc[14]), .CI(
        add_x_5_n493), .S(mem_br_target_14_) );
  OA22X1_LVT add_x_5_U451 ( .A1(n_T_914[14]), .A2(mem_reg_pc[14]), .A3(
        n_T_914[13]), .A4(mem_reg_pc[13]), .Y(add_x_5_n488) );
  AO21X1_LVT add_x_5_U450 ( .A1(add_x_5_n488), .A2(add_x_5_n491), .A3(
        add_x_5_n485), .Y(add_x_5_n490) );
  FADDX1_LVT add_x_5_U449 ( .A(n_T_914[15]), .B(mem_reg_pc[15]), .CI(
        add_x_5_n490), .S(mem_br_target_15_) );
  AND2X1_LVT add_x_5_U448 ( .A1(n_T_914[15]), .A2(mem_reg_pc[15]), .Y(
        add_x_5_n487) );
  OA22X1_LVT add_x_5_U447 ( .A1(add_x_5_n487), .A2(add_x_5_n490), .A3(
        n_T_914[15]), .A4(mem_reg_pc[15]), .Y(add_x_5_n489) );
  FADDX1_LVT add_x_5_U446 ( .A(n_T_914[16]), .B(mem_reg_pc[16]), .CI(
        add_x_5_n489), .S(mem_br_target_16_) );
  FADDX1_LVT add_x_5_U445 ( .A(n_T_914[17]), .B(mem_reg_pc[17]), .CI(
        add_x_5_n440), .S(mem_br_target_17_) );
  AND2X1_LVT add_x_5_U444 ( .A1(n_T_914[17]), .A2(mem_reg_pc[17]), .Y(
        add_x_5_n482) );
  OA22X1_LVT add_x_5_U443 ( .A1(n_T_914[17]), .A2(mem_reg_pc[17]), .A3(
        add_x_5_n482), .A4(add_x_5_n440), .Y(add_x_5_n483) );
  FADDX1_LVT add_x_5_U442 ( .A(n_T_914[18]), .B(mem_reg_pc[18]), .CI(
        add_x_5_n483), .S(mem_br_target_18_) );
  OA22X1_LVT add_x_5_U441 ( .A1(n_T_914[18]), .A2(mem_reg_pc[18]), .A3(
        n_T_914[17]), .A4(mem_reg_pc[17]), .Y(add_x_5_n479) );
  AO21X1_LVT add_x_5_U440 ( .A1(add_x_5_n479), .A2(add_x_5_n440), .A3(
        add_x_5_n478), .Y(add_x_5_n481) );
  FADDX1_LVT add_x_5_U439 ( .A(n_T_914[19]), .B(mem_reg_pc[19]), .CI(
        add_x_5_n481), .S(mem_br_target_19_) );
  NAND2X0_LVT add_x_5_U438 ( .A1(mem_reg_pc[1]), .A2(n_T_914[1]), .Y(
        add_x_5_n409) );
  OA21X1_LVT add_x_5_U437 ( .A1(mem_reg_pc[1]), .A2(n_T_914[1]), .A3(
        add_x_5_n409), .Y(mem_br_target_1_) );
  AND2X1_LVT add_x_5_U436 ( .A1(n_T_914[19]), .A2(mem_reg_pc[19]), .Y(
        add_x_5_n475) );
  AO221X1_LVT add_x_5_U435 ( .A1(add_x_5_n481), .A2(n_T_914[19]), .A3(
        add_x_5_n481), .A4(mem_reg_pc[19]), .A5(add_x_5_n475), .Y(add_x_5_n480) );
  FADDX1_LVT add_x_5_U434 ( .A(add_x_5_n403), .B(mem_reg_pc[20]), .CI(
        add_x_5_n480), .S(mem_br_target_20_) );
  OA22X1_LVT add_x_5_U433 ( .A1(n9427), .A2(mem_reg_pc[20]), .A3(n_T_914[19]), 
        .A4(mem_reg_pc[19]), .Y(add_x_5_n477) );
  AND2X1_LVT add_x_5_U432 ( .A1(add_x_5_n477), .A2(add_x_5_n479), .Y(
        add_x_5_n467) );
  OR2X1_LVT add_x_5_U431 ( .A1(mem_reg_pc[20]), .A2(add_x_5_n403), .Y(
        add_x_5_n476) );
  AO222X1_LVT add_x_5_U430 ( .A1(n9427), .A2(mem_reg_pc[20]), .A3(add_x_5_n475), .A4(add_x_5_n476), .A5(add_x_5_n477), .A6(add_x_5_n478), .Y(add_x_5_n465) );
  AO21X1_LVT add_x_5_U429 ( .A1(add_x_5_n467), .A2(add_x_5_n440), .A3(
        add_x_5_n465), .Y(add_x_5_n472) );
  FADDX1_LVT add_x_5_U428 ( .A(n9427), .B(mem_reg_pc[21]), .CI(add_x_5_n472), 
        .S(mem_br_target_21_) );
  OR2X1_LVT add_x_5_U427 ( .A1(add_x_5_n403), .A2(mem_reg_pc[21]), .Y(
        add_x_5_n474) );
  AO22X1_LVT add_x_5_U426 ( .A1(add_x_5_n403), .A2(mem_reg_pc[21]), .A3(
        add_x_5_n472), .A4(add_x_5_n474), .Y(add_x_5_n473) );
  FADDX1_LVT add_x_5_U425 ( .A(n9427), .B(mem_reg_pc[22]), .CI(add_x_5_n473), 
        .S(mem_br_target_22_) );
  OA21X1_LVT add_x_5_U424 ( .A1(mem_reg_pc[22]), .A2(mem_reg_pc[21]), .A3(
        add_x_5_n403), .Y(add_x_5_n466) );
  AO21X1_LVT add_x_5_U423 ( .A1(mem_reg_pc[22]), .A2(mem_reg_pc[21]), .A3(
        add_x_5_n403), .Y(add_x_5_n468) );
  OA21X1_LVT add_x_5_U422 ( .A1(add_x_5_n472), .A2(add_x_5_n466), .A3(
        add_x_5_n468), .Y(add_x_5_n470) );
  FADDX1_LVT add_x_5_U421 ( .A(add_x_5_n403), .B(mem_reg_pc[23]), .CI(
        add_x_5_n470), .S(mem_br_target_23_) );
  OR2X1_LVT add_x_5_U420 ( .A1(add_x_5_n403), .A2(mem_reg_pc[23]), .Y(
        add_x_5_n471) );
  AO22X1_LVT add_x_5_U419 ( .A1(n9427), .A2(mem_reg_pc[23]), .A3(add_x_5_n470), 
        .A4(add_x_5_n471), .Y(add_x_5_n469) );
  FADDX1_LVT add_x_5_U418 ( .A(add_x_5_n403), .B(mem_reg_pc[24]), .CI(
        add_x_5_n469), .S(mem_br_target_24_) );
  OA221X1_LVT add_x_5_U417 ( .A1(add_x_5_n403), .A2(mem_reg_pc[23]), .A3(
        add_x_5_n403), .A4(mem_reg_pc[24]), .A5(add_x_5_n468), .Y(add_x_5_n464) );
  AND2X1_LVT add_x_5_U416 ( .A1(add_x_5_n467), .A2(add_x_5_n464), .Y(
        add_x_5_n441) );
  AO21X1_LVT add_x_5_U415 ( .A1(add_x_5_n441), .A2(add_x_5_n440), .A3(
        add_x_5_n450), .Y(add_x_5_n456) );
  FADDX1_LVT add_x_5_U414 ( .A(n9427), .B(mem_reg_pc[25]), .CI(add_x_5_n456), 
        .S(mem_br_target_25_) );
  OR2X1_LVT add_x_5_U413 ( .A1(add_x_5_n403), .A2(mem_reg_pc[25]), .Y(
        add_x_5_n463) );
  AO22X1_LVT add_x_5_U412 ( .A1(add_x_5_n403), .A2(mem_reg_pc[25]), .A3(
        add_x_5_n456), .A4(add_x_5_n463), .Y(add_x_5_n462) );
  FADDX1_LVT add_x_5_U411 ( .A(n9427), .B(mem_reg_pc[26]), .CI(add_x_5_n462), 
        .S(mem_br_target_26_) );
  OA21X1_LVT add_x_5_U410 ( .A1(mem_reg_pc[26]), .A2(mem_reg_pc[25]), .A3(
        n9427), .Y(add_x_5_n458) );
  AO21X1_LVT add_x_5_U409 ( .A1(mem_reg_pc[26]), .A2(mem_reg_pc[25]), .A3(
        add_x_5_n403), .Y(add_x_5_n457) );
  OA21X1_LVT add_x_5_U408 ( .A1(add_x_5_n456), .A2(add_x_5_n458), .A3(
        add_x_5_n457), .Y(add_x_5_n460) );
  FADDX1_LVT add_x_5_U407 ( .A(n9427), .B(mem_reg_pc[27]), .CI(add_x_5_n460), 
        .S(mem_br_target_27_) );
  OR2X1_LVT add_x_5_U406 ( .A1(add_x_5_n403), .A2(mem_reg_pc[27]), .Y(
        add_x_5_n461) );
  AO22X1_LVT add_x_5_U405 ( .A1(n9427), .A2(mem_reg_pc[27]), .A3(add_x_5_n460), 
        .A4(add_x_5_n461), .Y(add_x_5_n459) );
  FADDX1_LVT add_x_5_U404 ( .A(n9427), .B(mem_reg_pc[28]), .CI(add_x_5_n459), 
        .S(mem_br_target_28_) );
  AO221X1_LVT add_x_5_U403 ( .A1(add_x_5_n403), .A2(mem_reg_pc[27]), .A3(
        add_x_5_n403), .A4(mem_reg_pc[28]), .A5(add_x_5_n458), .Y(add_x_5_n448) );
  OA221X1_LVT add_x_5_U402 ( .A1(add_x_5_n403), .A2(mem_reg_pc[27]), .A3(n9427), .A4(mem_reg_pc[28]), .A5(add_x_5_n457), .Y(add_x_5_n444) );
  OA21X1_LVT add_x_5_U401 ( .A1(add_x_5_n456), .A2(add_x_5_n448), .A3(
        add_x_5_n444), .Y(add_x_5_n453) );
  FADDX1_LVT add_x_5_U400 ( .A(n9427), .B(mem_reg_pc[29]), .CI(add_x_5_n453), 
        .S(mem_br_target_29_) );
  OR2X1_LVT add_x_5_U399 ( .A1(add_x_5_n403), .A2(mem_reg_pc[29]), .Y(
        add_x_5_n455) );
  AO22X1_LVT add_x_5_U398 ( .A1(add_x_5_n403), .A2(mem_reg_pc[29]), .A3(
        add_x_5_n453), .A4(add_x_5_n455), .Y(add_x_5_n454) );
  FADDX1_LVT add_x_5_U397 ( .A(n9427), .B(mem_reg_pc[30]), .CI(add_x_5_n454), 
        .S(mem_br_target_30_) );
  OA21X1_LVT add_x_5_U396 ( .A1(mem_reg_pc[30]), .A2(mem_reg_pc[29]), .A3(
        add_x_5_n403), .Y(add_x_5_n447) );
  AO21X1_LVT add_x_5_U395 ( .A1(mem_reg_pc[30]), .A2(mem_reg_pc[29]), .A3(
        n9427), .Y(add_x_5_n443) );
  OA21X1_LVT add_x_5_U394 ( .A1(add_x_5_n453), .A2(add_x_5_n447), .A3(
        add_x_5_n443), .Y(add_x_5_n452) );
  FADDX1_LVT add_x_5_U393 ( .A(add_x_5_n403), .B(mem_reg_pc[31]), .CI(
        add_x_5_n452), .S(mem_br_target_31_) );
  OR2X1_LVT add_x_5_U392 ( .A1(n9427), .A2(mem_reg_pc[31]), .Y(add_x_5_n445)
         );
  AO22X1_LVT add_x_5_U391 ( .A1(n9427), .A2(mem_reg_pc[31]), .A3(add_x_5_n452), 
        .A4(add_x_5_n445), .Y(add_x_5_n451) );
  FADDX1_LVT add_x_5_U390 ( .A(add_x_5_n403), .B(mem_reg_pc[32]), .CI(
        add_x_5_n451), .S(mem_br_target_32_) );
  AO221X1_LVT add_x_5_U389 ( .A1(n9427), .A2(mem_reg_pc[31]), .A3(n9427), .A4(
        mem_reg_pc[32]), .A5(add_x_5_n450), .Y(add_x_5_n449) );
  OR3X1_LVT add_x_5_U388 ( .A1(add_x_5_n447), .A2(add_x_5_n448), .A3(
        add_x_5_n449), .Y(add_x_5_n439) );
  OR2X1_LVT add_x_5_U387 ( .A1(n9427), .A2(mem_reg_pc[32]), .Y(add_x_5_n446)
         );
  AND4X1_LVT add_x_5_U386 ( .A1(add_x_5_n443), .A2(add_x_5_n444), .A3(
        add_x_5_n445), .A4(add_x_5_n446), .Y(add_x_5_n442) );
  FADDX1_LVT add_x_5_U385 ( .A(add_x_5_n403), .B(mem_reg_pc[33]), .CI(
        add_x_5_n429), .S(mem_br_target_33_) );
  OR2X1_LVT add_x_5_U384 ( .A1(add_x_5_n403), .A2(mem_reg_pc[33]), .Y(
        add_x_5_n438) );
  AO22X1_LVT add_x_5_U383 ( .A1(add_x_5_n403), .A2(mem_reg_pc[33]), .A3(
        add_x_5_n429), .A4(add_x_5_n438), .Y(add_x_5_n437) );
  FADDX1_LVT add_x_5_U382 ( .A(n9427), .B(mem_reg_pc[34]), .CI(add_x_5_n437), 
        .S(mem_br_target_34_) );
  AO21X1_LVT add_x_5_U381 ( .A1(mem_reg_pc[33]), .A2(mem_reg_pc[34]), .A3(
        n9427), .Y(add_x_5_n433) );
  OA21X1_LVT add_x_5_U380 ( .A1(mem_reg_pc[33]), .A2(mem_reg_pc[34]), .A3(
        n9427), .Y(add_x_5_n432) );
  AO21X1_LVT add_x_5_U379 ( .A1(add_x_5_n433), .A2(add_x_5_n429), .A3(
        add_x_5_n432), .Y(add_x_5_n436) );
  FADDX1_LVT add_x_5_U378 ( .A(add_x_5_n403), .B(mem_reg_pc[35]), .CI(
        add_x_5_n436), .S(mem_br_target_35_) );
  AND2X1_LVT add_x_5_U377 ( .A1(add_x_5_n403), .A2(mem_reg_pc[35]), .Y(
        add_x_5_n435) );
  OA22X1_LVT add_x_5_U376 ( .A1(add_x_5_n435), .A2(add_x_5_n436), .A3(n9427), 
        .A4(mem_reg_pc[35]), .Y(add_x_5_n434) );
  FADDX1_LVT add_x_5_U375 ( .A(add_x_5_n403), .B(add_x_5_n434), .CI(
        mem_reg_pc[36]), .S(mem_br_target_36_) );
  OA221X1_LVT add_x_5_U374 ( .A1(n9427), .A2(mem_reg_pc[35]), .A3(n9427), .A4(
        mem_reg_pc[36]), .A5(add_x_5_n433), .Y(add_x_5_n427) );
  AO221X1_LVT add_x_5_U373 ( .A1(n9427), .A2(mem_reg_pc[35]), .A3(n9427), .A4(
        mem_reg_pc[36]), .A5(add_x_5_n432), .Y(add_x_5_n430) );
  AO21X1_LVT add_x_5_U372 ( .A1(add_x_5_n427), .A2(add_x_5_n429), .A3(
        add_x_5_n430), .Y(add_x_5_n431) );
  FADDX1_LVT add_x_5_U371 ( .A(n9427), .B(mem_reg_pc[37]), .CI(add_x_5_n431), 
        .S(mem_br_target_37_) );
  AOI21X1_LVT add_x_5_U370 ( .A1(n9427), .A2(mem_reg_pc[37]), .A3(add_x_5_n430), .Y(add_x_5_n423) );
  OR2X1_LVT add_x_5_U369 ( .A1(mem_reg_pc[37]), .A2(add_x_5_n403), .Y(
        add_x_5_n428) );
  NAND3X0_LVT add_x_5_U368 ( .A1(add_x_5_n427), .A2(add_x_5_n428), .A3(
        add_x_5_n429), .Y(add_x_5_n424) );
  NAND2X0_LVT add_x_5_U367 ( .A1(add_x_5_n423), .A2(add_x_5_n424), .Y(
        add_x_5_n426) );
  FADDX1_LVT add_x_5_U366 ( .A(add_x_5_n403), .B(mem_reg_pc[38]), .CI(
        add_x_5_n426), .S(mem_br_target_38_) );
  NAND2X0_LVT add_x_5_U365 ( .A1(n9427), .A2(mem_reg_pc[38]), .Y(add_x_5_n425)
         );
  FADDX1_LVT add_x_5_U364 ( .A(add_x_5_n422), .B(mem_reg_pc[39]), .CI(
        add_x_5_n404), .S(mem_br_target_39_) );
  FADDX1_LVT add_x_5_U363 ( .A(add_x_5_n246), .B(mem_reg_pc[3]), .CI(
        n_T_914[3]), .S(mem_br_target_3_) );
  AO21X1_LVT add_x_5_U362 ( .A1(add_x_5_n246), .A2(add_x_5_n420), .A3(
        add_x_5_n421), .Y(add_x_5_n419) );
  FADDX1_LVT add_x_5_U361 ( .A(n_T_914[4]), .B(mem_reg_pc[4]), .CI(
        add_x_5_n419), .S(mem_br_target_4_) );
  FADDX1_LVT add_x_5_U360 ( .A(add_x_5_n415), .B(n_T_914[5]), .CI(
        mem_reg_pc[5]), .S(mem_br_target_5_) );
  OA22X1_LVT add_x_5_U359 ( .A1(add_x_5_n415), .A2(add_x_5_n418), .A3(
        n_T_914[5]), .A4(mem_reg_pc[5]), .Y(add_x_5_n417) );
  FADDX1_LVT add_x_5_U358 ( .A(n_T_914[6]), .B(mem_reg_pc[6]), .CI(
        add_x_5_n417), .S(mem_br_target_6_) );
  AO21X1_LVT add_x_5_U357 ( .A1(add_x_5_n414), .A2(add_x_5_n415), .A3(
        add_x_5_n416), .Y(add_x_5_n412) );
  FADDX1_LVT add_x_5_U356 ( .A(n_T_914[7]), .B(mem_reg_pc[7]), .CI(
        add_x_5_n412), .S(mem_br_target_7_) );
  AO221X1_LVT add_x_5_U355 ( .A1(add_x_5_n412), .A2(n_T_914[7]), .A3(
        add_x_5_n412), .A4(mem_reg_pc[7]), .A5(add_x_5_n413), .Y(add_x_5_n411)
         );
  FADDX1_LVT add_x_5_U354 ( .A(n_T_914[8]), .B(mem_reg_pc[8]), .CI(
        add_x_5_n411), .S(mem_br_target_8_) );
  FADDX1_LVT add_x_5_U353 ( .A(mem_reg_pc[9]), .B(n_T_914[9]), .CI(
        add_x_5_n410), .S(mem_br_target_9_) );
  INVX1_LVT add_x_5_U352 ( .A(add_x_5_n409), .Y(add_x_5_n408) );
  NAND2X0_LVT add_x_5_U351 ( .A1(add_x_5_n402), .A2(add_x_5_n407), .Y(
        add_x_5_n406) );
  AND2X1_LVT add_x_5_U350 ( .A1(add_x_5_n425), .A2(add_x_5_n423), .Y(
        add_x_5_n405) );
  AND2X1_LVT add_x_5_U349 ( .A1(add_x_5_n405), .A2(add_x_5_n406), .Y(
        add_x_5_n422) );
  OR2X1_LVT add_x_5_U348 ( .A1(add_x_5_n403), .A2(mem_reg_pc[38]), .Y(
        add_x_5_n402) );
  NBUFFX2_LVT add_x_5_U347 ( .A(n9427), .Y(add_x_5_n403) );
  OA221X1_LVT add_x_5_U346 ( .A1(add_x_5_n439), .A2(add_x_5_n440), .A3(
        add_x_5_n439), .A4(add_x_5_n441), .A5(add_x_5_n442), .Y(add_x_5_n429)
         );
  INVX0_LVT add_x_5_U345 ( .A(add_x_5_n424), .Y(add_x_5_n407) );
  INVX1_LVT add_x_5_U344 ( .A(n9427), .Y(add_x_5_n404) );
  AO222X1_LVT add_x_5_U343 ( .A1(n_T_914[6]), .A2(mem_reg_pc[6]), .A3(
        n_T_914[6]), .A4(add_x_5_n418), .A5(mem_reg_pc[6]), .A6(add_x_5_n418), 
        .Y(add_x_5_n416) );
  AO222X1_LVT add_x_5_U342 ( .A1(n_T_914[10]), .A2(mem_reg_pc[10]), .A3(
        n_T_914[10]), .A4(add_x_5_n501), .A5(mem_reg_pc[10]), .A6(add_x_5_n501), .Y(add_x_5_n497) );
  AO221X1_LVT add_x_5_U341 ( .A1(add_x_5_n403), .A2(mem_reg_pc[23]), .A3(
        add_x_5_n403), .A4(mem_reg_pc[24]), .A5(add_x_5_n401), .Y(add_x_5_n450) );
  AO21X1_LVT add_x_5_U340 ( .A1(add_x_5_n465), .A2(add_x_5_n464), .A3(
        add_x_5_n466), .Y(add_x_5_n401) );
  AO222X1_LVT add_x_5_U339 ( .A1(n_T_914[18]), .A2(mem_reg_pc[18]), .A3(
        n_T_914[18]), .A4(add_x_5_n482), .A5(mem_reg_pc[18]), .A6(add_x_5_n482), .Y(add_x_5_n478) );
  AO222X1_LVT add_x_5_U338 ( .A1(n_T_914[14]), .A2(mem_reg_pc[14]), .A3(
        n_T_914[14]), .A4(add_x_5_n492), .A5(mem_reg_pc[14]), .A6(add_x_5_n492), .Y(add_x_5_n485) );
  AO222X1_LVT add_x_5_U337 ( .A1(add_x_5_n398), .A2(add_x_5_n399), .A3(
        add_x_5_n400), .A4(add_x_5_n413), .A5(mem_reg_pc[8]), .A6(n_T_914[8]), 
        .Y(add_x_5_n410) );
  OR2X1_LVT add_x_5_U336 ( .A1(n_T_914[8]), .A2(mem_reg_pc[8]), .Y(
        add_x_5_n400) );
  OA22X1_LVT add_x_5_U335 ( .A1(n_T_914[7]), .A2(mem_reg_pc[7]), .A3(
        n_T_914[8]), .A4(mem_reg_pc[8]), .Y(add_x_5_n399) );
  AO21X1_LVT add_x_5_U334 ( .A1(add_x_5_n415), .A2(add_x_5_n414), .A3(
        add_x_5_n416), .Y(add_x_5_n398) );
  OR3X1_LVT add_x_5_U333 ( .A1(add_x_5_n395), .A2(add_x_5_n396), .A3(
        add_x_5_n397), .Y(add_x_5_n440) );
  AO222X1_LVT add_x_5_U332 ( .A1(n_T_914[16]), .A2(mem_reg_pc[16]), .A3(
        n_T_914[16]), .A4(add_x_5_n487), .A5(mem_reg_pc[16]), .A6(add_x_5_n487), .Y(add_x_5_n397) );
  OA221X1_LVT add_x_5_U331 ( .A1(add_x_5_n485), .A2(add_x_5_n488), .A3(
        add_x_5_n485), .A4(add_x_5_n486), .A5(add_x_5_n394), .Y(add_x_5_n396)
         );
  AND4X1_LVT add_x_5_U330 ( .A1(add_x_5_n410), .A2(add_x_5_n484), .A3(
        add_x_5_n394), .A4(add_x_5_n488), .Y(add_x_5_n395) );
  OA22X1_LVT add_x_5_U329 ( .A1(n_T_914[15]), .A2(mem_reg_pc[15]), .A3(
        n_T_914[16]), .A4(mem_reg_pc[16]), .Y(add_x_5_n394) );
  FADDX1_LVT add_x_5_U319 ( .A(n_T_914[2]), .B(mem_reg_pc[2]), .CI(
        add_x_5_n408), .CO(add_x_5_n246), .S(mem_br_target_2_) );
endmodule

