
module PlusArgTimeout ( clock, reset, io_count );
  input [31:0] io_count;
  input clock, reset;


endmodule


module RVCExpander ( io_in, io_out_bits, io_out_rd, io_out_rs1, io_out_rs2, 
        io_out_rs3, io_rvc_BAR );
  input [31:0] io_in;
  output [31:0] io_out_bits;
  output [4:0] io_out_rd;
  output [4:0] io_out_rs1;
  output [4:0] io_out_rs2;
  output [4:0] io_out_rs3;
  output io_rvc_BAR;
  wire   n354, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n32,
         n34, n35, n36, n37, n38, n39, n40, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353;

  AO221X1_LVT U3 ( .A1(1'b1), .A2(n223), .A3(n66), .A4(n221), .A5(n32), .Y(
        io_out_bits[17]) );
  AO221X1_LVT U4 ( .A1(1'b1), .A2(n30), .A3(n63), .A4(n265), .A5(n354), .Y(
        io_out_bits[24]) );
  OA221X1_LVT U5 ( .A1(1'b0), .A2(n40), .A3(io_in[13]), .A4(n288), .A5(n169), 
        .Y(n17) );
  OA221X1_LVT U6 ( .A1(1'b0), .A2(n335), .A3(n289), .A4(n161), .A5(n13), .Y(
        n15) );
  NOR2X2_LVT U7 ( .A1(io_in[6]), .A2(n2), .Y(n342) );
  OR2X1_LVT U8 ( .A1(n344), .A2(n203), .Y(n226) );
  AND3X1_LVT U9 ( .A1(n342), .A2(n74), .A3(n290), .Y(n110) );
  AO21X1_LVT U10 ( .A1(n66), .A2(n83), .A3(n223), .Y(io_out_rs1[2]) );
  OA21X1_LVT U11 ( .A1(n70), .A2(n46), .A3(n248), .Y(n141) );
  AND3X1_LVT U12 ( .A1(n46), .A2(n77), .A3(n180), .Y(n205) );
  OAI21X2_LVT U13 ( .A1(n290), .A2(n73), .A3(n234), .Y(io_out_rs2[0]) );
  NAND3X0_LVT U14 ( .A1(n133), .A2(n342), .A3(n152), .Y(n121) );
  NBUFFX2_LVT U15 ( .A(io_in[2]), .Y(n1) );
  NBUFFX2_LVT U16 ( .A(io_in[5]), .Y(n2) );
  AND2X1_LVT U17 ( .A1(n56), .A2(n172), .Y(n3) );
  AND3X2_LVT U18 ( .A1(n154), .A2(n109), .A3(n300), .Y(n163) );
  AO22X2_LVT U19 ( .A1(n320), .A2(n9), .A3(io_rvc_BAR), .A4(io_in[24]), .Y(
        io_out_rs2[4]) );
  AO22X1_LVT U20 ( .A1(n320), .A2(n9), .A3(io_rvc_BAR), .A4(io_in[24]), .Y(
        n354) );
  NBUFFX2_LVT U21 ( .A(io_in[9]), .Y(n5) );
  OR2X4_LVT U22 ( .A1(io_in[10]), .A2(io_in[7]), .Y(n116) );
  AO21X2_LVT U23 ( .A1(n83), .A2(n62), .A3(n204), .Y(io_out_rs1[0]) );
  NAND2X0_LVT U24 ( .A1(n88), .A2(n190), .Y(n6) );
  NAND2X0_LVT U25 ( .A1(n88), .A2(n190), .Y(n7) );
  NAND2X0_LVT U26 ( .A1(n7), .A2(n333), .Y(n279) );
  OR2X4_LVT U27 ( .A1(n179), .A2(n6), .Y(n343) );
  NAND3X2_LVT U28 ( .A1(n154), .A2(n153), .A3(n152), .Y(n8) );
  AND2X4_LVT U29 ( .A1(io_rvc_BAR), .A2(io_in[17]), .Y(n223) );
  NBUFFX2_LVT U30 ( .A(io_in[6]), .Y(n9) );
  NAND3X2_LVT U31 ( .A1(n56), .A2(n48), .A3(n350), .Y(n111) );
  AND3X2_LVT U32 ( .A1(n342), .A2(n300), .A3(n350), .Y(n132) );
  NAND3X2_LVT U33 ( .A1(n203), .A2(n68), .A3(n202), .Y(n221) );
  OA22X2_LVT U34 ( .A1(n71), .A2(n86), .A3(n120), .A4(n203), .Y(n227) );
  AND2X4_LVT U35 ( .A1(n180), .A2(n302), .Y(n91) );
  IBUFFX2_LVT U36 ( .A(n162), .Y(n10) );
  DELLN2X2_LVT U37 ( .A(io_in[6]), .Y(n63) );
  IBUFFX2_LVT U38 ( .A(n320), .Y(n285) );
  AO21X2_LVT U39 ( .A1(n283), .A2(n216), .A3(n279), .Y(n213) );
  NAND2X0_LVT U40 ( .A1(n353), .A2(n352), .Y(io_out_bits[31]) );
  AND2X4_LVT U41 ( .A1(n101), .A2(n93), .Y(n283) );
  NAND3X0_LVT U42 ( .A1(n140), .A2(n329), .A3(n328), .Y(n144) );
  NAND3X2_LVT U43 ( .A1(n10), .A2(n244), .A3(n243), .Y(n254) );
  NAND3X0_LVT U44 ( .A1(n144), .A2(n143), .A3(n142), .Y(io_out_bits[3]) );
  NAND3X2_LVT U45 ( .A1(n330), .A2(n329), .A3(n328), .Y(n331) );
  NOR2X2_LVT U46 ( .A1(io_in[13]), .A2(n57), .Y(n190) );
  OR2X2_LVT U47 ( .A1(io_in[13]), .A2(n57), .Y(n90) );
  IBUFFX2_LVT U48 ( .A(n101), .Y(n78) );
  AO21X1_LVT U49 ( .A1(n70), .A2(n163), .A3(n49), .Y(n127) );
  INVX1_LVT U50 ( .A(io_rvc_BAR), .Y(n71) );
  INVX1_LVT U51 ( .A(n245), .Y(n52) );
  NAND4X0_LVT U52 ( .A1(n155), .A2(n157), .A3(n156), .A4(n260), .Y(
        io_out_bits[5]) );
  INVX1_LVT U53 ( .A(n248), .Y(n35) );
  OA21X1_LVT U54 ( .A1(n270), .A2(n325), .A3(n343), .Y(n271) );
  INVX1_LVT U55 ( .A(n162), .Y(n329) );
  NAND3X0_LVT U56 ( .A1(n185), .A2(n186), .A3(n200), .Y(io_out_bits[12]) );
  INVX1_LVT U57 ( .A(n289), .Y(n62) );
  IBUFFX2_LVT U58 ( .A(io_in[8]), .Y(n300) );
  INVX1_LVT U59 ( .A(io_in[15]), .Y(n89) );
  INVX0_LVT U60 ( .A(n62), .Y(n11) );
  INVX0_LVT U61 ( .A(n164), .Y(n12) );
  NAND3X0_LVT U62 ( .A1(n266), .A2(n1), .A3(n264), .Y(n13) );
  OAI222X1_LVT U64 ( .A1(n11), .A2(n12), .A3(n163), .A4(n232), .A5(n162), .A6(
        n15), .Y(io_out_bits[7]) );
  NAND3X0_LVT U66 ( .A1(n349), .A2(n52), .A3(n264), .Y(n18) );
  NAND3X0_LVT U67 ( .A1(n174), .A2(n216), .A3(n63), .Y(n19) );
  NAND2X0_LVT U68 ( .A1(n66), .A2(n279), .Y(n20) );
  NAND3X0_LVT U69 ( .A1(n20), .A2(n19), .A3(n18), .Y(n21) );
  NAND2X0_LVT U70 ( .A1(n10), .A2(n21), .Y(n22) );
  NAND2X0_LVT U71 ( .A1(n283), .A2(n52), .Y(n23) );
  OR2X1_LVT U72 ( .A1(n168), .A2(n17), .Y(n24) );
  NAND3X0_LVT U73 ( .A1(n24), .A2(n23), .A3(n22), .Y(io_out_bits[9]) );
  NAND4X0_LVT U74 ( .A1(n242), .A2(n210), .A3(n317), .A4(n328), .Y(n25) );
  OA21X1_LVT U75 ( .A1(n178), .A2(n25), .A3(n39), .Y(io_out_bits[11]) );
  AOI22X1_LVT U76 ( .A1(n62), .A2(n221), .A3(n64), .A4(n38), .Y(n26) );
  INVX0_LVT U77 ( .A(n204), .Y(n27) );
  NAND3X0_LVT U78 ( .A1(n222), .A2(n26), .A3(n27), .Y(io_out_bits[15]) );
  AND4X1_LVT U79 ( .A1(n224), .A2(n328), .A3(n225), .A4(n235), .Y(n28) );
  NAND2X0_LVT U80 ( .A1(n226), .A2(n28), .Y(io_out_bits[18]) );
  NAND2X0_LVT U81 ( .A1(n67), .A2(n242), .Y(n29) );
  AND2X4_LVT U82 ( .A1(n300), .A2(n29), .Y(n212) );
  OA221X1_LVT U83 ( .A1(n263), .A2(n264), .A3(n263), .A4(n39), .A5(n336), .Y(
        n30) );
  INVX0_LVT U85 ( .A(n235), .Y(n32) );
  INVX1_LVT U87 ( .A(n151), .Y(n38) );
  OR3X2_LVT U88 ( .A1(n146), .A2(n171), .A3(n145), .Y(n150) );
  NAND2X2_LVT U89 ( .A1(n274), .A2(n273), .Y(io_out_bits[25]) );
  OR2X4_LVT U90 ( .A1(n343), .A2(n344), .Y(n345) );
  NAND3X1_LVT U91 ( .A1(n277), .A2(n317), .A3(n343), .Y(n265) );
  AND2X1_LVT U92 ( .A1(n101), .A2(io_in[15]), .Y(n34) );
  NAND3X2_LVT U93 ( .A1(n318), .A2(n317), .A3(n334), .Y(n319) );
  AND2X4_LVT U94 ( .A1(n334), .A2(n317), .Y(n276) );
  OA21X2_LVT U95 ( .A1(n53), .A2(n301), .A3(n334), .Y(n194) );
  AND4X2_LVT U96 ( .A1(io_in[13]), .A2(n120), .A3(n168), .A4(n344), .Y(n114)
         );
  IBUFFX2_LVT U97 ( .A(n120), .Y(n39) );
  OR2X2_LVT U98 ( .A1(n172), .A2(n171), .Y(n309) );
  AOI21X1_LVT U99 ( .A1(n35), .A2(n163), .A3(n36), .Y(n119) );
  AND4X2_LVT U100 ( .A1(n115), .A2(n114), .A3(n300), .A4(n289), .Y(n36) );
  AND2X4_LVT U101 ( .A1(n168), .A2(n120), .Y(n153) );
  AO22X2_LVT U102 ( .A1(n241), .A2(n52), .A3(n100), .A4(n66), .Y(io_out_rd[2])
         );
  NAND3X2_LVT U103 ( .A1(n101), .A2(io_in[15]), .A3(io_in[13]), .Y(n102) );
  OR3X2_LVT U104 ( .A1(n101), .A2(n290), .A3(n162), .Y(n98) );
  AND3X4_LVT U105 ( .A1(n229), .A2(n228), .A3(n242), .Y(n250) );
  OR2X2_LVT U106 ( .A1(n188), .A2(n229), .Y(n334) );
  NAND2X0_LVT U107 ( .A1(n332), .A2(n331), .Y(io_out_bits[28]) );
  NAND2X0_LVT U108 ( .A1(n92), .A2(n320), .Y(n37) );
  IBUFFX2_LVT U109 ( .A(io_in[11]), .Y(n120) );
  NAND3X2_LVT U110 ( .A1(n90), .A2(n320), .A3(n70), .Y(n268) );
  IBUFFX2_LVT U111 ( .A(n163), .Y(n233) );
  IBUFFX2_LVT U112 ( .A(n2), .Y(n151) );
  NAND3X2_LVT U113 ( .A1(n270), .A2(n9), .A3(n38), .Y(n183) );
  NAND3X1_LVT U114 ( .A1(n320), .A2(io_in[15]), .A3(n190), .Y(n61) );
  AND3X4_LVT U115 ( .A1(n320), .A2(io_in[15]), .A3(n190), .Y(n172) );
  NAND3X2_LVT U116 ( .A1(n112), .A2(n113), .A3(n90), .Y(n302) );
  NOR2X4_LVT U117 ( .A1(io_in[1]), .A2(n60), .Y(n241) );
  NAND3X2_LVT U118 ( .A1(n75), .A2(n60), .A3(n89), .Y(n333) );
  AND3X2_LVT U119 ( .A1(n75), .A2(n60), .A3(n89), .Y(n47) );
  OR2X2_LVT U120 ( .A1(n97), .A2(n51), .Y(n162) );
  NAND2X1_LVT U121 ( .A1(n227), .A2(n87), .Y(io_out_rs1[4]) );
  INVX1_LVT U122 ( .A(n211), .Y(n115) );
  OR2X1_LVT U123 ( .A1(n117), .A2(n333), .Y(n210) );
  NOR2X1_LVT U124 ( .A1(n117), .A2(n333), .Y(n48) );
  INVX0_LVT U125 ( .A(io_in[1]), .Y(n75) );
  IBUFFX2_LVT U126 ( .A(io_rvc_BAR), .Y(n40) );
  INVX0_LVT U127 ( .A(io_in[10]), .Y(n344) );
  INVX1_LVT U128 ( .A(io_in[12]), .Y(n350) );
  NAND3X0_LVT U129 ( .A1(n99), .A2(n232), .A3(n98), .Y(io_out_rd[0]) );
  AO22X1_LVT U130 ( .A1(n107), .A2(n106), .A3(io_in[10]), .A4(n105), .Y(
        io_out_rd[3]) );
  NAND3X1_LVT U131 ( .A1(n194), .A2(n193), .A3(n192), .Y(io_out_bits[13]) );
  INVX0_LVT U132 ( .A(n104), .Y(n107) );
  NOR2X1_LVT U133 ( .A1(n280), .A2(n279), .Y(n337) );
  INVX0_LVT U134 ( .A(n279), .Y(n161) );
  NOR2X1_LVT U135 ( .A1(n174), .A2(n279), .Y(n264) );
  OR2X1_LVT U136 ( .A1(n261), .A2(n336), .Y(io_out_rs2[3]) );
  INVX0_LVT U137 ( .A(n317), .Y(n257) );
  INVX1_LVT U138 ( .A(n277), .Y(n325) );
  NOR2X1_LVT U139 ( .A1(io_rvc_BAR), .A2(n291), .Y(n96) );
  AND2X1_LVT U140 ( .A1(n190), .A2(n34), .Y(n270) );
  OR2X1_LVT U141 ( .A1(n61), .A2(n110), .Y(n170) );
  AND2X1_LVT U142 ( .A1(n211), .A2(n177), .Y(n317) );
  OR2X1_LVT U143 ( .A1(n350), .A2(n53), .Y(n275) );
  OAI21X1_LVT U144 ( .A1(n301), .A2(n73), .A3(n237), .Y(io_out_rs2[1]) );
  NOR2X1_LVT U145 ( .A1(n5), .A2(n39), .Y(n109) );
  NOR2X1_LVT U146 ( .A1(n89), .A2(n71), .Y(n204) );
  OR2X1_LVT U147 ( .A1(n1), .A2(n40), .Y(n129) );
  OR2X1_LVT U148 ( .A1(n72), .A2(n40), .Y(n237) );
  OAI21X1_LVT U149 ( .A1(n245), .A2(n73), .A3(n246), .Y(io_out_rs2[2]) );
  INVX1_LVT U150 ( .A(n241), .Y(n182) );
  NAND3X0_LVT U151 ( .A1(io_in[8]), .A2(n216), .A3(io_in[15]), .Y(n217) );
  INVX0_LVT U152 ( .A(n342), .Y(n196) );
  INVX0_LVT U153 ( .A(n63), .Y(n298) );
  NOR2X1_LVT U154 ( .A1(io_in[4]), .A2(n55), .Y(n74) );
  INVX0_LVT U155 ( .A(io_in[27]), .Y(n303) );
  INVX1_LVT U156 ( .A(io_in[21]), .Y(n72) );
  NAND3X0_LVT U157 ( .A1(n121), .A2(n216), .A3(n242), .Y(n122) );
  AND2X4_LVT U158 ( .A1(n60), .A2(io_in[1]), .Y(io_rvc_BAR) );
  NAND2X0_LVT U159 ( .A1(n56), .A2(n172), .Y(n46) );
  OR2X1_LVT U160 ( .A1(io_in[13]), .A2(n333), .Y(n177) );
  AND2X1_LVT U161 ( .A1(n92), .A2(n101), .Y(n340) );
  NOR3X0_LVT U162 ( .A1(n89), .A2(n216), .A3(n57), .Y(n92) );
  NAND2X0_LVT U163 ( .A1(n110), .A2(n172), .Y(n49) );
  NAND2X0_LVT U164 ( .A1(n110), .A2(n172), .Y(n50) );
  NAND4X0_LVT U165 ( .A1(n82), .A2(n207), .A3(n81), .A4(n80), .Y(io_out_rs1[1]) );
  IBUFFX2_LVT U166 ( .A(io_in[2]), .Y(n290) );
  NAND2X0_LVT U167 ( .A1(n288), .A2(n96), .Y(n51) );
  OA22X1_LVT U168 ( .A1(n290), .A2(n302), .A3(n289), .A4(n288), .Y(n294) );
  INVX1_LVT U169 ( .A(n168), .Y(n66) );
  NAND3X0_LVT U170 ( .A1(n209), .A2(n47), .A3(n118), .Y(n53) );
  NAND3X0_LVT U171 ( .A1(n209), .A2(n47), .A3(n118), .Y(n54) );
  OR3X2_LVT U172 ( .A1(n5), .A2(io_in[11]), .A3(n116), .Y(n209) );
  NAND3X0_LVT U173 ( .A1(n209), .A2(n47), .A3(n118), .Y(n316) );
  NOR2X2_LVT U174 ( .A1(n283), .A2(n340), .Y(n349) );
  NAND3X0_LVT U175 ( .A1(n160), .A2(n349), .A3(n159), .Y(io_out_bits[6]) );
  NBUFFX2_LVT U176 ( .A(io_in[3]), .Y(n55) );
  AND3X1_LVT U177 ( .A1(n342), .A2(n74), .A3(n290), .Y(n56) );
  NBUFFX2_LVT U178 ( .A(io_in[14]), .Y(n57) );
  OR2X1_LVT U179 ( .A1(n58), .A2(n90), .Y(n59) );
  NAND2X0_LVT U180 ( .A1(n320), .A2(n89), .Y(n58) );
  NBUFFX2_LVT U181 ( .A(io_in[0]), .Y(n60) );
  OA21X2_LVT U182 ( .A1(io_in[1]), .A2(n93), .A3(n60), .Y(n73) );
  AND3X1_LVT U183 ( .A1(n209), .A2(n47), .A3(n118), .Y(n64) );
  NAND4X0_LVT U184 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .Y(
        io_out_bits[14]) );
  NAND2X0_LVT U185 ( .A1(n92), .A2(n101), .Y(n65) );
  OA21X1_LVT U186 ( .A1(n172), .A2(n340), .A3(n170), .Y(n176) );
  OR2X1_LVT U187 ( .A1(n340), .A2(n215), .Y(n218) );
  NAND2X0_LVT U188 ( .A1(n288), .A2(n96), .Y(n171) );
  NAND3X0_LVT U189 ( .A1(n154), .A2(n153), .A3(n152), .Y(n158) );
  IBUFFX2_LVT U190 ( .A(n60), .Y(n113) );
  INVX1_LVT U191 ( .A(n270), .Y(n201) );
  OA21X1_LVT U192 ( .A1(n216), .A2(n184), .A3(n183), .Y(n185) );
  AND2X1_LVT U193 ( .A1(n75), .A2(n60), .Y(n101) );
  NAND3X0_LVT U194 ( .A1(n67), .A2(n38), .A3(n333), .Y(n255) );
  NAND2X0_LVT U195 ( .A1(n241), .A2(n90), .Y(n67) );
  AND2X1_LVT U196 ( .A1(n256), .A2(n242), .Y(n68) );
  NAND4X1_LVT U197 ( .A1(n329), .A2(n55), .A3(n264), .A4(n65), .Y(n165) );
  AND2X1_LVT U198 ( .A1(n101), .A2(io_in[15]), .Y(n88) );
  NAND4X0_LVT U199 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(
        io_out_bits[30]) );
  INVX1_LVT U200 ( .A(io_in[4]), .Y(n245) );
  NAND3X1_LVT U201 ( .A1(n321), .A2(io_in[13]), .A3(n320), .Y(n323) );
  IBUFFX2_LVT U202 ( .A(io_in[13]), .Y(n216) );
  OR2X2_LVT U203 ( .A1(n283), .A2(n340), .Y(n296) );
  AOI22X1_LVT U204 ( .A1(io_rvc_BAR), .A2(io_in[30]), .A3(n340), .A4(io_in[8]), 
        .Y(n347) );
  AO22X1_LVT U205 ( .A1(n241), .A2(n55), .A3(n100), .A4(io_in[8]), .Y(
        io_out_rd[1]) );
  AND3X1_LVT U206 ( .A1(n286), .A2(n333), .A3(n59), .Y(n106) );
  NAND3X0_LVT U207 ( .A1(n328), .A2(n228), .A3(n40), .Y(n206) );
  NAND3X0_LVT U208 ( .A1(n348), .A2(n339), .A3(n338), .Y(io_out_bits[29]) );
  NOR2X0_LVT U209 ( .A1(io_in[1]), .A2(n283), .Y(n336) );
  OR2X1_LVT U210 ( .A1(n350), .A2(n49), .Y(n232) );
  AND2X1_LVT U211 ( .A1(n315), .A2(n314), .Y(io_out_bits[27]) );
  INVX1_LVT U212 ( .A(n55), .Y(n301) );
  INVX1_LVT U213 ( .A(n296), .Y(n266) );
  AND3X2_LVT U214 ( .A1(n130), .A2(n129), .A3(n128), .Y(io_out_bits[2]) );
  OR2X1_LVT U215 ( .A1(n195), .A2(n173), .Y(n248) );
  INVX1_LVT U216 ( .A(n350), .Y(n70) );
  NAND3X2_LVT U217 ( .A1(n226), .A2(n225), .A3(n85), .Y(io_out_rs1[3]) );
  INVX1_LVT U218 ( .A(n283), .Y(n328) );
  INVX1_LVT U219 ( .A(n242), .Y(n174) );
  OA21X2_LVT U220 ( .A1(n47), .A2(n178), .A3(n39), .Y(io_out_rd[4]) );
  OR2X2_LVT U221 ( .A1(n210), .A2(n209), .Y(n277) );
  AND2X1_LVT U222 ( .A1(n57), .A2(io_in[15]), .Y(n93) );
  OR2X2_LVT U223 ( .A1(n89), .A2(n182), .Y(n242) );
  OR2X2_LVT U224 ( .A1(n57), .A2(n333), .Y(n211) );
  AND2X2_LVT U225 ( .A1(n113), .A2(io_in[1]), .Y(n320) );
  NAND3X0_LVT U226 ( .A1(n203), .A2(n68), .A3(n244), .Y(n83) );
  AND4X1_LVT U227 ( .A1(n317), .A2(n63), .A3(n242), .A4(n297), .Y(n243) );
  AND2X1_LVT U228 ( .A1(n96), .A2(n288), .Y(n94) );
  OA21X1_LVT U229 ( .A1(n350), .A2(n71), .A3(n59), .Y(n181) );
  AND2X1_LVT U230 ( .A1(n153), .A2(n154), .Y(n133) );
  NAND2X0_LVT U231 ( .A1(io_rvc_BAR), .A2(io_in[20]), .Y(n234) );
  NAND2X0_LVT U232 ( .A1(io_rvc_BAR), .A2(io_in[22]), .Y(n246) );
  AO22X1_LVT U233 ( .A1(n320), .A2(n38), .A3(io_rvc_BAR), .A4(io_in[23]), .Y(
        n261) );
  AND2X1_LVT U234 ( .A1(n320), .A2(n190), .Y(n126) );
  NAND2X0_LVT U235 ( .A1(n126), .A2(n89), .Y(n180) );
  AND2X1_LVT U236 ( .A1(n180), .A2(n211), .Y(n76) );
  NAND2X0_LVT U237 ( .A1(io_in[12]), .A2(n172), .Y(n77) );
  AND3X1_LVT U238 ( .A1(n50), .A2(n76), .A3(n77), .Y(n203) );
  NAND2X0_LVT U239 ( .A1(n241), .A2(n90), .Y(n256) );
  NAND2X0_LVT U240 ( .A1(n67), .A2(n242), .Y(n280) );
  NAND2X0_LVT U241 ( .A1(n57), .A2(io_in[13]), .Y(n117) );
  NOR3X0_LVT U242 ( .A1(n48), .A2(n270), .A3(n296), .Y(n244) );
  AO21X1_LVT U243 ( .A1(n244), .A2(n211), .A3(n300), .Y(n82) );
  NAND2X0_LVT U244 ( .A1(io_rvc_BAR), .A2(io_in[16]), .Y(n207) );
  OR2X1_LVT U245 ( .A1(n300), .A2(n205), .Y(n81) );
  INVX1_LVT U246 ( .A(n212), .Y(n79) );
  INVX1_LVT U247 ( .A(n126), .Y(n228) );
  NAND4X0_LVT U248 ( .A1(n79), .A2(n78), .A3(n228), .A4(n40), .Y(n80) );
  AND2X1_LVT U249 ( .A1(n201), .A2(n68), .Y(n225) );
  NAND2X0_LVT U250 ( .A1(io_in[10]), .A2(n48), .Y(n84) );
  NAND2X0_LVT U251 ( .A1(io_rvc_BAR), .A2(io_in[18]), .Y(n224) );
  AND3X1_LVT U252 ( .A1(n349), .A2(n84), .A3(n224), .Y(n85) );
  INVX1_LVT U253 ( .A(io_in[19]), .Y(n86) );
  OR2X1_LVT U254 ( .A1(n120), .A2(n210), .Y(n87) );
  NAND2X0_LVT U255 ( .A1(n88), .A2(n190), .Y(n229) );
  INVX1_LVT U256 ( .A(n213), .Y(n95) );
  AND2X1_LVT U257 ( .A1(io_in[1]), .A2(n89), .Y(n112) );
  AND2X1_LVT U258 ( .A1(n91), .A2(n170), .Y(n169) );
  AND2X1_LVT U259 ( .A1(n92), .A2(n320), .Y(n291) );
  NAND2X0_LVT U260 ( .A1(n93), .A2(n320), .Y(n288) );
  AND2X1_LVT U261 ( .A1(n169), .A2(n94), .Y(n108) );
  NAND2X0_LVT U262 ( .A1(n95), .A2(n108), .Y(n100) );
  NAND2X0_LVT U263 ( .A1(n62), .A2(n100), .Y(n99) );
  NAND2X0_LVT U264 ( .A1(n302), .A2(n228), .Y(n97) );
  AND2X1_LVT U265 ( .A1(n37), .A2(n302), .Y(n103) );
  NAND3X0_LVT U266 ( .A1(n103), .A2(n61), .A3(n102), .Y(n104) );
  AND2X1_LVT U267 ( .A1(n288), .A2(n40), .Y(n286) );
  NAND3X0_LVT U268 ( .A1(n104), .A2(n103), .A3(n170), .Y(n105) );
  INVX1_LVT U269 ( .A(n108), .Y(n178) );
  AND2X1_LVT U270 ( .A1(n111), .A2(n65), .Y(n138) );
  AND2X1_LVT U271 ( .A1(n127), .A2(n138), .Y(n125) );
  INVX1_LVT U272 ( .A(n57), .Y(n195) );
  NAND2X0_LVT U273 ( .A1(n113), .A2(n112), .Y(n173) );
  INVX1_LVT U274 ( .A(io_in[7]), .Y(n289) );
  INVX1_LVT U275 ( .A(n117), .Y(n118) );
  AND3X1_LVT U276 ( .A1(n119), .A2(n71), .A3(n54), .Y(n124) );
  INVX1_LVT U277 ( .A(n5), .Y(n168) );
  NOR2X0_LVT U278 ( .A1(io_in[10]), .A2(n62), .Y(n154) );
  AND2X1_LVT U279 ( .A1(n300), .A2(n350), .Y(n152) );
  NAND3X0_LVT U280 ( .A1(n122), .A2(n161), .A3(n195), .Y(n123) );
  NAND3X0_LVT U281 ( .A1(n125), .A2(n124), .A3(n123), .Y(n130) );
  NAND2X0_LVT U282 ( .A1(n127), .A2(n126), .Y(n128) );
  NAND2X0_LVT U283 ( .A1(io_in[11]), .A2(io_in[10]), .Y(n187) );
  INVX1_LVT U284 ( .A(n187), .Y(n179) );
  AND2X1_LVT U285 ( .A1(n270), .A2(n179), .Y(n341) );
  NAND2X0_LVT U286 ( .A1(n341), .A2(n70), .Y(n131) );
  OA21X1_LVT U287 ( .A1(n211), .A2(n216), .A3(n131), .Y(n139) );
  NAND2X0_LVT U288 ( .A1(n190), .A2(io_in[15]), .Y(n136) );
  NAND3X0_LVT U289 ( .A1(n133), .A2(n132), .A3(n256), .Y(n135) );
  NAND3X0_LVT U290 ( .A1(n201), .A2(n210), .A3(n177), .Y(n134) );
  AO21X1_LVT U291 ( .A1(n135), .A2(n136), .A3(n134), .Y(n137) );
  NAND3X0_LVT U292 ( .A1(n139), .A2(n138), .A3(n137), .Y(n140) );
  OR2X1_LVT U293 ( .A1(n233), .A2(n141), .Y(n143) );
  NAND2X0_LVT U294 ( .A1(io_rvc_BAR), .A2(n55), .Y(n142) );
  NAND2X0_LVT U295 ( .A1(n302), .A2(n67), .Y(n146) );
  NAND2X0_LVT U296 ( .A1(n61), .A2(n349), .Y(n145) );
  OA21X1_LVT U297 ( .A1(n40), .A2(n245), .A3(n170), .Y(n149) );
  NAND2X0_LVT U298 ( .A1(n61), .A2(n248), .Y(n147) );
  NAND2X0_LVT U299 ( .A1(n163), .A2(n147), .Y(n148) );
  NAND3X0_LVT U300 ( .A1(n150), .A2(n149), .A3(n148), .Y(io_out_bits[4]) );
  NOR2X0_LVT U301 ( .A1(n174), .A2(n341), .Y(n260) );
  AND3X1_LVT U302 ( .A1(n170), .A2(n266), .A3(n54), .Y(n157) );
  AND2X1_LVT U303 ( .A1(n37), .A2(n288), .Y(n299) );
  OA21X1_LVT U304 ( .A1(n71), .A2(n151), .A3(n299), .Y(n156) );
  NAND2X0_LVT U305 ( .A1(n8), .A2(n172), .Y(n155) );
  NAND2X0_LVT U306 ( .A1(n158), .A2(n3), .Y(n160) );
  NAND2X0_LVT U307 ( .A1(n63), .A2(io_rvc_BAR), .Y(n159) );
  NAND2X0_LVT U308 ( .A1(n283), .A2(n70), .Y(n335) );
  NAND2X0_LVT U309 ( .A1(n169), .A2(n40), .Y(n164) );
  NAND2X0_LVT U310 ( .A1(n164), .A2(io_in[8]), .Y(n167) );
  NAND2X0_LVT U311 ( .A1(n279), .A2(io_in[8]), .Y(n166) );
  NAND3X0_LVT U312 ( .A1(n167), .A2(n166), .A3(n165), .Y(io_out_bits[8]) );
  NAND2X0_LVT U313 ( .A1(n349), .A2(n173), .Y(n310) );
  OR3X1_LVT U314 ( .A1(n174), .A2(n47), .A3(n310), .Y(n175) );
  OAI22X1_LVT U315 ( .A1(n176), .A2(n344), .A3(n309), .A4(n175), .Y(
        io_out_bits[10]) );
  NAND2X0_LVT U316 ( .A1(n340), .A2(n70), .Y(n222) );
  AND2X1_LVT U317 ( .A1(n222), .A2(n343), .Y(n200) );
  OA21X1_LVT U318 ( .A1(n316), .A2(n290), .A3(n181), .Y(n186) );
  AND3X1_LVT U319 ( .A1(n328), .A2(n285), .A3(n182), .Y(n184) );
  NAND2X0_LVT U320 ( .A1(io_in[11]), .A2(n187), .Y(n188) );
  OR2X1_LVT U321 ( .A1(n216), .A2(n40), .Y(n189) );
  OA21X1_LVT U322 ( .A1(n190), .A2(n285), .A3(n189), .Y(n191) );
  AND3X1_LVT U323 ( .A1(n68), .A2(n191), .A3(n222), .Y(n193) );
  NAND2X0_LVT U324 ( .A1(n63), .A2(n341), .Y(n192) );
  OR2X1_LVT U325 ( .A1(n195), .A2(n40), .Y(n199) );
  NAND2X0_LVT U326 ( .A1(n52), .A2(n64), .Y(n198) );
  NAND3X0_LVT U327 ( .A1(n270), .A2(n196), .A3(n350), .Y(n197) );
  AND2X1_LVT U328 ( .A1(n201), .A2(n328), .Y(n202) );
  AO21X1_LVT U329 ( .A1(n205), .A2(n328), .A3(n300), .Y(n208) );
  NAND3X0_LVT U330 ( .A1(n208), .A2(n207), .A3(n206), .Y(n220) );
  AND2X1_LVT U331 ( .A1(n211), .A2(n277), .Y(n214) );
  OA222X1_LVT U332 ( .A1(n298), .A2(n53), .A3(n300), .A4(n214), .A5(n213), 
        .A6(n212), .Y(n215) );
  NAND3X0_LVT U333 ( .A1(n218), .A2(n222), .A3(n217), .Y(n219) );
  AND2X1_LVT U334 ( .A1(n220), .A2(n219), .Y(io_out_bits[16]) );
  AND2X1_LVT U335 ( .A1(n275), .A2(n222), .Y(n235) );
  NAND2X0_LVT U336 ( .A1(n227), .A2(n235), .Y(io_out_bits[19]) );
  NAND3X0_LVT U337 ( .A1(n250), .A2(n317), .A3(n299), .Y(n230) );
  NAND2X0_LVT U338 ( .A1(n1), .A2(n230), .Y(n231) );
  OA21X1_LVT U339 ( .A1(n233), .A2(n232), .A3(n231), .Y(n236) );
  NAND3X0_LVT U340 ( .A1(n236), .A2(n235), .A3(n234), .Y(io_out_bits[20]) );
  NAND2X0_LVT U341 ( .A1(n237), .A2(n301), .Y(n240) );
  INVX1_LVT U342 ( .A(n275), .Y(n263) );
  NAND4X0_LVT U343 ( .A1(n299), .A2(n317), .A3(n65), .A4(n237), .Y(n239) );
  NAND2X0_LVT U344 ( .A1(n275), .A2(n250), .Y(n238) );
  OA22X1_LVT U345 ( .A1(n240), .A2(n263), .A3(n239), .A4(n238), .Y(
        io_out_bits[21]) );
  NAND2X0_LVT U346 ( .A1(io_in[13]), .A2(n241), .Y(n297) );
  OR2X1_LVT U347 ( .A1(n245), .A2(n299), .Y(n247) );
  AND3X1_LVT U348 ( .A1(n247), .A2(n275), .A3(n246), .Y(n253) );
  OA21X1_LVT U349 ( .A1(io_in[13]), .A2(n248), .A3(n65), .Y(n249) );
  NAND3X0_LVT U350 ( .A1(n250), .A2(n317), .A3(n249), .Y(n251) );
  NAND2X0_LVT U351 ( .A1(n52), .A2(n251), .Y(n252) );
  NAND3X0_LVT U352 ( .A1(n254), .A2(n253), .A3(n252), .Y(io_out_bits[22]) );
  OA21X1_LVT U353 ( .A1(n344), .A2(n256), .A3(n255), .Y(n259) );
  NAND2X0_LVT U354 ( .A1(n257), .A2(n38), .Y(n258) );
  NAND4X0_LVT U355 ( .A1(n260), .A2(n259), .A3(n275), .A4(n258), .Y(n262) );
  AO21X1_LVT U356 ( .A1(n262), .A2(n336), .A3(n261), .Y(io_out_bits[23]) );
  AO21X1_LVT U357 ( .A1(n266), .A2(n277), .A3(n290), .Y(n269) );
  NAND2X0_LVT U358 ( .A1(io_in[25]), .A2(io_rvc_BAR), .Y(n267) );
  AND3X1_LVT U359 ( .A1(n269), .A2(n268), .A3(n267), .Y(n274) );
  OR2X1_LVT U360 ( .A1(n350), .A2(n296), .Y(n272) );
  OR3X1_LVT U361 ( .A1(n272), .A2(n271), .A3(n309), .Y(n273) );
  OA21X1_LVT U362 ( .A1(n350), .A2(n276), .A3(n275), .Y(n307) );
  NAND3X0_LVT U363 ( .A1(n277), .A2(n68), .A3(n328), .Y(n278) );
  NAND2X0_LVT U364 ( .A1(n38), .A2(n278), .Y(n282) );
  NAND2X0_LVT U365 ( .A1(n62), .A2(n337), .Y(n281) );
  NAND3X0_LVT U366 ( .A1(n307), .A2(n282), .A3(n281), .Y(n287) );
  NAND2X0_LVT U367 ( .A1(n283), .A2(n282), .Y(n284) );
  NAND4X0_LVT U368 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .Y(n295) );
  NAND2X0_LVT U369 ( .A1(n62), .A2(n291), .Y(n293) );
  NAND2X0_LVT U370 ( .A1(io_in[26]), .A2(io_rvc_BAR), .Y(n292) );
  NAND4X0_LVT U371 ( .A1(n295), .A2(n294), .A3(n293), .A4(n292), .Y(
        io_out_bits[26]) );
  NAND2X0_LVT U372 ( .A1(n296), .A2(n9), .Y(n311) );
  OA21X1_LVT U373 ( .A1(n298), .A2(n297), .A3(n311), .Y(n305) );
  OA222X1_LVT U374 ( .A1(n40), .A2(n303), .A3(n302), .A4(n301), .A5(n300), 
        .A6(n299), .Y(n312) );
  NAND2X0_LVT U375 ( .A1(n325), .A2(n55), .Y(n304) );
  AND3X1_LVT U376 ( .A1(n305), .A2(n312), .A3(n304), .Y(n308) );
  NAND2X0_LVT U377 ( .A1(n337), .A2(io_in[8]), .Y(n306) );
  NAND3X0_LVT U378 ( .A1(n308), .A2(n307), .A3(n306), .Y(n315) );
  AO21X1_LVT U379 ( .A1(n311), .A2(n310), .A3(n309), .Y(n313) );
  NAND2X0_LVT U380 ( .A1(n313), .A2(n312), .Y(n314) );
  AND2X1_LVT U381 ( .A1(n54), .A2(n328), .Y(n318) );
  NAND2X0_LVT U382 ( .A1(n70), .A2(n319), .Y(n324) );
  MUX21X1_LVT U383 ( .A1(n52), .A2(n66), .S0(io_in[15]), .Y(n321) );
  NAND2X0_LVT U384 ( .A1(io_in[28]), .A2(io_rvc_BAR), .Y(n322) );
  AND3X1_LVT U385 ( .A1(n324), .A2(n323), .A3(n322), .Y(n332) );
  NAND2X0_LVT U386 ( .A1(n52), .A2(n325), .Y(n327) );
  NAND2X0_LVT U387 ( .A1(n66), .A2(n337), .Y(n326) );
  NAND2X0_LVT U388 ( .A1(n327), .A2(n326), .Y(n330) );
  AO21X1_LVT U389 ( .A1(n333), .A2(n334), .A3(n350), .Y(n353) );
  AND2X1_LVT U390 ( .A1(n353), .A2(n335), .Y(n348) );
  NAND2X0_LVT U391 ( .A1(io_in[29]), .A2(io_rvc_BAR), .Y(n339) );
  NAND3X0_LVT U392 ( .A1(n337), .A2(io_in[10]), .A3(n336), .Y(n338) );
  NAND2X0_LVT U393 ( .A1(n342), .A2(n341), .Y(n346) );
  INVX1_LVT U394 ( .A(io_in[31]), .Y(n351) );
  OA22X1_LVT U395 ( .A1(n40), .A2(n351), .A3(n350), .A4(n349), .Y(n352) );
endmodule


module SNPS_CLOCK_GATE_HIGH_IBuf ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module IBuf ( clock, reset, io_imem_ready, io_imem_valid, 
        io_imem_bits_btb_taken, io_imem_bits_btb_bridx, io_imem_bits_btb_entry, 
        io_imem_bits_btb_bht_history, io_imem_bits_pc, io_imem_bits_data, 
        io_imem_bits_xcpt_pf_inst, io_imem_bits_xcpt_ae_inst, 
        io_imem_bits_replay, io_kill, io_pc, io_btb_resp_entry, 
        io_btb_resp_bht_history, io_inst_0_ready, io_inst_0_valid, 
        io_inst_0_bits_xcpt0_pf_inst, io_inst_0_bits_xcpt0_ae_inst, 
        io_inst_0_bits_xcpt1_pf_inst, io_inst_0_bits_xcpt1_ae_inst, 
        io_inst_0_bits_replay, io_inst_0_bits_inst_bits, 
        io_inst_0_bits_inst_rd, io_inst_0_bits_inst_rs1, 
        io_inst_0_bits_inst_rs2, io_inst_0_bits_inst_rs3, io_inst_0_bits_raw, 
        io_inst_0_bits_rvc );
  input [4:0] io_imem_bits_btb_entry;
  input [7:0] io_imem_bits_btb_bht_history;
  input [39:0] io_imem_bits_pc;
  input [31:0] io_imem_bits_data;
  output [39:0] io_pc;
  output [4:0] io_btb_resp_entry;
  output [7:0] io_btb_resp_bht_history;
  output [31:0] io_inst_0_bits_inst_bits;
  output [4:0] io_inst_0_bits_inst_rd;
  output [4:0] io_inst_0_bits_inst_rs1;
  output [4:0] io_inst_0_bits_inst_rs2;
  output [4:0] io_inst_0_bits_inst_rs3;
  output [31:0] io_inst_0_bits_raw;
  input clock, reset, io_imem_valid, io_imem_bits_btb_taken,
         io_imem_bits_btb_bridx, io_imem_bits_xcpt_pf_inst,
         io_imem_bits_xcpt_ae_inst, io_imem_bits_replay, io_kill,
         io_inst_0_ready;
  output io_imem_ready, io_inst_0_valid, io_inst_0_bits_xcpt0_pf_inst,
         io_inst_0_bits_xcpt0_ae_inst, io_inst_0_bits_xcpt1_pf_inst,
         io_inst_0_bits_xcpt1_ae_inst, io_inst_0_bits_replay,
         io_inst_0_bits_rvc;
  wire   n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         buf__replay, n_T_27_0_, n_T_55_91_, n_T_55_85_, n_T_55_84_,
         buf__xcpt_pf_inst, buf__xcpt_ae_inst, N51, net35341, n12, n40, n5, n7,
         n8, n9, n10, n11, n18, n19, n20, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         io_inst_0_bits_inst_rs3_4, io_inst_0_bits_inst_rs3_2,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7;
  wire   [15:0] n_T_34;
  wire   [15:0] buf__data;
  wire   [39:0] buf__pc;
  wire   [4:0] ibufBTBResp_entry;
  wire   [7:0] ibufBTBResp_bht_history;

  RVCExpander RVCExpander ( .io_in({io_inst_0_bits_raw[31:28], n_T_55_91_, 
        io_inst_0_bits_raw[26:22], n_T_55_85_, n_T_55_84_, 
        io_inst_0_bits_raw[19:16], n123, n124, n125, n126, 
        io_inst_0_bits_raw[11], n127, io_inst_0_bits_raw[9:7], n128, 
        io_inst_0_bits_raw[5:4], n129, io_inst_0_bits_raw[2], n130, n131}), 
        .io_out_bits({io_inst_0_bits_inst_bits[31:2], SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .io_out_rd(io_inst_0_bits_inst_rd), 
        .io_out_rs1(io_inst_0_bits_inst_rs1), .io_out_rs2(
        io_inst_0_bits_inst_rs2), .io_out_rs3({SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7}), .io_rvc_BAR(n122) );
  SNPS_CLOCK_GATE_HIGH_IBuf clk_gate_ibufBTBResp_bht_history_reg ( .CLK(clock), 
        .EN(N51), .ENCLK(net35341), .TE(1'b0) );
  DFFX1_LVT buf__data_reg_0_ ( .D(n_T_34[0]), .CLK(n43), .Q(buf__data[0]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_7_ ( .D(
        io_imem_bits_btb_bht_history[7]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[7]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_6_ ( .D(
        io_imem_bits_btb_bht_history[6]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[6]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_5_ ( .D(
        io_imem_bits_btb_bht_history[5]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[5]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_4_ ( .D(
        io_imem_bits_btb_bht_history[4]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[4]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_3_ ( .D(
        io_imem_bits_btb_bht_history[3]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[3]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_2_ ( .D(
        io_imem_bits_btb_bht_history[2]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[2]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_1_ ( .D(
        io_imem_bits_btb_bht_history[1]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[1]) );
  DFFX1_LVT ibufBTBResp_bht_history_reg_0_ ( .D(
        io_imem_bits_btb_bht_history[0]), .CLK(n43), .Q(
        ibufBTBResp_bht_history[0]) );
  DFFX1_LVT ibufBTBResp_entry_reg_4_ ( .D(io_imem_bits_btb_entry[4]), .CLK(n43), .Q(ibufBTBResp_entry[4]) );
  DFFX1_LVT ibufBTBResp_entry_reg_3_ ( .D(io_imem_bits_btb_entry[3]), .CLK(n43), .Q(ibufBTBResp_entry[3]) );
  DFFX1_LVT ibufBTBResp_entry_reg_2_ ( .D(io_imem_bits_btb_entry[2]), .CLK(n43), .Q(ibufBTBResp_entry[2]) );
  DFFX1_LVT ibufBTBResp_entry_reg_1_ ( .D(io_imem_bits_btb_entry[1]), .CLK(n42), .Q(ibufBTBResp_entry[1]) );
  DFFX1_LVT ibufBTBResp_entry_reg_0_ ( .D(io_imem_bits_btb_entry[0]), .CLK(n42), .Q(ibufBTBResp_entry[0]) );
  DFFX1_LVT buf__replay_reg ( .D(io_imem_bits_replay), .CLK(n42), .Q(
        buf__replay) );
  DFFX1_LVT buf__pc_reg_39_ ( .D(io_imem_bits_pc[39]), .CLK(n42), .Q(
        buf__pc[39]) );
  DFFX1_LVT buf__pc_reg_38_ ( .D(io_imem_bits_pc[38]), .CLK(n42), .Q(
        buf__pc[38]) );
  DFFX1_LVT buf__pc_reg_37_ ( .D(io_imem_bits_pc[37]), .CLK(n42), .Q(
        buf__pc[37]) );
  DFFX1_LVT buf__pc_reg_36_ ( .D(io_imem_bits_pc[36]), .CLK(n42), .Q(
        buf__pc[36]) );
  DFFX1_LVT buf__pc_reg_35_ ( .D(io_imem_bits_pc[35]), .CLK(n42), .Q(
        buf__pc[35]) );
  DFFX1_LVT buf__pc_reg_34_ ( .D(io_imem_bits_pc[34]), .CLK(n42), .Q(
        buf__pc[34]) );
  DFFX1_LVT buf__pc_reg_33_ ( .D(io_imem_bits_pc[33]), .CLK(n42), .Q(
        buf__pc[33]) );
  DFFX1_LVT buf__pc_reg_32_ ( .D(io_imem_bits_pc[32]), .CLK(n42), .Q(
        buf__pc[32]) );
  DFFX1_LVT buf__pc_reg_31_ ( .D(io_imem_bits_pc[31]), .CLK(n42), .Q(
        buf__pc[31]) );
  DFFX1_LVT buf__pc_reg_30_ ( .D(io_imem_bits_pc[30]), .CLK(n41), .Q(
        buf__pc[30]) );
  DFFX1_LVT buf__pc_reg_29_ ( .D(io_imem_bits_pc[29]), .CLK(n41), .Q(
        buf__pc[29]) );
  DFFX1_LVT buf__pc_reg_28_ ( .D(io_imem_bits_pc[28]), .CLK(n41), .Q(
        buf__pc[28]) );
  DFFX1_LVT buf__pc_reg_27_ ( .D(io_imem_bits_pc[27]), .CLK(n41), .Q(
        buf__pc[27]) );
  DFFX1_LVT buf__pc_reg_26_ ( .D(io_imem_bits_pc[26]), .CLK(n41), .Q(
        buf__pc[26]) );
  DFFX1_LVT buf__pc_reg_25_ ( .D(io_imem_bits_pc[25]), .CLK(n41), .Q(
        buf__pc[25]) );
  DFFX1_LVT buf__pc_reg_24_ ( .D(io_imem_bits_pc[24]), .CLK(n41), .Q(
        buf__pc[24]) );
  DFFX1_LVT buf__pc_reg_23_ ( .D(io_imem_bits_pc[23]), .CLK(n41), .Q(
        buf__pc[23]) );
  DFFX1_LVT buf__pc_reg_22_ ( .D(io_imem_bits_pc[22]), .CLK(n41), .Q(
        buf__pc[22]) );
  DFFX1_LVT buf__pc_reg_21_ ( .D(io_imem_bits_pc[21]), .CLK(n41), .Q(
        buf__pc[21]) );
  DFFX1_LVT buf__pc_reg_20_ ( .D(io_imem_bits_pc[20]), .CLK(n41), .Q(
        buf__pc[20]) );
  DFFX1_LVT buf__pc_reg_19_ ( .D(io_imem_bits_pc[19]), .CLK(n41), .Q(
        buf__pc[19]) );
  DFFX1_LVT buf__pc_reg_18_ ( .D(io_imem_bits_pc[18]), .CLK(n39), .Q(
        buf__pc[18]) );
  DFFX1_LVT buf__pc_reg_17_ ( .D(io_imem_bits_pc[17]), .CLK(n39), .Q(
        buf__pc[17]) );
  DFFX1_LVT buf__pc_reg_16_ ( .D(io_imem_bits_pc[16]), .CLK(n39), .Q(
        buf__pc[16]) );
  DFFX1_LVT buf__pc_reg_15_ ( .D(io_imem_bits_pc[15]), .CLK(n39), .Q(
        buf__pc[15]) );
  DFFX1_LVT buf__pc_reg_14_ ( .D(io_imem_bits_pc[14]), .CLK(n39), .Q(
        buf__pc[14]) );
  DFFX1_LVT buf__pc_reg_13_ ( .D(io_imem_bits_pc[13]), .CLK(n39), .Q(
        buf__pc[13]) );
  DFFX1_LVT buf__pc_reg_12_ ( .D(io_imem_bits_pc[12]), .CLK(n39), .Q(
        buf__pc[12]) );
  DFFX1_LVT buf__pc_reg_11_ ( .D(io_imem_bits_pc[11]), .CLK(n39), .Q(
        buf__pc[11]) );
  DFFX1_LVT buf__pc_reg_10_ ( .D(io_imem_bits_pc[10]), .CLK(n39), .Q(
        buf__pc[10]) );
  DFFX1_LVT buf__pc_reg_9_ ( .D(io_imem_bits_pc[9]), .CLK(n39), .Q(buf__pc[9])
         );
  DFFX1_LVT buf__pc_reg_8_ ( .D(io_imem_bits_pc[8]), .CLK(n39), .Q(buf__pc[8])
         );
  DFFX1_LVT buf__pc_reg_7_ ( .D(io_imem_bits_pc[7]), .CLK(n39), .Q(buf__pc[7])
         );
  DFFX1_LVT buf__pc_reg_6_ ( .D(io_imem_bits_pc[6]), .CLK(n38), .Q(buf__pc[6])
         );
  DFFX1_LVT buf__pc_reg_5_ ( .D(io_imem_bits_pc[5]), .CLK(n38), .Q(buf__pc[5])
         );
  DFFX1_LVT buf__pc_reg_4_ ( .D(io_imem_bits_pc[4]), .CLK(n38), .Q(buf__pc[4])
         );
  DFFX1_LVT buf__pc_reg_3_ ( .D(io_imem_bits_pc[3]), .CLK(n38), .Q(buf__pc[3])
         );
  DFFX1_LVT buf__pc_reg_2_ ( .D(io_imem_bits_pc[2]), .CLK(n38), .Q(buf__pc[2])
         );
  DFFX1_LVT buf__pc_reg_1_ ( .D(n_T_27_0_), .CLK(n38), .Q(buf__pc[1]) );
  DFFX1_LVT buf__pc_reg_0_ ( .D(io_imem_bits_pc[0]), .CLK(n38), .Q(buf__pc[0])
         );
  DFFX1_LVT buf__data_reg_15_ ( .D(n_T_34[15]), .CLK(n38), .Q(buf__data[15])
         );
  DFFX1_LVT buf__data_reg_14_ ( .D(n_T_34[14]), .CLK(n38), .Q(buf__data[14])
         );
  DFFX1_LVT buf__data_reg_13_ ( .D(n_T_34[13]), .CLK(n38), .Q(buf__data[13])
         );
  DFFX1_LVT buf__data_reg_12_ ( .D(n_T_34[12]), .CLK(n38), .Q(buf__data[12])
         );
  DFFX1_LVT buf__data_reg_11_ ( .D(n_T_34[11]), .CLK(n38), .Q(buf__data[11])
         );
  DFFX1_LVT buf__data_reg_10_ ( .D(n_T_34[10]), .CLK(n37), .Q(buf__data[10])
         );
  DFFX1_LVT buf__data_reg_9_ ( .D(n_T_34[9]), .CLK(n37), .Q(buf__data[9]) );
  DFFX1_LVT buf__data_reg_8_ ( .D(n_T_34[8]), .CLK(n37), .Q(buf__data[8]) );
  DFFX1_LVT buf__data_reg_7_ ( .D(n_T_34[7]), .CLK(n37), .Q(buf__data[7]) );
  DFFX1_LVT buf__data_reg_6_ ( .D(n_T_34[6]), .CLK(n37), .Q(buf__data[6]) );
  DFFX1_LVT buf__data_reg_5_ ( .D(n_T_34[5]), .CLK(n37), .Q(buf__data[5]) );
  DFFX1_LVT buf__data_reg_4_ ( .D(n_T_34[4]), .CLK(n37), .Q(buf__data[4]) );
  DFFX1_LVT buf__data_reg_3_ ( .D(n_T_34[3]), .CLK(n37), .Q(buf__data[3]) );
  DFFX1_LVT buf__data_reg_2_ ( .D(n_T_34[2]), .CLK(n37), .Q(buf__data[2]) );
  DFFX1_LVT buf__data_reg_1_ ( .D(n_T_34[1]), .CLK(n37), .Q(buf__data[1]) );
  DFFX1_LVT buf__xcpt_pf_inst_reg ( .D(io_imem_bits_xcpt_pf_inst), .CLK(n37), 
        .Q(buf__xcpt_pf_inst) );
  DFFX1_LVT buf__xcpt_ae_inst_reg ( .D(io_imem_bits_xcpt_ae_inst), .CLK(n37), 
        .Q(buf__xcpt_ae_inst) );
  DFFX2_LVT nBufValid_reg ( .D(n40), .CLK(clock), .Q(n34), .QN(n12) );
  MUX21X2_LVT U3 ( .A1(io_imem_bits_data[4]), .A2(io_imem_bits_data[20]), .S0(
        n23), .Y(io_inst_0_bits_raw[20]) );
  MUX21X1_LVT U4 ( .A1(io_imem_bits_data[4]), .A2(io_imem_bits_data[20]), .S0(
        n23), .Y(n_T_55_84_) );
  NAND3X0_LVT U5 ( .A1(n68), .A2(n67), .A3(n66), .Y(io_inst_0_bits_raw[3]) );
  NAND3X2_LVT U6 ( .A1(n77), .A2(n76), .A3(n75), .Y(io_inst_0_bits_raw[6]) );
  NAND3X1_LVT U7 ( .A1(n114), .A2(n12), .A3(io_imem_bits_data[14]), .Y(n98) );
  NAND3X1_LVT U8 ( .A1(n114), .A2(n36), .A3(io_imem_bits_data[0]), .Y(n58) );
  NAND3X0_LVT U9 ( .A1(n98), .A2(n99), .A3(n97), .Y(io_inst_0_bits_raw[14]) );
  AND2X1_LVT U10 ( .A1(io_imem_bits_data[8]), .A2(n12), .Y(n5) );
  NAND3X0_LVT U11 ( .A1(n58), .A2(n59), .A3(n57), .Y(io_inst_0_bits_raw[0]) );
  NAND3X2_LVT U12 ( .A1(n83), .A2(n82), .A3(n81), .Y(io_inst_0_bits_raw[8]) );
  NAND3X0_LVT U13 ( .A1(n12), .A2(n20), .A3(io_imem_bits_data[30]), .Y(n97) );
  AND2X1_LVT U14 ( .A1(n12), .A2(io_imem_bits_data[11]), .Y(n27) );
  AND2X1_LVT U15 ( .A1(n12), .A2(io_imem_bits_data[10]), .Y(n30) );
  AND2X1_LVT U16 ( .A1(n12), .A2(io_imem_bits_data[7]), .Y(n31) );
  AND2X1_LVT U17 ( .A1(n12), .A2(io_imem_bits_data[6]), .Y(n26) );
  AND2X1_LVT U18 ( .A1(n12), .A2(io_imem_bits_data[4]), .Y(n24) );
  MUX21X1_LVT U19 ( .A1(buf__pc[39]), .A2(io_imem_bits_pc[39]), .S0(n36), .Y(
        io_pc[39]) );
  MUX21X1_LVT U20 ( .A1(buf__pc[38]), .A2(io_imem_bits_pc[38]), .S0(n36), .Y(
        io_pc[38]) );
  MUX21X1_LVT U21 ( .A1(buf__pc[37]), .A2(io_imem_bits_pc[37]), .S0(n36), .Y(
        io_pc[37]) );
  MUX21X1_LVT U22 ( .A1(buf__pc[36]), .A2(io_imem_bits_pc[36]), .S0(n36), .Y(
        io_pc[36]) );
  MUX21X1_LVT U23 ( .A1(buf__pc[35]), .A2(io_imem_bits_pc[35]), .S0(n36), .Y(
        io_pc[35]) );
  MUX21X1_LVT U24 ( .A1(buf__pc[34]), .A2(io_imem_bits_pc[34]), .S0(n36), .Y(
        io_pc[34]) );
  MUX21X1_LVT U25 ( .A1(buf__pc[33]), .A2(io_imem_bits_pc[33]), .S0(n36), .Y(
        io_pc[33]) );
  MUX21X1_LVT U26 ( .A1(buf__pc[32]), .A2(io_imem_bits_pc[32]), .S0(n36), .Y(
        io_pc[32]) );
  MUX21X1_LVT U27 ( .A1(buf__pc[31]), .A2(io_imem_bits_pc[31]), .S0(n36), .Y(
        io_pc[31]) );
  MUX21X1_LVT U28 ( .A1(buf__pc[30]), .A2(io_imem_bits_pc[30]), .S0(n36), .Y(
        io_pc[30]) );
  MUX21X1_LVT U29 ( .A1(buf__pc[29]), .A2(io_imem_bits_pc[29]), .S0(n36), .Y(
        io_pc[29]) );
  MUX21X1_LVT U30 ( .A1(buf__pc[28]), .A2(io_imem_bits_pc[28]), .S0(n36), .Y(
        io_pc[28]) );
  MUX21X1_LVT U31 ( .A1(buf__pc[27]), .A2(io_imem_bits_pc[27]), .S0(n36), .Y(
        io_pc[27]) );
  MUX21X1_LVT U32 ( .A1(buf__pc[26]), .A2(io_imem_bits_pc[26]), .S0(n36), .Y(
        io_pc[26]) );
  MUX21X1_LVT U33 ( .A1(buf__pc[25]), .A2(io_imem_bits_pc[25]), .S0(n36), .Y(
        io_pc[25]) );
  MUX21X1_LVT U34 ( .A1(buf__pc[24]), .A2(io_imem_bits_pc[24]), .S0(n36), .Y(
        io_pc[24]) );
  MUX21X1_LVT U35 ( .A1(buf__pc[23]), .A2(io_imem_bits_pc[23]), .S0(n36), .Y(
        io_pc[23]) );
  MUX21X1_LVT U36 ( .A1(buf__pc[22]), .A2(io_imem_bits_pc[22]), .S0(n36), .Y(
        io_pc[22]) );
  MUX21X1_LVT U37 ( .A1(buf__pc[21]), .A2(io_imem_bits_pc[21]), .S0(n36), .Y(
        io_pc[21]) );
  MUX21X1_LVT U38 ( .A1(buf__pc[20]), .A2(io_imem_bits_pc[20]), .S0(n36), .Y(
        io_pc[20]) );
  MUX21X1_LVT U39 ( .A1(buf__pc[19]), .A2(io_imem_bits_pc[19]), .S0(n36), .Y(
        io_pc[19]) );
  MUX21X1_LVT U40 ( .A1(buf__pc[18]), .A2(io_imem_bits_pc[18]), .S0(n36), .Y(
        io_pc[18]) );
  MUX21X1_LVT U41 ( .A1(buf__pc[17]), .A2(io_imem_bits_pc[17]), .S0(n36), .Y(
        io_pc[17]) );
  MUX21X1_LVT U42 ( .A1(buf__pc[16]), .A2(io_imem_bits_pc[16]), .S0(n36), .Y(
        io_pc[16]) );
  MUX21X1_LVT U43 ( .A1(buf__pc[15]), .A2(io_imem_bits_pc[15]), .S0(n36), .Y(
        io_pc[15]) );
  MUX21X1_LVT U44 ( .A1(buf__pc[14]), .A2(io_imem_bits_pc[14]), .S0(n36), .Y(
        io_pc[14]) );
  MUX21X1_LVT U45 ( .A1(buf__pc[13]), .A2(io_imem_bits_pc[13]), .S0(n36), .Y(
        io_pc[13]) );
  MUX21X1_LVT U46 ( .A1(buf__pc[12]), .A2(io_imem_bits_pc[12]), .S0(n36), .Y(
        io_pc[12]) );
  MUX21X1_LVT U47 ( .A1(buf__pc[11]), .A2(io_imem_bits_pc[11]), .S0(n36), .Y(
        io_pc[11]) );
  MUX21X1_LVT U48 ( .A1(buf__pc[10]), .A2(io_imem_bits_pc[10]), .S0(n36), .Y(
        io_pc[10]) );
  MUX21X1_LVT U49 ( .A1(buf__pc[9]), .A2(io_imem_bits_pc[9]), .S0(n36), .Y(
        io_pc[9]) );
  MUX21X1_LVT U50 ( .A1(buf__pc[8]), .A2(io_imem_bits_pc[8]), .S0(n36), .Y(
        io_pc[8]) );
  MUX21X1_LVT U51 ( .A1(buf__pc[7]), .A2(io_imem_bits_pc[7]), .S0(n36), .Y(
        io_pc[7]) );
  MUX21X1_LVT U52 ( .A1(buf__pc[6]), .A2(io_imem_bits_pc[6]), .S0(n36), .Y(
        io_pc[6]) );
  MUX21X1_LVT U53 ( .A1(buf__pc[5]), .A2(io_imem_bits_pc[5]), .S0(n36), .Y(
        io_pc[5]) );
  MUX21X1_LVT U54 ( .A1(buf__pc[4]), .A2(io_imem_bits_pc[4]), .S0(n36), .Y(
        io_pc[4]) );
  NAND2X0_LVT U55 ( .A1(n35), .A2(n114), .Y(n7) );
  AND2X1_LVT U56 ( .A1(n12), .A2(n7), .Y(n8) );
  NAND2X0_LVT U57 ( .A1(n20), .A2(n96), .Y(n9) );
  AO22X2_LVT U58 ( .A1(buf__data[13]), .A2(n34), .A3(n8), .A4(n9), .Y(n125) );
  NAND2X4_LVT U59 ( .A1(n105), .A2(n104), .Y(n123) );
  OR2X2_LVT U60 ( .A1(n20), .A2(n12), .Y(n10) );
  OR2X2_LVT U61 ( .A1(n20), .A2(n12), .Y(n11) );
  OR2X1_LVT U62 ( .A1(n20), .A2(n12), .Y(n106) );
  MUX21X2_LVT U63 ( .A1(io_imem_bits_data[15]), .A2(io_imem_bits_data[31]), 
        .S0(n106), .Y(io_inst_0_bits_raw[31]) );
  NAND3X1_LVT U64 ( .A1(n12), .A2(n20), .A3(io_imem_bits_data[17]), .Y(n60) );
  NAND3X2_LVT U65 ( .A1(n89), .A2(n88), .A3(n87), .Y(n127) );
  NAND3X0_LVT U66 ( .A1(n95), .A2(n94), .A3(n93), .Y(io_inst_0_bits_raw[12])
         );
  NAND3X0_LVT U67 ( .A1(n95), .A2(n94), .A3(n93), .Y(n126) );
  MUX21X2_LVT U68 ( .A1(io_imem_bits_data[12]), .A2(io_imem_bits_data[28]), 
        .S0(n10), .Y(io_inst_0_bits_raw[28]) );
  NBUFFX2_LVT U69 ( .A(n123), .Y(io_inst_0_bits_raw[15]) );
  NAND3X1_LVT U70 ( .A1(n114), .A2(n12), .A3(io_imem_bits_data[1]), .Y(n61) );
  NAND3X0_LVT U71 ( .A1(n90), .A2(n91), .A3(n92), .Y(io_inst_0_bits_raw[11])
         );
  NAND2X0_LVT U72 ( .A1(n56), .A2(n55), .Y(n100) );
  INVX1_LVT U73 ( .A(n122), .Y(io_inst_0_bits_rvc) );
  INVX0_LVT U74 ( .A(N51), .Y(n51) );
  INVX0_LVT U75 ( .A(n117), .Y(n49) );
  NAND2X0_LVT U76 ( .A1(n47), .A2(n113), .Y(n117) );
  NAND3X0_LVT U77 ( .A1(n80), .A2(n79), .A3(n78), .Y(io_inst_0_bits_raw[7]) );
  NAND3X0_LVT U78 ( .A1(n77), .A2(n76), .A3(n75), .Y(n128) );
  NAND3X0_LVT U79 ( .A1(n74), .A2(n73), .A3(n72), .Y(io_inst_0_bits_raw[5]) );
  NAND3X0_LVT U80 ( .A1(n69), .A2(n70), .A3(n71), .Y(io_inst_0_bits_raw[4]) );
  MUX21X1_LVT U81 ( .A1(io_imem_bits_data[13]), .A2(io_imem_bits_data[29]), 
        .S0(n23), .Y(io_inst_0_bits_raw[29]) );
  MUX21X1_LVT U82 ( .A1(io_imem_bits_data[14]), .A2(io_imem_bits_data[30]), 
        .S0(n11), .Y(io_inst_0_bits_raw[30]) );
  INVX0_LVT U83 ( .A(n116), .Y(n118) );
  INVX0_LVT U84 ( .A(n25), .Y(n19) );
  INVX0_LVT U85 ( .A(io_imem_bits_btb_bridx), .Y(n45) );
  NAND3X0_LVT U86 ( .A1(n98), .A2(n99), .A3(n97), .Y(n124) );
  NBUFFX2_LVT U87 ( .A(n_T_55_85_), .Y(io_inst_0_bits_raw[21]) );
  NAND3X0_LVT U88 ( .A1(n62), .A2(n61), .A3(n60), .Y(io_inst_0_bits_raw[1]) );
  NBUFFX2_LVT U89 ( .A(n125), .Y(io_inst_0_bits_raw[13]) );
  INVX1_LVT U90 ( .A(n32), .Y(n18) );
  IBUFFX2_LVT U91 ( .A(io_imem_bits_data[31]), .Y(n101) );
  NAND3X0_LVT U92 ( .A1(n12), .A2(n20), .A3(io_imem_bits_data[16]), .Y(n57) );
  OR2X1_LVT U93 ( .A1(n20), .A2(io_imem_bits_data[15]), .Y(n102) );
  AO21X1_LVT U94 ( .A1(io_imem_bits_btb_taken), .A2(n45), .A3(n19), .Y(n116)
         );
  NBUFFX2_LVT U95 ( .A(io_imem_bits_pc[1]), .Y(n20) );
  NAND2X0_LVT U96 ( .A1(n33), .A2(n86), .Y(io_inst_0_bits_raw[9]) );
  NBUFFX2_LVT U97 ( .A(n_T_55_91_), .Y(io_inst_0_bits_raw[27]) );
  MUX21X1_LVT U98 ( .A1(io_imem_bits_data[11]), .A2(io_imem_bits_data[27]), 
        .S0(n11), .Y(n_T_55_91_) );
  AND2X1_LVT U99 ( .A1(n114), .A2(n12), .Y(n28) );
  NBUFFX2_LVT U100 ( .A(n127), .Y(io_inst_0_bits_raw[10]) );
  NBUFFX2_LVT U101 ( .A(n10), .Y(n23) );
  INVX1_LVT U102 ( .A(n32), .Y(n115) );
  NAND2X0_LVT U103 ( .A1(n24), .A2(n114), .Y(n71) );
  NBUFFX2_LVT U104 ( .A(n114), .Y(n25) );
  NAND3X0_LVT U105 ( .A1(n62), .A2(n61), .A3(n60), .Y(n130) );
  NAND2X0_LVT U106 ( .A1(n25), .A2(n26), .Y(n77) );
  NAND2X0_LVT U107 ( .A1(n27), .A2(n114), .Y(n92) );
  NBUFFX2_LVT U108 ( .A(n11), .Y(n29) );
  MUX21X1_LVT U109 ( .A1(io_imem_bits_data[1]), .A2(io_imem_bits_data[17]), 
        .S0(n29), .Y(io_inst_0_bits_raw[17]) );
  MUX21X1_LVT U110 ( .A1(io_imem_bits_data[10]), .A2(io_imem_bits_data[26]), 
        .S0(n29), .Y(io_inst_0_bits_raw[26]) );
  MUX21X1_LVT U111 ( .A1(io_imem_bits_data[6]), .A2(io_imem_bits_data[22]), 
        .S0(n10), .Y(io_inst_0_bits_raw[22]) );
  MUX21X1_LVT U112 ( .A1(io_imem_bits_data[7]), .A2(io_imem_bits_data[23]), 
        .S0(n10), .Y(io_inst_0_bits_raw[23]) );
  MUX21X1_LVT U113 ( .A1(io_imem_bits_data[8]), .A2(io_imem_bits_data[24]), 
        .S0(n11), .Y(io_inst_0_bits_raw[24]) );
  MUX21X1_LVT U114 ( .A1(io_imem_bits_data[5]), .A2(io_imem_bits_data[21]), 
        .S0(n11), .Y(n_T_55_85_) );
  NAND2X0_LVT U115 ( .A1(n25), .A2(n30), .Y(n89) );
  NAND2X0_LVT U116 ( .A1(n31), .A2(n114), .Y(n80) );
  NAND2X0_LVT U117 ( .A1(n12), .A2(io_imem_bits_pc[1]), .Y(n32) );
  AND2X1_LVT U118 ( .A1(n85), .A2(n84), .Y(n33) );
  AO21X2_LVT U119 ( .A1(buf__pc[1]), .A2(n34), .A3(n18), .Y(io_pc[1]) );
  INVX1_LVT U120 ( .A(io_imem_bits_data[29]), .Y(n96) );
  INVX1_LVT U121 ( .A(io_imem_bits_data[13]), .Y(n35) );
  IBUFFX2_LVT U122 ( .A(io_imem_bits_pc[1]), .Y(n114) );
  NBUFFX2_LVT U123 ( .A(net35341), .Y(n43) );
  NBUFFX2_LVT U124 ( .A(net35341), .Y(n42) );
  NBUFFX2_LVT U125 ( .A(net35341), .Y(n41) );
  NBUFFX2_LVT U126 ( .A(net35341), .Y(n39) );
  NBUFFX2_LVT U127 ( .A(net35341), .Y(n38) );
  NBUFFX2_LVT U128 ( .A(net35341), .Y(n37) );
  MUX21X1_LVT U129 ( .A1(io_imem_bits_data[5]), .A2(io_imem_bits_data[21]), 
        .S0(n100), .Y(n_T_34[5]) );
  MUX21X1_LVT U130 ( .A1(io_imem_bits_data[12]), .A2(io_imem_bits_data[28]), 
        .S0(n100), .Y(n_T_34[12]) );
  MUX21X1_LVT U131 ( .A1(io_imem_bits_data[3]), .A2(io_imem_bits_data[19]), 
        .S0(n100), .Y(n_T_34[3]) );
  MUX21X1_LVT U132 ( .A1(io_imem_bits_data[15]), .A2(io_imem_bits_data[31]), 
        .S0(n100), .Y(n_T_34[15]) );
  MUX21X1_LVT U133 ( .A1(io_imem_bits_data[6]), .A2(io_imem_bits_data[22]), 
        .S0(n100), .Y(n_T_34[6]) );
  MUX21X1_LVT U134 ( .A1(io_imem_bits_data[1]), .A2(io_imem_bits_data[17]), 
        .S0(n100), .Y(n_T_34[1]) );
  MUX21X1_LVT U135 ( .A1(io_imem_bits_data[7]), .A2(io_imem_bits_data[23]), 
        .S0(n100), .Y(n_T_34[7]) );
  MUX21X1_LVT U136 ( .A1(io_imem_bits_data[14]), .A2(io_imem_bits_data[30]), 
        .S0(n100), .Y(n_T_34[14]) );
  MUX21X1_LVT U137 ( .A1(io_imem_bits_data[2]), .A2(io_imem_bits_data[18]), 
        .S0(n100), .Y(n_T_34[2]) );
  MUX21X1_LVT U138 ( .A1(io_imem_bits_data[11]), .A2(io_imem_bits_data[27]), 
        .S0(n100), .Y(n_T_34[11]) );
  MUX21X1_LVT U139 ( .A1(io_imem_bits_data[8]), .A2(io_imem_bits_data[24]), 
        .S0(n100), .Y(n_T_34[8]) );
  MUX21X1_LVT U140 ( .A1(io_imem_bits_data[4]), .A2(io_imem_bits_data[20]), 
        .S0(n100), .Y(n_T_34[4]) );
  MUX21X1_LVT U141 ( .A1(io_imem_bits_data[9]), .A2(io_imem_bits_data[25]), 
        .S0(n100), .Y(n_T_34[9]) );
  MUX21X1_LVT U142 ( .A1(io_imem_bits_data[10]), .A2(io_imem_bits_data[26]), 
        .S0(n100), .Y(n_T_34[10]) );
  MUX21X1_LVT U143 ( .A1(io_imem_bits_data[0]), .A2(io_imem_bits_data[16]), 
        .S0(n100), .Y(n_T_34[0]) );
  MUX21X1_LVT U144 ( .A1(io_imem_bits_data[13]), .A2(io_imem_bits_data[29]), 
        .S0(n100), .Y(n_T_34[13]) );
  MUX21X1_LVT U145 ( .A1(buf__pc[2]), .A2(io_imem_bits_pc[2]), .S0(n12), .Y(
        io_pc[2]) );
  MUX21X1_LVT U146 ( .A1(buf__pc[0]), .A2(io_imem_bits_pc[0]), .S0(n12), .Y(
        io_pc[0]) );
  MUX21X1_LVT U147 ( .A1(buf__pc[3]), .A2(io_imem_bits_pc[3]), .S0(n12), .Y(
        io_pc[3]) );
  MUX21X1_LVT U148 ( .A1(io_imem_bits_data[9]), .A2(io_imem_bits_data[25]), 
        .S0(n29), .Y(io_inst_0_bits_raw[25]) );
  NAND3X0_LVT U149 ( .A1(n68), .A2(n67), .A3(n66), .Y(n129) );
  MUX21X1_LVT U150 ( .A1(ibufBTBResp_bht_history[7]), .A2(
        io_imem_bits_btb_bht_history[7]), .S0(n113), .Y(
        io_btb_resp_bht_history[7]) );
  MUX21X1_LVT U151 ( .A1(ibufBTBResp_entry[1]), .A2(io_imem_bits_btb_entry[1]), 
        .S0(n113), .Y(io_btb_resp_entry[1]) );
  MUX21X1_LVT U152 ( .A1(ibufBTBResp_entry[0]), .A2(io_imem_bits_btb_entry[0]), 
        .S0(n113), .Y(io_btb_resp_entry[0]) );
  MUX21X1_LVT U153 ( .A1(ibufBTBResp_bht_history[1]), .A2(
        io_imem_bits_btb_bht_history[1]), .S0(n113), .Y(
        io_btb_resp_bht_history[1]) );
  MUX21X1_LVT U154 ( .A1(ibufBTBResp_entry[2]), .A2(io_imem_bits_btb_entry[2]), 
        .S0(n113), .Y(io_btb_resp_entry[2]) );
  MUX21X1_LVT U155 ( .A1(ibufBTBResp_entry[3]), .A2(io_imem_bits_btb_entry[3]), 
        .S0(n113), .Y(io_btb_resp_entry[3]) );
  MUX21X1_LVT U156 ( .A1(ibufBTBResp_bht_history[2]), .A2(
        io_imem_bits_btb_bht_history[2]), .S0(n113), .Y(
        io_btb_resp_bht_history[2]) );
  MUX21X1_LVT U157 ( .A1(ibufBTBResp_bht_history[4]), .A2(
        io_imem_bits_btb_bht_history[4]), .S0(n113), .Y(
        io_btb_resp_bht_history[4]) );
  MUX21X1_LVT U158 ( .A1(ibufBTBResp_bht_history[0]), .A2(
        io_imem_bits_btb_bht_history[0]), .S0(n113), .Y(
        io_btb_resp_bht_history[0]) );
  MUX21X1_LVT U159 ( .A1(ibufBTBResp_entry[4]), .A2(io_imem_bits_btb_entry[4]), 
        .S0(n113), .Y(io_btb_resp_entry[4]) );
  MUX21X1_LVT U160 ( .A1(ibufBTBResp_bht_history[5]), .A2(
        io_imem_bits_btb_bht_history[5]), .S0(n113), .Y(
        io_btb_resp_bht_history[5]) );
  MUX21X1_LVT U161 ( .A1(ibufBTBResp_bht_history[3]), .A2(
        io_imem_bits_btb_bht_history[3]), .S0(n113), .Y(
        io_btb_resp_bht_history[3]) );
  MUX21X1_LVT U162 ( .A1(ibufBTBResp_bht_history[6]), .A2(
        io_imem_bits_btb_bht_history[6]), .S0(n113), .Y(
        io_btb_resp_bht_history[6]) );
  XOR2X1_LVT U163 ( .A1(n117), .A2(n25), .Y(n_T_27_0_) );
  MUX21X1_LVT U164 ( .A1(n19), .A2(n117), .S0(n119), .Y(n56) );
  INVX1_LVT U165 ( .A(n34), .Y(n36) );
  NAND2X4_LVT U166 ( .A1(io_inst_0_bits_rvc), .A2(n34), .Y(n113) );
  NAND3X0_LVT U167 ( .A1(n102), .A2(n12), .A3(n103), .Y(n105) );
  NAND2X0_LVT U168 ( .A1(buf__data[1]), .A2(n34), .Y(n62) );
  NAND3X0_LVT U169 ( .A1(n58), .A2(n59), .A3(n57), .Y(n131) );
  NAND2X0_LVT U170 ( .A1(buf__data[0]), .A2(n34), .Y(n59) );
  NAND3X0_LVT U171 ( .A1(n45), .A2(io_imem_bits_btb_taken), .A3(n19), .Y(n107)
         );
  NAND2X0_LVT U172 ( .A1(io_imem_valid), .A2(n107), .Y(n110) );
  AO21X1_LVT U173 ( .A1(n12), .A2(n116), .A3(n110), .Y(n54) );
  NAND2X0_LVT U174 ( .A1(n34), .A2(buf__replay), .Y(n108) );
  NAND2X0_LVT U175 ( .A1(n54), .A2(n108), .Y(n46) );
  OR2X1_LVT U176 ( .A1(n46), .A2(io_inst_0_bits_rvc), .Y(n112) );
  OR2X1_LVT U177 ( .A1(n12), .A2(n112), .Y(n121) );
  OA21X1_LVT U178 ( .A1(n12), .A2(io_inst_0_ready), .A3(n121), .Y(n52) );
  OR2X1_LVT U179 ( .A1(n34), .A2(io_inst_0_bits_rvc), .Y(n47) );
  AND2X1_LVT U180 ( .A1(n107), .A2(n117), .Y(n48) );
  MUX21X1_LVT U181 ( .A1(n49), .A2(n48), .S0(n116), .Y(n50) );
  AND3X1_LVT U182 ( .A1(n50), .A2(io_imem_valid), .A3(io_inst_0_ready), .Y(N51) );
  AO21X1_LVT U183 ( .A1(n51), .A2(n52), .A3(reset), .Y(n53) );
  NOR2X0_LVT U184 ( .A1(n53), .A2(io_kill), .Y(n40) );
  OA21X1_LVT U185 ( .A1(n54), .A2(n34), .A3(n121), .Y(n119) );
  NAND2X0_LVT U186 ( .A1(n117), .A2(n19), .Y(n55) );
  NAND2X0_LVT U187 ( .A1(io_imem_bits_data[2]), .A2(n28), .Y(n65) );
  NAND2X0_LVT U188 ( .A1(buf__data[2]), .A2(n34), .Y(n64) );
  NAND2X0_LVT U189 ( .A1(io_imem_bits_data[18]), .A2(n115), .Y(n63) );
  NAND3X0_LVT U190 ( .A1(n65), .A2(n64), .A3(n63), .Y(io_inst_0_bits_raw[2])
         );
  NAND2X0_LVT U191 ( .A1(io_imem_bits_data[3]), .A2(n28), .Y(n68) );
  NAND2X0_LVT U192 ( .A1(buf__data[3]), .A2(n34), .Y(n67) );
  NAND2X0_LVT U193 ( .A1(io_imem_bits_data[19]), .A2(n18), .Y(n66) );
  NAND2X0_LVT U194 ( .A1(n34), .A2(buf__data[4]), .Y(n70) );
  NAND2X0_LVT U195 ( .A1(io_imem_bits_data[20]), .A2(n115), .Y(n69) );
  NAND2X0_LVT U196 ( .A1(n28), .A2(io_imem_bits_data[5]), .Y(n74) );
  NAND2X0_LVT U197 ( .A1(buf__data[5]), .A2(n34), .Y(n73) );
  NAND2X0_LVT U198 ( .A1(io_imem_bits_data[21]), .A2(n18), .Y(n72) );
  NAND2X0_LVT U199 ( .A1(buf__data[6]), .A2(n34), .Y(n76) );
  NAND2X0_LVT U200 ( .A1(io_imem_bits_data[22]), .A2(n115), .Y(n75) );
  NAND2X0_LVT U201 ( .A1(buf__data[7]), .A2(n34), .Y(n79) );
  NAND2X0_LVT U202 ( .A1(io_imem_bits_data[23]), .A2(n115), .Y(n78) );
  NAND2X0_LVT U203 ( .A1(n5), .A2(n114), .Y(n83) );
  NAND2X0_LVT U204 ( .A1(buf__data[8]), .A2(n34), .Y(n82) );
  NAND2X0_LVT U205 ( .A1(io_imem_bits_data[24]), .A2(n18), .Y(n81) );
  NAND2X0_LVT U206 ( .A1(io_imem_bits_data[9]), .A2(n28), .Y(n86) );
  NAND2X0_LVT U207 ( .A1(buf__data[9]), .A2(n34), .Y(n85) );
  NAND2X0_LVT U208 ( .A1(io_imem_bits_data[25]), .A2(n115), .Y(n84) );
  NAND2X0_LVT U209 ( .A1(buf__data[10]), .A2(n34), .Y(n88) );
  NAND2X0_LVT U210 ( .A1(io_imem_bits_data[26]), .A2(n18), .Y(n87) );
  NAND2X0_LVT U211 ( .A1(buf__data[11]), .A2(n34), .Y(n91) );
  NAND2X0_LVT U212 ( .A1(io_imem_bits_data[27]), .A2(n115), .Y(n90) );
  NAND2X0_LVT U213 ( .A1(io_imem_bits_data[12]), .A2(n28), .Y(n95) );
  NAND2X0_LVT U214 ( .A1(buf__data[12]), .A2(n34), .Y(n94) );
  NAND2X0_LVT U215 ( .A1(io_imem_bits_data[28]), .A2(n18), .Y(n93) );
  NAND2X0_LVT U216 ( .A1(buf__data[14]), .A2(n34), .Y(n99) );
  NAND2X0_LVT U217 ( .A1(n101), .A2(n20), .Y(n103) );
  NAND2X0_LVT U218 ( .A1(n34), .A2(buf__data[15]), .Y(n104) );
  MUX21X1_LVT U219 ( .A1(io_imem_bits_data[0]), .A2(io_imem_bits_data[16]), 
        .S0(n29), .Y(io_inst_0_bits_raw[16]) );
  MUX21X1_LVT U220 ( .A1(io_imem_bits_data[2]), .A2(io_imem_bits_data[18]), 
        .S0(n23), .Y(io_inst_0_bits_raw[18]) );
  MUX21X1_LVT U221 ( .A1(io_imem_bits_data[3]), .A2(io_imem_bits_data[19]), 
        .S0(n29), .Y(io_inst_0_bits_raw[19]) );
  NAND4X0_LVT U222 ( .A1(n113), .A2(io_imem_valid), .A3(io_imem_bits_replay), 
        .A4(n107), .Y(n109) );
  NAND2X0_LVT U223 ( .A1(n109), .A2(n108), .Y(io_inst_0_bits_replay) );
  AND2X1_LVT U224 ( .A1(io_imem_bits_xcpt_ae_inst), .A2(n122), .Y(
        io_inst_0_bits_xcpt1_ae_inst) );
  AND2X1_LVT U225 ( .A1(io_imem_bits_xcpt_pf_inst), .A2(n122), .Y(
        io_inst_0_bits_xcpt1_pf_inst) );
  MUX21X1_LVT U226 ( .A1(buf__xcpt_ae_inst), .A2(io_imem_bits_xcpt_ae_inst), 
        .S0(n12), .Y(io_inst_0_bits_xcpt0_ae_inst) );
  MUX21X1_LVT U227 ( .A1(buf__xcpt_pf_inst), .A2(io_imem_bits_xcpt_pf_inst), 
        .S0(n12), .Y(io_inst_0_bits_xcpt0_pf_inst) );
  NAND2X0_LVT U228 ( .A1(n110), .A2(n12), .Y(n111) );
  AND2X1_LVT U229 ( .A1(n112), .A2(n111), .Y(io_inst_0_valid) );
  NAND3X0_LVT U230 ( .A1(n119), .A2(n118), .A3(n117), .Y(n120) );
  AND3X1_LVT U231 ( .A1(n120), .A2(n121), .A3(io_inst_0_ready), .Y(
        io_imem_ready) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module CSRFile_DW01_inc_J38_0 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(A[24]), .Y(n159) );
  INVX1_LVT U127 ( .A(n183), .Y(n160) );
  INVX1_LVT U128 ( .A(A[20]), .Y(n161) );
  INVX1_LVT U129 ( .A(n187), .Y(n162) );
  INVX1_LVT U130 ( .A(A[16]), .Y(n163) );
  INVX1_LVT U131 ( .A(n192), .Y(n164) );
  INVX1_LVT U132 ( .A(A[12]), .Y(n165) );
  INVX1_LVT U133 ( .A(n196), .Y(n166) );
  INVX1_LVT U134 ( .A(A[8]), .Y(n167) );
  INVX1_LVT U135 ( .A(n172), .Y(n168) );
  INVX1_LVT U136 ( .A(A[4]), .Y(n169) );
  INVX1_LVT U137 ( .A(n176), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n168), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n168), .A2(n167), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n170), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n169), .A4(n170), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n160), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n160), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n159), .A4(n160), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n162), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n162), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n161), .A4(n162), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n164), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n164), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n164), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n164), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n163), .A4(n164), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n166), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n166), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n166), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n165), .A4(n166), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n168), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n168), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n168), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n170), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_1 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(A[24]), .Y(n159) );
  INVX1_LVT U127 ( .A(n183), .Y(n160) );
  INVX1_LVT U128 ( .A(A[20]), .Y(n161) );
  INVX1_LVT U129 ( .A(n187), .Y(n162) );
  INVX1_LVT U130 ( .A(A[16]), .Y(n163) );
  INVX1_LVT U131 ( .A(n192), .Y(n164) );
  INVX1_LVT U132 ( .A(A[12]), .Y(n165) );
  INVX1_LVT U133 ( .A(n196), .Y(n166) );
  INVX1_LVT U134 ( .A(A[8]), .Y(n167) );
  INVX1_LVT U135 ( .A(n172), .Y(n168) );
  INVX1_LVT U136 ( .A(A[4]), .Y(n169) );
  INVX1_LVT U137 ( .A(n176), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n168), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n168), .A2(n167), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n170), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n169), .A4(n170), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n160), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n160), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n159), .A4(n160), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n162), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n162), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n161), .A4(n162), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n164), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n164), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n164), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n164), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n163), .A4(n164), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n166), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n166), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n166), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n165), .A4(n166), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n168), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n168), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n168), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n170), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_2 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(A[24]), .Y(n159) );
  INVX1_LVT U127 ( .A(n183), .Y(n160) );
  INVX1_LVT U128 ( .A(A[20]), .Y(n161) );
  INVX1_LVT U129 ( .A(n187), .Y(n162) );
  INVX1_LVT U130 ( .A(A[16]), .Y(n163) );
  INVX1_LVT U131 ( .A(n192), .Y(n164) );
  INVX1_LVT U132 ( .A(A[12]), .Y(n165) );
  INVX1_LVT U133 ( .A(n196), .Y(n166) );
  INVX1_LVT U134 ( .A(A[8]), .Y(n167) );
  INVX1_LVT U135 ( .A(n172), .Y(n168) );
  INVX1_LVT U136 ( .A(A[4]), .Y(n169) );
  INVX1_LVT U137 ( .A(n176), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n168), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n168), .A2(n167), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n170), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n169), .A4(n170), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n160), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n160), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n159), .A4(n160), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n162), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n162), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n161), .A4(n162), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n164), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n164), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n164), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n164), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n163), .A4(n164), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n166), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n166), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n166), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n165), .A4(n166), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n168), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n168), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n168), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n170), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_3 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(A[24]), .Y(n159) );
  INVX1_LVT U127 ( .A(n183), .Y(n160) );
  INVX1_LVT U128 ( .A(A[20]), .Y(n161) );
  INVX1_LVT U129 ( .A(n187), .Y(n162) );
  INVX1_LVT U130 ( .A(A[16]), .Y(n163) );
  INVX1_LVT U131 ( .A(n192), .Y(n164) );
  INVX1_LVT U132 ( .A(A[12]), .Y(n165) );
  INVX1_LVT U133 ( .A(n196), .Y(n166) );
  INVX1_LVT U134 ( .A(A[8]), .Y(n167) );
  INVX1_LVT U135 ( .A(n172), .Y(n168) );
  INVX1_LVT U136 ( .A(A[4]), .Y(n169) );
  INVX1_LVT U137 ( .A(n176), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n168), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n168), .A2(n167), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n170), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n169), .A4(n170), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n160), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n160), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n159), .A4(n160), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n162), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n162), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n161), .A4(n162), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n164), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n164), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n164), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n164), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n163), .A4(n164), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n166), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n166), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n166), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n165), .A4(n166), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n168), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n168), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n168), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n170), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_4 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(n183), .Y(n159) );
  INVX1_LVT U127 ( .A(n187), .Y(n160) );
  INVX1_LVT U128 ( .A(n192), .Y(n161) );
  INVX1_LVT U129 ( .A(n196), .Y(n162) );
  INVX1_LVT U130 ( .A(n172), .Y(n163) );
  INVX1_LVT U131 ( .A(n176), .Y(n164) );
  INVX1_LVT U132 ( .A(A[24]), .Y(n165) );
  INVX1_LVT U133 ( .A(A[20]), .Y(n166) );
  INVX1_LVT U134 ( .A(A[16]), .Y(n167) );
  INVX1_LVT U135 ( .A(A[12]), .Y(n168) );
  INVX1_LVT U136 ( .A(A[8]), .Y(n169) );
  INVX1_LVT U137 ( .A(A[4]), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n163), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n163), .A2(n169), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n164), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n170), .A4(n164), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n159), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n159), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n165), .A4(n159), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n160), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n160), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n166), .A4(n160), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n161), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n161), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n161), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n161), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n167), .A4(n161), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n162), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n162), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n162), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n168), .A4(n162), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n163), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n163), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n163), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n164), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_5 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(n183), .Y(n159) );
  INVX1_LVT U127 ( .A(n187), .Y(n160) );
  INVX1_LVT U128 ( .A(n192), .Y(n161) );
  INVX1_LVT U129 ( .A(n196), .Y(n162) );
  INVX1_LVT U130 ( .A(n172), .Y(n163) );
  INVX1_LVT U131 ( .A(n176), .Y(n164) );
  INVX1_LVT U132 ( .A(A[24]), .Y(n165) );
  INVX1_LVT U133 ( .A(A[20]), .Y(n166) );
  INVX1_LVT U134 ( .A(A[16]), .Y(n167) );
  INVX1_LVT U135 ( .A(A[12]), .Y(n168) );
  INVX1_LVT U136 ( .A(A[8]), .Y(n169) );
  INVX1_LVT U137 ( .A(A[4]), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n163), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n163), .A2(n169), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n164), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n170), .A4(n164), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n159), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n159), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n165), .A4(n159), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n160), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n160), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n166), .A4(n160), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n161), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n161), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n161), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n161), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n167), .A4(n161), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n162), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n162), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n162), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n168), .A4(n162), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n163), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n163), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n163), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n164), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_6 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(A[24]), .Y(n159) );
  INVX1_LVT U127 ( .A(n183), .Y(n160) );
  INVX1_LVT U128 ( .A(A[20]), .Y(n161) );
  INVX1_LVT U129 ( .A(n187), .Y(n162) );
  INVX1_LVT U130 ( .A(A[16]), .Y(n163) );
  INVX1_LVT U131 ( .A(n192), .Y(n164) );
  INVX1_LVT U132 ( .A(A[12]), .Y(n165) );
  INVX1_LVT U133 ( .A(n196), .Y(n166) );
  INVX1_LVT U134 ( .A(A[8]), .Y(n167) );
  INVX1_LVT U135 ( .A(n172), .Y(n168) );
  INVX1_LVT U136 ( .A(A[4]), .Y(n169) );
  INVX1_LVT U137 ( .A(n176), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n168), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n168), .A2(n167), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n170), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n169), .A4(n170), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n160), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n160), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n159), .A4(n160), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n162), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n162), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n161), .A4(n162), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n164), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n164), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n164), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n164), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n163), .A4(n164), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n166), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n166), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n166), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n165), .A4(n166), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n168), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n168), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n168), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n170), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_7 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;
  wire   n93, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199;

  HADDX1_LVT U121 ( .A0(A[1]), .B0(A[0]), .C1(n93), .SO(SUM[1]) );
  INVX1_LVT U126 ( .A(n183), .Y(n159) );
  INVX1_LVT U127 ( .A(n187), .Y(n160) );
  INVX1_LVT U128 ( .A(n192), .Y(n161) );
  INVX1_LVT U129 ( .A(n196), .Y(n162) );
  INVX1_LVT U130 ( .A(n172), .Y(n163) );
  INVX1_LVT U131 ( .A(n176), .Y(n164) );
  INVX1_LVT U132 ( .A(A[24]), .Y(n165) );
  INVX1_LVT U133 ( .A(A[20]), .Y(n166) );
  INVX1_LVT U134 ( .A(A[16]), .Y(n167) );
  INVX1_LVT U135 ( .A(A[12]), .Y(n168) );
  INVX1_LVT U136 ( .A(A[8]), .Y(n169) );
  INVX1_LVT U137 ( .A(A[4]), .Y(n170) );
  HADDX1_LVT U138 ( .A0(n171), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U139 ( .A1(A[8]), .A2(n163), .Y(n171) );
  AO22X1_LVT U140 ( .A1(n163), .A2(n169), .A3(n172), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U141 ( .A0(A[7]), .B0(n173), .SO(SUM[7]) );
  AND2X1_LVT U142 ( .A1(A[6]), .A2(n174), .Y(n173) );
  HADDX1_LVT U143 ( .A0(A[6]), .B0(n174), .SO(SUM[6]) );
  HADDX1_LVT U144 ( .A0(n175), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U145 ( .A1(n164), .A2(A[4]), .Y(n175) );
  AO22X1_LVT U146 ( .A1(A[4]), .A2(n176), .A3(n170), .A4(n164), .Y(SUM[4]) );
  HADDX1_LVT U147 ( .A0(A[3]), .B0(n177), .SO(SUM[3]) );
  AND2X1_LVT U148 ( .A1(n93), .A2(A[2]), .Y(n177) );
  HADDX1_LVT U149 ( .A0(n93), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U150 ( .A0(n178), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U151 ( .A1(n179), .A2(A[27]), .A3(A[28]), .Y(n178) );
  HADDX1_LVT U152 ( .A0(n180), .B0(A[28]), .SO(SUM[28]) );
  AND2X1_LVT U153 ( .A1(A[27]), .A2(n179), .Y(n180) );
  HADDX1_LVT U154 ( .A0(A[27]), .B0(n179), .SO(SUM[27]) );
  AND2X1_LVT U155 ( .A1(A[26]), .A2(n181), .Y(n179) );
  HADDX1_LVT U156 ( .A0(A[26]), .B0(n181), .SO(SUM[26]) );
  AND3X1_LVT U157 ( .A1(A[24]), .A2(A[25]), .A3(n159), .Y(n181) );
  HADDX1_LVT U158 ( .A0(n182), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U159 ( .A1(n159), .A2(A[24]), .Y(n182) );
  AO22X1_LVT U160 ( .A1(A[24]), .A2(n183), .A3(n165), .A4(n159), .Y(SUM[24])
         );
  NAND3X0_LVT U161 ( .A1(A[23]), .A2(A[22]), .A3(n184), .Y(n183) );
  HADDX1_LVT U162 ( .A0(n185), .B0(A[23]), .SO(SUM[23]) );
  AND2X1_LVT U163 ( .A1(n184), .A2(A[22]), .Y(n185) );
  HADDX1_LVT U164 ( .A0(A[22]), .B0(n184), .SO(SUM[22]) );
  AND3X1_LVT U165 ( .A1(A[20]), .A2(A[21]), .A3(n160), .Y(n184) );
  HADDX1_LVT U166 ( .A0(n186), .B0(A[21]), .SO(SUM[21]) );
  AND2X1_LVT U167 ( .A1(n160), .A2(A[20]), .Y(n186) );
  AO22X1_LVT U168 ( .A1(A[20]), .A2(n187), .A3(n166), .A4(n160), .Y(SUM[20])
         );
  NAND2X0_LVT U169 ( .A1(n188), .A2(n161), .Y(n187) );
  AND4X1_LVT U170 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n188)
         );
  HADDX1_LVT U171 ( .A0(A[19]), .B0(n189), .SO(SUM[19]) );
  AND4X1_LVT U172 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n161), .Y(n189) );
  HADDX1_LVT U173 ( .A0(A[18]), .B0(n190), .SO(SUM[18]) );
  AND3X1_LVT U174 ( .A1(A[16]), .A2(A[17]), .A3(n161), .Y(n190) );
  HADDX1_LVT U175 ( .A0(n191), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U176 ( .A1(n161), .A2(A[16]), .Y(n191) );
  AO22X1_LVT U177 ( .A1(A[16]), .A2(n192), .A3(n167), .A4(n161), .Y(SUM[16])
         );
  NAND3X0_LVT U178 ( .A1(A[14]), .A2(A[15]), .A3(n193), .Y(n192) );
  HADDX1_LVT U179 ( .A0(A[15]), .B0(n194), .SO(SUM[15]) );
  AND4X1_LVT U180 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n162), .Y(n194) );
  HADDX1_LVT U181 ( .A0(A[14]), .B0(n193), .SO(SUM[14]) );
  AND3X1_LVT U182 ( .A1(A[12]), .A2(A[13]), .A3(n162), .Y(n193) );
  HADDX1_LVT U183 ( .A0(n195), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U184 ( .A1(n162), .A2(A[12]), .Y(n195) );
  AO22X1_LVT U185 ( .A1(A[12]), .A2(n196), .A3(n168), .A4(n162), .Y(SUM[12])
         );
  NAND2X0_LVT U186 ( .A1(n163), .A2(n197), .Y(n196) );
  AND4X1_LVT U187 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n197) );
  HADDX1_LVT U188 ( .A0(A[11]), .B0(n198), .SO(SUM[11]) );
  AND4X1_LVT U189 ( .A1(n163), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n198) );
  HADDX1_LVT U190 ( .A0(A[10]), .B0(n199), .SO(SUM[10]) );
  AND3X1_LVT U191 ( .A1(n163), .A2(A[9]), .A3(A[8]), .Y(n199) );
  NAND3X0_LVT U192 ( .A1(A[6]), .A2(A[7]), .A3(n174), .Y(n172) );
  AND3X1_LVT U193 ( .A1(A[4]), .A2(A[5]), .A3(n164), .Y(n174) );
  NAND3X0_LVT U194 ( .A1(n93), .A2(A[2]), .A3(A[3]), .Y(n176) );
endmodule


module CSRFile_DW01_inc_J38_8 ( A, SUM );
  input [57:0] A;
  output [57:0] SUM;
  wire   n203, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  HADDX1_LVT U259 ( .A0(A[1]), .B0(A[0]), .C1(n203), .SO(SUM[1]) );
  INVX0_LVT U264 ( .A(A[32]), .Y(n325) );
  AO22X1_LVT U265 ( .A1(A[32]), .A2(n383), .A3(n325), .A4(n334), .Y(SUM[32])
         );
  INVX0_LVT U266 ( .A(A[44]), .Y(n326) );
  AO22X1_LVT U267 ( .A1(A[44]), .A2(n367), .A3(n326), .A4(n331), .Y(SUM[44])
         );
  INVX0_LVT U268 ( .A(A[52]), .Y(n327) );
  AO22X1_LVT U269 ( .A1(A[52]), .A2(n355), .A3(n327), .A4(n329), .Y(SUM[52])
         );
  INVX0_LVT U270 ( .A(A[48]), .Y(n328) );
  AO22X1_LVT U271 ( .A1(A[48]), .A2(n361), .A3(n328), .A4(n330), .Y(SUM[48])
         );
  INVX1_LVT U272 ( .A(A[24]), .Y(n335) );
  INVX1_LVT U273 ( .A(A[8]), .Y(n341) );
  INVX1_LVT U274 ( .A(A[4]), .Y(n343) );
  INVX1_LVT U275 ( .A(A[12]), .Y(n339) );
  INVX1_LVT U276 ( .A(A[16]), .Y(n337) );
  INVX0_LVT U277 ( .A(A[40]), .Y(n332) );
  INVX1_LVT U278 ( .A(n383), .Y(n334) );
  INVX1_LVT U279 ( .A(n393), .Y(n336) );
  INVX1_LVT U280 ( .A(n404), .Y(n338) );
  INVX1_LVT U281 ( .A(n355), .Y(n329) );
  INVX1_LVT U282 ( .A(n361), .Y(n330) );
  INVX1_LVT U283 ( .A(n367), .Y(n331) );
  INVX1_LVT U284 ( .A(n371), .Y(n333) );
  INVX1_LVT U285 ( .A(n408), .Y(n340) );
  INVX1_LVT U286 ( .A(n346), .Y(n342) );
  INVX1_LVT U287 ( .A(n359), .Y(n344) );
  HADDX1_LVT U288 ( .A0(n345), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U289 ( .A1(A[8]), .A2(n342), .Y(n345) );
  AO22X1_LVT U290 ( .A1(n342), .A2(n341), .A3(n346), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U291 ( .A0(A[7]), .B0(n347), .SO(SUM[7]) );
  AND2X1_LVT U292 ( .A1(A[6]), .A2(n348), .Y(n347) );
  HADDX1_LVT U293 ( .A0(A[6]), .B0(n348), .SO(SUM[6]) );
  HADDX1_LVT U294 ( .A0(n349), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U295 ( .A1(n344), .A2(A[4]), .Y(n349) );
  HADDX1_LVT U296 ( .A0(A[57]), .B0(n350), .SO(SUM[57]) );
  AND4X1_LVT U297 ( .A1(A[55]), .A2(A[54]), .A3(n351), .A4(A[56]), .Y(n350) );
  HADDX1_LVT U298 ( .A0(n352), .B0(A[56]), .SO(SUM[56]) );
  AND3X1_LVT U299 ( .A1(A[55]), .A2(A[54]), .A3(n351), .Y(n352) );
  HADDX1_LVT U300 ( .A0(n353), .B0(A[55]), .SO(SUM[55]) );
  AND2X1_LVT U301 ( .A1(n351), .A2(A[54]), .Y(n353) );
  HADDX1_LVT U302 ( .A0(A[54]), .B0(n351), .SO(SUM[54]) );
  AND3X1_LVT U303 ( .A1(A[52]), .A2(A[53]), .A3(n329), .Y(n351) );
  HADDX1_LVT U304 ( .A0(n354), .B0(A[53]), .SO(SUM[53]) );
  AND2X1_LVT U305 ( .A1(n329), .A2(A[52]), .Y(n354) );
  NAND2X0_LVT U306 ( .A1(n356), .A2(n330), .Y(n355) );
  AND4X1_LVT U307 ( .A1(A[48]), .A2(A[49]), .A3(A[51]), .A4(A[50]), .Y(n356)
         );
  HADDX1_LVT U308 ( .A0(A[51]), .B0(n357), .SO(SUM[51]) );
  AND4X1_LVT U309 ( .A1(A[48]), .A2(A[49]), .A3(A[50]), .A4(n330), .Y(n357) );
  HADDX1_LVT U310 ( .A0(A[50]), .B0(n358), .SO(SUM[50]) );
  AND3X1_LVT U311 ( .A1(A[48]), .A2(A[49]), .A3(n330), .Y(n358) );
  AO22X1_LVT U312 ( .A1(A[4]), .A2(n359), .A3(n343), .A4(n344), .Y(SUM[4]) );
  HADDX1_LVT U313 ( .A0(n360), .B0(A[49]), .SO(SUM[49]) );
  AND2X1_LVT U314 ( .A1(n330), .A2(A[48]), .Y(n360) );
  NAND3X0_LVT U315 ( .A1(A[47]), .A2(A[46]), .A3(n362), .Y(n361) );
  AND4X1_LVT U316 ( .A1(A[44]), .A2(A[45]), .A3(n363), .A4(n333), .Y(n362) );
  HADDX1_LVT U317 ( .A0(A[47]), .B0(n364), .SO(SUM[47]) );
  AND4X1_LVT U318 ( .A1(A[46]), .A2(A[44]), .A3(A[45]), .A4(n331), .Y(n364) );
  HADDX1_LVT U319 ( .A0(A[46]), .B0(n365), .SO(SUM[46]) );
  AND3X1_LVT U320 ( .A1(A[44]), .A2(A[45]), .A3(n331), .Y(n365) );
  HADDX1_LVT U321 ( .A0(n366), .B0(A[45]), .SO(SUM[45]) );
  AND2X1_LVT U322 ( .A1(n331), .A2(A[44]), .Y(n366) );
  NAND2X0_LVT U323 ( .A1(n363), .A2(n333), .Y(n367) );
  AND4X1_LVT U324 ( .A1(A[40]), .A2(A[41]), .A3(A[43]), .A4(A[42]), .Y(n363)
         );
  HADDX1_LVT U325 ( .A0(A[43]), .B0(n368), .SO(SUM[43]) );
  AND4X1_LVT U326 ( .A1(A[40]), .A2(A[41]), .A3(A[42]), .A4(n333), .Y(n368) );
  HADDX1_LVT U327 ( .A0(A[42]), .B0(n369), .SO(SUM[42]) );
  AND3X1_LVT U328 ( .A1(A[40]), .A2(A[41]), .A3(n333), .Y(n369) );
  HADDX1_LVT U329 ( .A0(n370), .B0(A[41]), .SO(SUM[41]) );
  AND2X1_LVT U330 ( .A1(n333), .A2(A[40]), .Y(n370) );
  AO22X1_LVT U331 ( .A1(A[40]), .A2(n371), .A3(n332), .A4(n333), .Y(SUM[40])
         );
  NAND2X0_LVT U332 ( .A1(n334), .A2(n372), .Y(n371) );
  AND4X1_LVT U333 ( .A1(A[38]), .A2(A[39]), .A3(n373), .A4(n374), .Y(n372) );
  HADDX1_LVT U334 ( .A0(A[3]), .B0(n375), .SO(SUM[3]) );
  AND2X1_LVT U335 ( .A1(n203), .A2(A[2]), .Y(n375) );
  HADDX1_LVT U336 ( .A0(A[39]), .B0(n376), .SO(SUM[39]) );
  AND4X1_LVT U337 ( .A1(n334), .A2(A[38]), .A3(n373), .A4(n374), .Y(n376) );
  HADDX1_LVT U338 ( .A0(A[38]), .B0(n377), .SO(SUM[38]) );
  AND3X1_LVT U339 ( .A1(n334), .A2(n373), .A3(n374), .Y(n377) );
  AND2X1_LVT U340 ( .A1(A[36]), .A2(A[37]), .Y(n373) );
  HADDX1_LVT U341 ( .A0(n378), .B0(A[37]), .SO(SUM[37]) );
  AND3X1_LVT U342 ( .A1(A[36]), .A2(n334), .A3(n374), .Y(n378) );
  HADDX1_LVT U343 ( .A0(A[36]), .B0(n379), .SO(SUM[36]) );
  AND2X1_LVT U344 ( .A1(n334), .A2(n374), .Y(n379) );
  AND4X1_LVT U345 ( .A1(A[32]), .A2(A[33]), .A3(A[35]), .A4(A[34]), .Y(n374)
         );
  HADDX1_LVT U346 ( .A0(A[35]), .B0(n380), .SO(SUM[35]) );
  AND4X1_LVT U347 ( .A1(n334), .A2(A[32]), .A3(A[33]), .A4(A[34]), .Y(n380) );
  HADDX1_LVT U348 ( .A0(A[34]), .B0(n381), .SO(SUM[34]) );
  AND3X1_LVT U349 ( .A1(n334), .A2(A[32]), .A3(A[33]), .Y(n381) );
  HADDX1_LVT U350 ( .A0(n382), .B0(A[33]), .SO(SUM[33]) );
  AND2X1_LVT U351 ( .A1(A[32]), .A2(n334), .Y(n382) );
  NAND4X0_LVT U352 ( .A1(A[31]), .A2(A[30]), .A3(n384), .A4(n385), .Y(n383) );
  HADDX1_LVT U353 ( .A0(A[31]), .B0(n386), .SO(SUM[31]) );
  AND4X1_LVT U354 ( .A1(n387), .A2(A[30]), .A3(n384), .A4(n336), .Y(n386) );
  HADDX1_LVT U355 ( .A0(A[30]), .B0(n388), .SO(SUM[30]) );
  AND3X1_LVT U356 ( .A1(n387), .A2(n384), .A3(n336), .Y(n388) );
  AND2X1_LVT U357 ( .A1(A[28]), .A2(A[29]), .Y(n384) );
  HADDX1_LVT U358 ( .A0(n203), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U359 ( .A0(n389), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U360 ( .A1(A[28]), .A2(n387), .A3(n336), .Y(n389) );
  HADDX1_LVT U361 ( .A0(A[28]), .B0(n385), .SO(SUM[28]) );
  AND2X1_LVT U362 ( .A1(n387), .A2(n336), .Y(n385) );
  AND4X1_LVT U363 ( .A1(A[24]), .A2(A[25]), .A3(A[27]), .A4(A[26]), .Y(n387)
         );
  HADDX1_LVT U364 ( .A0(A[27]), .B0(n390), .SO(SUM[27]) );
  AND4X1_LVT U365 ( .A1(A[24]), .A2(A[25]), .A3(A[26]), .A4(n336), .Y(n390) );
  HADDX1_LVT U366 ( .A0(A[26]), .B0(n391), .SO(SUM[26]) );
  AND3X1_LVT U367 ( .A1(A[24]), .A2(A[25]), .A3(n336), .Y(n391) );
  HADDX1_LVT U368 ( .A0(n392), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U369 ( .A1(n336), .A2(A[24]), .Y(n392) );
  AO22X1_LVT U370 ( .A1(A[24]), .A2(n393), .A3(n335), .A4(n336), .Y(SUM[24])
         );
  NAND2X0_LVT U371 ( .A1(n394), .A2(n338), .Y(n393) );
  AND4X1_LVT U372 ( .A1(A[22]), .A2(A[23]), .A3(n395), .A4(n396), .Y(n394) );
  HADDX1_LVT U373 ( .A0(A[23]), .B0(n397), .SO(SUM[23]) );
  AND4X1_LVT U374 ( .A1(A[22]), .A2(n395), .A3(n396), .A4(n338), .Y(n397) );
  HADDX1_LVT U375 ( .A0(A[22]), .B0(n398), .SO(SUM[22]) );
  AND3X1_LVT U376 ( .A1(n395), .A2(n396), .A3(n338), .Y(n398) );
  AND2X1_LVT U377 ( .A1(A[20]), .A2(A[21]), .Y(n395) );
  HADDX1_LVT U378 ( .A0(n399), .B0(A[21]), .SO(SUM[21]) );
  AND3X1_LVT U379 ( .A1(n396), .A2(A[20]), .A3(n338), .Y(n399) );
  HADDX1_LVT U380 ( .A0(A[20]), .B0(n400), .SO(SUM[20]) );
  AND2X1_LVT U381 ( .A1(n396), .A2(n338), .Y(n400) );
  AND4X1_LVT U382 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n396)
         );
  HADDX1_LVT U383 ( .A0(A[19]), .B0(n401), .SO(SUM[19]) );
  AND4X1_LVT U384 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n338), .Y(n401) );
  HADDX1_LVT U385 ( .A0(A[18]), .B0(n402), .SO(SUM[18]) );
  AND3X1_LVT U386 ( .A1(A[16]), .A2(A[17]), .A3(n338), .Y(n402) );
  HADDX1_LVT U387 ( .A0(n403), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U388 ( .A1(n338), .A2(A[16]), .Y(n403) );
  AO22X1_LVT U389 ( .A1(A[16]), .A2(n404), .A3(n337), .A4(n338), .Y(SUM[16])
         );
  NAND3X0_LVT U390 ( .A1(A[14]), .A2(A[15]), .A3(n405), .Y(n404) );
  HADDX1_LVT U391 ( .A0(A[15]), .B0(n406), .SO(SUM[15]) );
  AND4X1_LVT U392 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n340), .Y(n406) );
  HADDX1_LVT U393 ( .A0(A[14]), .B0(n405), .SO(SUM[14]) );
  AND3X1_LVT U394 ( .A1(A[12]), .A2(A[13]), .A3(n340), .Y(n405) );
  HADDX1_LVT U395 ( .A0(n407), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U396 ( .A1(n340), .A2(A[12]), .Y(n407) );
  AO22X1_LVT U397 ( .A1(A[12]), .A2(n408), .A3(n339), .A4(n340), .Y(SUM[12])
         );
  NAND2X0_LVT U398 ( .A1(n342), .A2(n409), .Y(n408) );
  AND4X1_LVT U399 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n409) );
  HADDX1_LVT U400 ( .A0(A[11]), .B0(n410), .SO(SUM[11]) );
  AND4X1_LVT U401 ( .A1(n342), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n410) );
  HADDX1_LVT U402 ( .A0(A[10]), .B0(n411), .SO(SUM[10]) );
  AND3X1_LVT U403 ( .A1(n342), .A2(A[9]), .A3(A[8]), .Y(n411) );
  NAND3X0_LVT U404 ( .A1(A[6]), .A2(A[7]), .A3(n348), .Y(n346) );
  AND3X1_LVT U405 ( .A1(A[4]), .A2(A[5]), .A3(n344), .Y(n348) );
  NAND3X0_LVT U406 ( .A1(n203), .A2(A[2]), .A3(A[3]), .Y(n359) );
endmodule


module CSRFile_DW01_inc_J38_9 ( A, SUM );
  input [57:0] A;
  output [57:0] SUM;
  wire   n203, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  HADDX1_LVT U259 ( .A0(A[1]), .B0(A[0]), .C1(n203), .SO(SUM[1]) );
  INVX0_LVT U264 ( .A(A[52]), .Y(n325) );
  AO22X1_LVT U265 ( .A1(A[52]), .A2(n355), .A3(n325), .A4(n328), .Y(SUM[52])
         );
  INVX0_LVT U266 ( .A(A[44]), .Y(n326) );
  AO22X1_LVT U267 ( .A1(A[44]), .A2(n367), .A3(n326), .A4(n331), .Y(SUM[44])
         );
  INVX0_LVT U268 ( .A(A[32]), .Y(n327) );
  AO22X1_LVT U269 ( .A1(A[32]), .A2(n383), .A3(n327), .A4(n334), .Y(SUM[32])
         );
  INVX0_LVT U270 ( .A(A[24]), .Y(n335) );
  INVX0_LVT U271 ( .A(A[8]), .Y(n341) );
  INVX0_LVT U272 ( .A(A[48]), .Y(n329) );
  INVX0_LVT U273 ( .A(A[40]), .Y(n332) );
  INVX1_LVT U274 ( .A(n383), .Y(n334) );
  INVX1_LVT U275 ( .A(n393), .Y(n336) );
  INVX1_LVT U276 ( .A(n404), .Y(n338) );
  INVX1_LVT U277 ( .A(n355), .Y(n328) );
  INVX1_LVT U278 ( .A(n361), .Y(n330) );
  INVX1_LVT U279 ( .A(n367), .Y(n331) );
  INVX1_LVT U280 ( .A(n371), .Y(n333) );
  INVX1_LVT U281 ( .A(A[16]), .Y(n337) );
  INVX1_LVT U282 ( .A(A[12]), .Y(n339) );
  INVX1_LVT U283 ( .A(n408), .Y(n340) );
  INVX1_LVT U284 ( .A(n346), .Y(n342) );
  INVX1_LVT U285 ( .A(A[4]), .Y(n343) );
  INVX1_LVT U286 ( .A(n359), .Y(n344) );
  HADDX1_LVT U287 ( .A0(n345), .B0(A[9]), .SO(SUM[9]) );
  AND2X1_LVT U288 ( .A1(A[8]), .A2(n342), .Y(n345) );
  AO22X1_LVT U289 ( .A1(n342), .A2(n341), .A3(n346), .A4(A[8]), .Y(SUM[8]) );
  HADDX1_LVT U290 ( .A0(A[7]), .B0(n347), .SO(SUM[7]) );
  AND2X1_LVT U291 ( .A1(A[6]), .A2(n348), .Y(n347) );
  HADDX1_LVT U292 ( .A0(A[6]), .B0(n348), .SO(SUM[6]) );
  HADDX1_LVT U293 ( .A0(n349), .B0(A[5]), .SO(SUM[5]) );
  AND2X1_LVT U294 ( .A1(n344), .A2(A[4]), .Y(n349) );
  HADDX1_LVT U295 ( .A0(A[57]), .B0(n350), .SO(SUM[57]) );
  AND4X1_LVT U296 ( .A1(A[55]), .A2(A[54]), .A3(n351), .A4(A[56]), .Y(n350) );
  HADDX1_LVT U297 ( .A0(n352), .B0(A[56]), .SO(SUM[56]) );
  AND3X1_LVT U298 ( .A1(A[55]), .A2(A[54]), .A3(n351), .Y(n352) );
  HADDX1_LVT U299 ( .A0(n353), .B0(A[55]), .SO(SUM[55]) );
  AND2X1_LVT U300 ( .A1(n351), .A2(A[54]), .Y(n353) );
  HADDX1_LVT U301 ( .A0(A[54]), .B0(n351), .SO(SUM[54]) );
  AND3X1_LVT U302 ( .A1(A[52]), .A2(A[53]), .A3(n328), .Y(n351) );
  HADDX1_LVT U303 ( .A0(n354), .B0(A[53]), .SO(SUM[53]) );
  AND2X1_LVT U304 ( .A1(n328), .A2(A[52]), .Y(n354) );
  NAND2X0_LVT U305 ( .A1(n356), .A2(n330), .Y(n355) );
  AND4X1_LVT U306 ( .A1(A[48]), .A2(A[49]), .A3(A[51]), .A4(A[50]), .Y(n356)
         );
  HADDX1_LVT U307 ( .A0(A[51]), .B0(n357), .SO(SUM[51]) );
  AND4X1_LVT U308 ( .A1(A[48]), .A2(A[49]), .A3(A[50]), .A4(n330), .Y(n357) );
  HADDX1_LVT U309 ( .A0(A[50]), .B0(n358), .SO(SUM[50]) );
  AND3X1_LVT U310 ( .A1(A[48]), .A2(A[49]), .A3(n330), .Y(n358) );
  AO22X1_LVT U311 ( .A1(A[4]), .A2(n359), .A3(n343), .A4(n344), .Y(SUM[4]) );
  HADDX1_LVT U312 ( .A0(n360), .B0(A[49]), .SO(SUM[49]) );
  AND2X1_LVT U313 ( .A1(n330), .A2(A[48]), .Y(n360) );
  AO22X1_LVT U314 ( .A1(A[48]), .A2(n361), .A3(n329), .A4(n330), .Y(SUM[48])
         );
  NAND3X0_LVT U315 ( .A1(A[47]), .A2(A[46]), .A3(n362), .Y(n361) );
  AND4X1_LVT U316 ( .A1(A[44]), .A2(A[45]), .A3(n363), .A4(n333), .Y(n362) );
  HADDX1_LVT U317 ( .A0(A[47]), .B0(n364), .SO(SUM[47]) );
  AND4X1_LVT U318 ( .A1(A[46]), .A2(A[44]), .A3(A[45]), .A4(n331), .Y(n364) );
  HADDX1_LVT U319 ( .A0(A[46]), .B0(n365), .SO(SUM[46]) );
  AND3X1_LVT U320 ( .A1(A[44]), .A2(A[45]), .A3(n331), .Y(n365) );
  HADDX1_LVT U321 ( .A0(n366), .B0(A[45]), .SO(SUM[45]) );
  AND2X1_LVT U322 ( .A1(n331), .A2(A[44]), .Y(n366) );
  NAND2X0_LVT U323 ( .A1(n363), .A2(n333), .Y(n367) );
  AND4X1_LVT U324 ( .A1(A[40]), .A2(A[41]), .A3(A[43]), .A4(A[42]), .Y(n363)
         );
  HADDX1_LVT U325 ( .A0(A[43]), .B0(n368), .SO(SUM[43]) );
  AND4X1_LVT U326 ( .A1(A[40]), .A2(A[41]), .A3(A[42]), .A4(n333), .Y(n368) );
  HADDX1_LVT U327 ( .A0(A[42]), .B0(n369), .SO(SUM[42]) );
  AND3X1_LVT U328 ( .A1(A[40]), .A2(A[41]), .A3(n333), .Y(n369) );
  HADDX1_LVT U329 ( .A0(n370), .B0(A[41]), .SO(SUM[41]) );
  AND2X1_LVT U330 ( .A1(n333), .A2(A[40]), .Y(n370) );
  AO22X1_LVT U331 ( .A1(A[40]), .A2(n371), .A3(n332), .A4(n333), .Y(SUM[40])
         );
  NAND2X0_LVT U332 ( .A1(n334), .A2(n372), .Y(n371) );
  AND4X1_LVT U333 ( .A1(A[38]), .A2(A[39]), .A3(n373), .A4(n374), .Y(n372) );
  HADDX1_LVT U334 ( .A0(A[3]), .B0(n375), .SO(SUM[3]) );
  AND2X1_LVT U335 ( .A1(n203), .A2(A[2]), .Y(n375) );
  HADDX1_LVT U336 ( .A0(A[39]), .B0(n376), .SO(SUM[39]) );
  AND4X1_LVT U337 ( .A1(n334), .A2(A[38]), .A3(n373), .A4(n374), .Y(n376) );
  HADDX1_LVT U338 ( .A0(A[38]), .B0(n377), .SO(SUM[38]) );
  AND3X1_LVT U339 ( .A1(n334), .A2(n373), .A3(n374), .Y(n377) );
  AND2X1_LVT U340 ( .A1(A[36]), .A2(A[37]), .Y(n373) );
  HADDX1_LVT U341 ( .A0(n378), .B0(A[37]), .SO(SUM[37]) );
  AND3X1_LVT U342 ( .A1(A[36]), .A2(n334), .A3(n374), .Y(n378) );
  HADDX1_LVT U343 ( .A0(A[36]), .B0(n379), .SO(SUM[36]) );
  AND2X1_LVT U344 ( .A1(n334), .A2(n374), .Y(n379) );
  AND4X1_LVT U345 ( .A1(A[32]), .A2(A[33]), .A3(A[35]), .A4(A[34]), .Y(n374)
         );
  HADDX1_LVT U346 ( .A0(A[35]), .B0(n380), .SO(SUM[35]) );
  AND4X1_LVT U347 ( .A1(n334), .A2(A[32]), .A3(A[33]), .A4(A[34]), .Y(n380) );
  HADDX1_LVT U348 ( .A0(A[34]), .B0(n381), .SO(SUM[34]) );
  AND3X1_LVT U349 ( .A1(n334), .A2(A[32]), .A3(A[33]), .Y(n381) );
  HADDX1_LVT U350 ( .A0(n382), .B0(A[33]), .SO(SUM[33]) );
  AND2X1_LVT U351 ( .A1(A[32]), .A2(n334), .Y(n382) );
  NAND4X0_LVT U352 ( .A1(A[31]), .A2(A[30]), .A3(n384), .A4(n385), .Y(n383) );
  HADDX1_LVT U353 ( .A0(A[31]), .B0(n386), .SO(SUM[31]) );
  AND4X1_LVT U354 ( .A1(n387), .A2(A[30]), .A3(n384), .A4(n336), .Y(n386) );
  HADDX1_LVT U355 ( .A0(A[30]), .B0(n388), .SO(SUM[30]) );
  AND3X1_LVT U356 ( .A1(n387), .A2(n384), .A3(n336), .Y(n388) );
  AND2X1_LVT U357 ( .A1(A[28]), .A2(A[29]), .Y(n384) );
  HADDX1_LVT U358 ( .A0(n203), .B0(A[2]), .SO(SUM[2]) );
  HADDX1_LVT U359 ( .A0(n389), .B0(A[29]), .SO(SUM[29]) );
  AND3X1_LVT U360 ( .A1(A[28]), .A2(n387), .A3(n336), .Y(n389) );
  HADDX1_LVT U361 ( .A0(A[28]), .B0(n385), .SO(SUM[28]) );
  AND2X1_LVT U362 ( .A1(n387), .A2(n336), .Y(n385) );
  AND4X1_LVT U363 ( .A1(A[24]), .A2(A[25]), .A3(A[27]), .A4(A[26]), .Y(n387)
         );
  HADDX1_LVT U364 ( .A0(A[27]), .B0(n390), .SO(SUM[27]) );
  AND4X1_LVT U365 ( .A1(A[24]), .A2(A[25]), .A3(A[26]), .A4(n336), .Y(n390) );
  HADDX1_LVT U366 ( .A0(A[26]), .B0(n391), .SO(SUM[26]) );
  AND3X1_LVT U367 ( .A1(A[24]), .A2(A[25]), .A3(n336), .Y(n391) );
  HADDX1_LVT U368 ( .A0(n392), .B0(A[25]), .SO(SUM[25]) );
  AND2X1_LVT U369 ( .A1(n336), .A2(A[24]), .Y(n392) );
  AO22X1_LVT U370 ( .A1(A[24]), .A2(n393), .A3(n335), .A4(n336), .Y(SUM[24])
         );
  NAND2X0_LVT U371 ( .A1(n394), .A2(n338), .Y(n393) );
  AND4X1_LVT U372 ( .A1(A[22]), .A2(A[23]), .A3(n395), .A4(n396), .Y(n394) );
  HADDX1_LVT U373 ( .A0(A[23]), .B0(n397), .SO(SUM[23]) );
  AND4X1_LVT U374 ( .A1(A[22]), .A2(n395), .A3(n396), .A4(n338), .Y(n397) );
  HADDX1_LVT U375 ( .A0(A[22]), .B0(n398), .SO(SUM[22]) );
  AND3X1_LVT U376 ( .A1(n395), .A2(n396), .A3(n338), .Y(n398) );
  AND2X1_LVT U377 ( .A1(A[20]), .A2(A[21]), .Y(n395) );
  HADDX1_LVT U378 ( .A0(n399), .B0(A[21]), .SO(SUM[21]) );
  AND3X1_LVT U379 ( .A1(n396), .A2(A[20]), .A3(n338), .Y(n399) );
  HADDX1_LVT U380 ( .A0(A[20]), .B0(n400), .SO(SUM[20]) );
  AND2X1_LVT U381 ( .A1(n396), .A2(n338), .Y(n400) );
  AND4X1_LVT U382 ( .A1(A[16]), .A2(A[17]), .A3(A[19]), .A4(A[18]), .Y(n396)
         );
  HADDX1_LVT U383 ( .A0(A[19]), .B0(n401), .SO(SUM[19]) );
  AND4X1_LVT U384 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n338), .Y(n401) );
  HADDX1_LVT U385 ( .A0(A[18]), .B0(n402), .SO(SUM[18]) );
  AND3X1_LVT U386 ( .A1(A[16]), .A2(A[17]), .A3(n338), .Y(n402) );
  HADDX1_LVT U387 ( .A0(n403), .B0(A[17]), .SO(SUM[17]) );
  AND2X1_LVT U388 ( .A1(n338), .A2(A[16]), .Y(n403) );
  AO22X1_LVT U389 ( .A1(A[16]), .A2(n404), .A3(n337), .A4(n338), .Y(SUM[16])
         );
  NAND3X0_LVT U390 ( .A1(A[14]), .A2(A[15]), .A3(n405), .Y(n404) );
  HADDX1_LVT U391 ( .A0(A[15]), .B0(n406), .SO(SUM[15]) );
  AND4X1_LVT U392 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n340), .Y(n406) );
  HADDX1_LVT U393 ( .A0(A[14]), .B0(n405), .SO(SUM[14]) );
  AND3X1_LVT U394 ( .A1(A[12]), .A2(A[13]), .A3(n340), .Y(n405) );
  HADDX1_LVT U395 ( .A0(n407), .B0(A[13]), .SO(SUM[13]) );
  AND2X1_LVT U396 ( .A1(n340), .A2(A[12]), .Y(n407) );
  AO22X1_LVT U397 ( .A1(A[12]), .A2(n408), .A3(n339), .A4(n340), .Y(SUM[12])
         );
  NAND2X0_LVT U398 ( .A1(n342), .A2(n409), .Y(n408) );
  AND4X1_LVT U399 ( .A1(A[9]), .A2(A[8]), .A3(A[11]), .A4(A[10]), .Y(n409) );
  HADDX1_LVT U400 ( .A0(A[11]), .B0(n410), .SO(SUM[11]) );
  AND4X1_LVT U401 ( .A1(n342), .A2(A[9]), .A3(A[8]), .A4(A[10]), .Y(n410) );
  HADDX1_LVT U402 ( .A0(A[10]), .B0(n411), .SO(SUM[10]) );
  AND3X1_LVT U403 ( .A1(n342), .A2(A[9]), .A3(A[8]), .Y(n411) );
  NAND3X0_LVT U404 ( .A1(A[6]), .A2(A[7]), .A3(n348), .Y(n346) );
  AND3X1_LVT U405 ( .A1(A[4]), .A2(A[5]), .A3(n344), .Y(n348) );
  NAND3X0_LVT U406 ( .A1(n203), .A2(A[2]), .A3(A[3]), .Y(n359) );
endmodule


module SNPS_CLOCK_GATE_HIGH_CSRFile_0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module CSRFile ( clock, reset, io_ungated_clock, io_interrupts_debug, 
        io_interrupts_mtip, io_interrupts_msip, io_interrupts_meip, 
        io_interrupts_seip, io_rw_addr, io_rw_cmd, io_rw_rdata, io_rw_wdata, 
        io_decode_0_csr, io_decode_0_fp_illegal, io_decode_0_fp_csr, 
        io_decode_0_read_illegal, io_decode_0_write_illegal, 
        io_decode_0_write_flush, io_decode_0_system_illegal, io_csr_stall, 
        io_eret, io_singleStep, io_status_cease, io_status_wfi, io_status_dprv, 
        io_status_prv, io_status_sd, io_status_zero2, io_status_sxl, 
        io_status_uxl, io_status_sd_rv32, io_status_zero1, io_status_tsr, 
        io_status_tw, io_status_tvm, io_status_mxr, io_status_sum, 
        io_status_mprv, io_status_xs, io_status_fs, io_status_mpp, 
        io_status_vs, io_status_spp, io_status_mpie, io_status_hpie, 
        io_status_spie, io_status_upie, io_status_mie, io_status_hie, 
        io_status_sie, io_status_uie, io_ptbr_mode, io_ptbr_ppn, io_evec, 
        io_exception, io_retire, io_cause, io_pc, io_tval, io_time, io_fcsr_rm, 
        io_fcsr_flags_valid, io_fcsr_flags_bits, io_interrupt, 
        io_interrupt_cause, io_bp_0_control_action, io_bp_0_control_tmatch, 
        io_bp_0_control_m, io_bp_0_control_s, io_bp_0_control_u, 
        io_bp_0_control_x, io_bp_0_control_w, io_bp_0_control_r, 
        io_bp_0_address, io_pmp_0_cfg_l, io_pmp_0_cfg_a, io_pmp_0_cfg_x, 
        io_pmp_0_cfg_w, io_pmp_0_cfg_r, io_pmp_0_addr, io_pmp_0_mask, 
        io_pmp_1_cfg_l, io_pmp_1_cfg_a, io_pmp_1_cfg_x, io_pmp_1_cfg_w, 
        io_pmp_1_cfg_r, io_pmp_1_addr, io_pmp_1_mask, io_pmp_2_cfg_l, 
        io_pmp_2_cfg_a, io_pmp_2_cfg_x, io_pmp_2_cfg_w, io_pmp_2_cfg_r, 
        io_pmp_2_addr, io_pmp_2_mask, io_pmp_3_cfg_l, io_pmp_3_cfg_a, 
        io_pmp_3_cfg_x, io_pmp_3_cfg_w, io_pmp_3_cfg_r, io_pmp_3_addr, 
        io_pmp_3_mask, io_pmp_4_cfg_l, io_pmp_4_cfg_a, io_pmp_4_cfg_x, 
        io_pmp_4_cfg_w, io_pmp_4_cfg_r, io_pmp_4_addr, io_pmp_4_mask, 
        io_pmp_5_cfg_l, io_pmp_5_cfg_a, io_pmp_5_cfg_x, io_pmp_5_cfg_w, 
        io_pmp_5_cfg_r, io_pmp_5_addr, io_pmp_5_mask, io_pmp_6_cfg_l, 
        io_pmp_6_cfg_a, io_pmp_6_cfg_x, io_pmp_6_cfg_w, io_pmp_6_cfg_r, 
        io_pmp_6_addr, io_pmp_6_mask, io_pmp_7_cfg_l, io_pmp_7_cfg_a, 
        io_pmp_7_cfg_x, io_pmp_7_cfg_w, io_pmp_7_cfg_r, io_pmp_7_addr, 
        io_pmp_7_mask, io_inst_0, io_trace_0_valid, io_trace_0_iaddr, 
        io_trace_0_insn, io_trace_0_exception, io_customCSRs_0_value, 
        io_status_debug_BAR, io_status_isa_31_, io_status_isa_30_, 
        io_status_isa_29_, io_status_isa_28_, io_status_isa_27_, 
        io_status_isa_26_, io_status_isa_25_, io_status_isa_24_, 
        io_status_isa_23_, io_status_isa_22_, io_status_isa_21_, 
        io_status_isa_20_, io_status_isa_19_, io_status_isa_18_, 
        io_status_isa_17_, io_status_isa_16_, io_status_isa_15_, 
        io_status_isa_14_, io_status_isa_13_, io_status_isa_12__BAR, 
        io_status_isa_11_, io_status_isa_10_, io_status_isa_9_, 
        io_status_isa_8_, io_status_isa_7_, io_status_isa_6_, io_status_isa_5_, 
        io_status_isa_4_, io_status_isa_3_, io_status_isa_2_, io_status_isa_1_, 
        io_status_isa_0__BAR );
  input [11:0] io_rw_addr;
  input [2:0] io_rw_cmd;
  output [63:0] io_rw_rdata;
  input [63:0] io_rw_wdata;
  input [11:0] io_decode_0_csr;
  output [1:0] io_status_dprv;
  output [1:0] io_status_prv;
  output [26:0] io_status_zero2;
  output [1:0] io_status_sxl;
  output [1:0] io_status_uxl;
  output [7:0] io_status_zero1;
  output [1:0] io_status_xs;
  output [1:0] io_status_fs;
  output [1:0] io_status_mpp;
  output [1:0] io_status_vs;
  output [3:0] io_ptbr_mode;
  output [43:0] io_ptbr_ppn;
  output [39:0] io_evec;
  input [63:0] io_cause;
  input [39:0] io_pc;
  input [39:0] io_tval;
  output [63:0] io_time;
  output [2:0] io_fcsr_rm;
  input [4:0] io_fcsr_flags_bits;
  output [63:0] io_interrupt_cause;
  output [1:0] io_bp_0_control_tmatch;
  output [38:0] io_bp_0_address;
  output [1:0] io_pmp_0_cfg_a;
  output [29:0] io_pmp_0_addr;
  output [31:0] io_pmp_0_mask;
  output [1:0] io_pmp_1_cfg_a;
  output [29:0] io_pmp_1_addr;
  output [31:0] io_pmp_1_mask;
  output [1:0] io_pmp_2_cfg_a;
  output [29:0] io_pmp_2_addr;
  output [31:0] io_pmp_2_mask;
  output [1:0] io_pmp_3_cfg_a;
  output [29:0] io_pmp_3_addr;
  output [31:0] io_pmp_3_mask;
  output [1:0] io_pmp_4_cfg_a;
  output [29:0] io_pmp_4_addr;
  output [31:0] io_pmp_4_mask;
  output [1:0] io_pmp_5_cfg_a;
  output [29:0] io_pmp_5_addr;
  output [31:0] io_pmp_5_mask;
  output [1:0] io_pmp_6_cfg_a;
  output [29:0] io_pmp_6_addr;
  output [31:0] io_pmp_6_mask;
  output [1:0] io_pmp_7_cfg_a;
  output [29:0] io_pmp_7_addr;
  output [31:0] io_pmp_7_mask;
  input [31:0] io_inst_0;
  output [39:0] io_trace_0_iaddr;
  output [31:0] io_trace_0_insn;
  output [63:0] io_customCSRs_0_value;
  input clock, reset, io_ungated_clock, io_interrupts_debug,
         io_interrupts_mtip, io_interrupts_msip, io_interrupts_meip,
         io_interrupts_seip, io_exception, io_retire, io_fcsr_flags_valid;
  output io_decode_0_fp_illegal, io_decode_0_fp_csr, io_decode_0_read_illegal,
         io_decode_0_write_illegal, io_decode_0_write_flush,
         io_decode_0_system_illegal, io_csr_stall, io_eret, io_singleStep,
         io_status_cease, io_status_wfi, io_status_sd, io_status_sd_rv32,
         io_status_tsr, io_status_tw, io_status_tvm, io_status_mxr,
         io_status_sum, io_status_mprv, io_status_spp, io_status_mpie,
         io_status_hpie, io_status_spie, io_status_upie, io_status_mie,
         io_status_hie, io_status_sie, io_status_uie, io_interrupt,
         io_bp_0_control_action, io_bp_0_control_m, io_bp_0_control_s,
         io_bp_0_control_u, io_bp_0_control_x, io_bp_0_control_w,
         io_bp_0_control_r, io_pmp_0_cfg_l, io_pmp_0_cfg_x, io_pmp_0_cfg_w,
         io_pmp_0_cfg_r, io_pmp_1_cfg_l, io_pmp_1_cfg_x, io_pmp_1_cfg_w,
         io_pmp_1_cfg_r, io_pmp_2_cfg_l, io_pmp_2_cfg_x, io_pmp_2_cfg_w,
         io_pmp_2_cfg_r, io_pmp_3_cfg_l, io_pmp_3_cfg_x, io_pmp_3_cfg_w,
         io_pmp_3_cfg_r, io_pmp_4_cfg_l, io_pmp_4_cfg_x, io_pmp_4_cfg_w,
         io_pmp_4_cfg_r, io_pmp_5_cfg_l, io_pmp_5_cfg_x, io_pmp_5_cfg_w,
         io_pmp_5_cfg_r, io_pmp_6_cfg_l, io_pmp_6_cfg_x, io_pmp_6_cfg_w,
         io_pmp_6_cfg_r, io_pmp_7_cfg_l, io_pmp_7_cfg_x, io_pmp_7_cfg_w,
         io_pmp_7_cfg_r, io_trace_0_valid, io_trace_0_exception,
         io_status_debug_BAR, io_status_isa_31_, io_status_isa_30_,
         io_status_isa_29_, io_status_isa_28_, io_status_isa_27_,
         io_status_isa_26_, io_status_isa_25_, io_status_isa_24_,
         io_status_isa_23_, io_status_isa_22_, io_status_isa_21_,
         io_status_isa_20_, io_status_isa_19_, io_status_isa_18_,
         io_status_isa_17_, io_status_isa_16_, io_status_isa_15_,
         io_status_isa_14_, io_status_isa_13_, io_status_isa_12__BAR,
         io_status_isa_11_, io_status_isa_10_, io_status_isa_9_,
         io_status_isa_8_, io_status_isa_7_, io_status_isa_6_,
         io_status_isa_5_, io_status_isa_4_, io_status_isa_3_,
         io_status_isa_2_, io_status_isa_1_, io_status_isa_0__BAR;
  wire   io_status_debug, n1918, n1919, n1920, n1921, io_status_isa_12_, n1922,
         n1923, io_status_isa_0_, n1924, n1925, n1926, n1927, n1928, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n_T_1155_3, read_mideleg_9_,
         read_mideleg_5, read_mideleg_1, read_medeleg_15, read_medeleg_13,
         read_medeleg_12, read_medeleg_8, read_medeleg_6, read_medeleg_0,
         n_T_61_5_, n_T_61_1, n_T_366_59_, n_T_389_2, n_T_389_1, n_T_389_0,
         n_T_3678_63_, n_T_3694_9_, N276, N290, N333, N334, N335, N360, N435,
         N438, N459, N460, N467, N469, N475, N479, N485, N487, N515, N518,
         N527, N531, N539, N542, N551, N556, N559, N568, N575, N580, N587,
         N592, N595, N604, N607, N609, N611, N613, N615, N617, N670, N880,
         N881, N882, N883, N884, N944, N992, N993, N994, N995, N996, N997,
         N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017,
         N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027,
         N1028, N1029, N1030, N1031, N1032, N1033, N1269, N1270, N1271, N1272,
         N1273, N1274, N1333, N1381, N1382, N1383, N1384, N1385, N1386, N1387,
         N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397,
         N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407,
         N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417,
         N1418, N1419, N1420, N1421, N1422, N1426, N1428, N1429, N1430, N1431,
         N1432, N1433, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503,
         N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513,
         N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523,
         N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533,
         N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543,
         N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553,
         N1554, N1558, N1567, N1577, N1579, N1582, N1622, N1691, N1692, N1693,
         N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1890, N1891, N1892,
         N1893, N1894, N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902,
         N1903, N1904, N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912,
         N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922,
         N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932,
         N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942,
         N1943, N1944, N1945, N1946, N1947, N1948, net34722, net34728,
         net34733, net34738, net34743, net34748, net34753, net34759, net34763,
         net34766, net34769, net34772, net34775, net34778, net34781, net34784,
         net34787, net34790, net34793, net34796, net34799, net34802, net34805,
         net34808, net34811, net34814, net34817, net34820, net34823, net34826,
         net34829, net34832, net34835, net34838, net34841, net34844, net34847,
         net34850, net34853, net34856, net34859, net34862, net34865, net34868,
         net34871, net34874, net34877, net34880, net34885, net34890, net34895,
         net34900, net34905, net34910, net34915, net34920, net34925, net34930,
         net34935, net34940, net34945, net34950, net34955, net34961, net34965,
         net34968, net34971, net34974, net34977, net34980, net34983, net34986,
         net34989, net34992, net34995, net34998, net35001, net35004, net35007,
         net35010, net35013, net35016, net35019, net35022, net35025, net35028,
         net35031, net35034, net35037, net35040, net35043, net35046, net35049,
         net35052, net35055, net35058, net35061, net35064, net35067, net35070,
         net35073, net35076, net35079, net35082, net35087, net35092, net35097,
         net35102, net35107, net35112, net35117, net35122, net35127, net35132,
         net35137, net35147, net35152, net35157, net35162, net35167, net35172,
         net35177, net35183, net35187, net35190, net35193, net35196, net35199,
         net35202, net35205, net35208, net35211, net35214, net35217, net35220,
         net35223, net35226, net35229, net35232, net35235, net35238, net35241,
         net35244, net35247, net35250, net35253, net35256, net35259, net35262,
         net35265, net35268, net35271, net35274, net35277, net35280, net35283,
         net35286, net35289, net35292, net35295, net35298, net35301, net35304,
         net35309, net35314, net35319, net35324, n51, n194, n199, n200, n658,
         n659, n860, n1041, n1062, n1346, n2155, n2156, n2157, n2160, n2161,
         n2162, n2163, n2165, n2166, n2167, n2168, n2169, n1, n2, n3, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n195, n196, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n258, n259, n260, n261, n262,
         n263, n264, n265, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n280, n281, n282, n283, n284, n285, n286,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1917, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10;
  wire   [1929:1930] n;
  wire   [1:0] n_T_1155;
  wire   [4:2] read_medeleg;
  wire   [2:0] read_mcounteren;
  wire   [2:0] read_scounteren;
  wire   [57:1] n_T_44;
  wire   [63:0] n_T_45;
  wire   [57:1] n_T_52;
  wire   [11:1] reg_mie;
  wire   [29:1] n_T_241;
  wire   [29:1] n_T_250;
  wire   [29:1] n_T_259;
  wire   [29:1] n_T_268;
  wire   [29:1] n_T_277;
  wire   [29:1] n_T_286;
  wire   [29:1] n_T_295;
  wire   [29:1] n_T_304;
  wire   [31:2] reg_mtvec;
  wire   [38:2] reg_stvec;
  wire   [39:1] reg_mepc;
  wire   [39:0] n_T_383;
  wire   [8:6] n_T_389;
  wire   [39:1] reg_dpc;
  wire   [4:0] read_fcsr;
  wire   [39:0] n_T_444;
  wire   [39:1] reg_sepc;
  wire   [63:0] wdata;
  wire   [63:0] reg_mscratch;
  wire   [63:0] reg_mcause;
  wire   [63:0] reg_dscratch;
  wire   [63:0] reg_sscratch;
  wire   [63:0] reg_scause;
  wire   [2:0] n_GEN_155;
  wire   [29:0] n_GEN_258;
  wire   [29:0] n_GEN_265;
  wire   [29:0] n_GEN_272;
  wire   [29:0] n_GEN_279;
  wire   [29:0] n_GEN_286;
  wire   [29:0] n_GEN_293;
  wire   [29:0] n_GEN_300;
  wire   [29:0] n_GEN_307;
  wire   [4:0] n_GEN_345;
  assign io_pmp_0_mask[2] = io_pmp_0_cfg_a[0];
  assign io_pmp_1_mask[2] = io_pmp_1_cfg_a[0];
  assign io_pmp_2_mask[2] = io_pmp_2_cfg_a[0];
  assign io_pmp_3_mask[2] = io_pmp_3_cfg_a[0];
  assign io_pmp_4_mask[2] = io_pmp_4_cfg_a[0];
  assign io_pmp_5_mask[2] = io_pmp_5_cfg_a[0];
  assign io_pmp_6_mask[2] = io_pmp_6_cfg_a[0];
  assign io_pmp_7_mask[2] = io_pmp_7_cfg_a[0];

  SNPS_CLOCK_GATE_HIGH_CSRFile_0 clk_gate_reg_bp_0_address_reg ( .CLK(n594), 
        .EN(n2163), .ENCLK(net34722), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_47 clk_gate_reg_mie_reg ( .CLK(n594), .EN(N670), 
        .ENCLK(net34728), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_46 clk_gate_reg_pmp_0_cfg_x_reg ( .CLK(n594), 
        .EN(N518), .ENCLK(net34733), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_45 clk_gate_reg_pmp_7_cfg_r_reg ( .CLK(n593), 
        .EN(N604), .ENCLK(net34738), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_44 clk_gate_reg_pmp_7_cfg_l_reg ( .CLK(n593), 
        .EN(N595), .ENCLK(net34743), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_43 clk_gate_reg_pmp_2_cfg_x_reg ( .CLK(n593), 
        .EN(N542), .ENCLK(net34748), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_42 clk_gate_reg_pmp_2_cfg_a_reg ( .CLK(n593), 
        .EN(N539), .ENCLK(net34753), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_41 clk_gate_reg_sepc_reg ( .CLK(n593), .EN(
        net34759), .ENCLK(net34880), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_40 clk_gate_reg_mcause_reg ( .CLK(n593), .EN(
        N880), .ENCLK(net34885), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_39 clk_gate__T_41_reg ( .CLK(n593), .EN(N1496), 
        .ENCLK(net34890), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_38 clk_gate_reg_mtval_reg ( .CLK(n593), .EN(
        N992), .ENCLK(net34895), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_37 clk_gate_reg_frm_reg ( .CLK(n593), .EN(n2166), .ENCLK(net34900), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_36 clk_gate_reg_pmp_0_cfg_a_reg ( .CLK(n593), 
        .EN(N515), .ENCLK(net34905), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_35 clk_gate_reg_pmp_4_cfg_l_reg ( .CLK(n593), 
        .EN(N559), .ENCLK(net34910), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_34 clk_gate_reg_satp_ppn_reg ( .CLK(n593), .EN(
        N1426), .ENCLK(net34915), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_33 clk_gate_reg_stvec_reg ( .CLK(n593), .EN(
        n2167), .ENCLK(net34920), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_32 clk_gate_reg_sscratch_reg ( .CLK(n593), .EN(
        N1422), .ENCLK(net34925), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_31 clk_gate_reg_stval_reg ( .CLK(n593), .EN(
        N1381), .ENCLK(net34930), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_30 clk_gate_reg_scause_reg ( .CLK(n593), .EN(
        N1269), .ENCLK(net34935), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_29 clk_gate_reg_scounteren_reg ( .CLK(n593), 
        .EN(n2168), .ENCLK(net34940), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_28 clk_gate_reg_mcounteren_reg ( .CLK(n593), 
        .EN(n2169), .ENCLK(net34945), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_27 clk_gate_reg_mtvec_reg ( .CLK(n593), .EN(
        n2165), .ENCLK(net34950), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_26 clk_gate_reg_mscratch_reg ( .CLK(n593), .EN(
        N1033), .ENCLK(net34955), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_25 clk_gate_reg_mepc_reg ( .CLK(n593), .EN(
        net34961), .ENCLK(net35082), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_24 clk_gate_reg_pmp_1_cfg_w_reg ( .CLK(n593), 
        .EN(N531), .ENCLK(net35087), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_23 clk_gate_reg_pmp_6_addr_reg ( .CLK(n592), 
        .EN(n504), .ENCLK(net35092), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_22 clk_gate_reg_pmp_5_cfg_r_reg ( .CLK(n592), 
        .EN(N580), .ENCLK(net35097), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_21 clk_gate_reg_pmp_6_cfg_a_reg ( .CLK(n592), 
        .EN(N587), .ENCLK(net35102), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_20 clk_gate_reg_pmp_6_cfg_r_reg ( .CLK(n592), 
        .EN(N592), .ENCLK(net35107), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_19 clk_gate_reg_pmp_5_cfg_a_reg ( .CLK(n592), 
        .EN(N575), .ENCLK(net35112), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_18 clk_gate_reg_pmp_4_cfg_r_reg ( .CLK(n592), 
        .EN(N568), .ENCLK(net35117), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_17 clk_gate_reg_pmp_3_cfg_r_reg ( .CLK(n592), 
        .EN(N556), .ENCLK(net35122), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_16 clk_gate_reg_pmp_3_cfg_a_reg ( .CLK(n592), 
        .EN(N551), .ENCLK(net35127), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_15 clk_gate_reg_pmp_1_cfg_a_reg ( .CLK(n592), 
        .EN(N527), .ENCLK(net35132), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_14 clk_gate_reg_misa_reg ( .CLK(n592), .EN(
        N1558), .ENCLK(net35137), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_12 clk_gate_reg_mstatus_mpp_reg ( .CLK(n592), 
        .EN(N335), .ENCLK(net35147), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_11 clk_gate_reg_mstatus_tsr_reg ( .CLK(n593), 
        .EN(N276), .ENCLK(net35152), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_10 clk_gate_reg_mstatus_mxr_reg ( .CLK(n593), 
        .EN(N290), .ENCLK(net35157), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_9 clk_gate_reg_dcsr_ebreakm_reg ( .CLK(n593), 
        .EN(N438), .ENCLK(net35162), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_8 clk_gate_reg_mideleg_reg ( .CLK(n593), .EN(
        N459), .ENCLK(net35167), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_7 clk_gate_reg_medeleg_reg ( .CLK(n593), .EN(
        N460), .ENCLK(net35172), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_6 clk_gate_reg_dcsr_cause_reg ( .CLK(n593), 
        .EN(N467), .ENCLK(net35177), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_5 clk_gate_reg_dpc_reg ( .CLK(n593), .EN(
        net35183), .ENCLK(net35304), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_4 clk_gate_reg_dscratch_reg ( .CLK(n593), .EN(
        N475), .ENCLK(net35309), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_3 clk_gate_reg_bp_0_control_dmode_reg ( .CLK(
        n593), .EN(N479), .ENCLK(net35314), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_2 clk_gate_reg_bp_0_control_tmatch_reg ( .CLK(
        n593), .EN(N487), .ENCLK(net35319), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_1 clk_gate__T_49_reg ( .CLK(n591), .EN(N1890), 
        .ENCLK(net35324), .TE(1'b0) );
  CSRFile_DW01_inc_J38_0 add_x_427 ( .A({io_pmp_7_addr[28:0], 
        io_pmp_7_cfg_a[0]}), .SUM({n_T_304, SYNOPSYS_UNCONNECTED_1}) );
  CSRFile_DW01_inc_J38_1 add_x_426 ( .A({io_pmp_6_addr[28:0], 
        io_pmp_6_cfg_a[0]}), .SUM({n_T_295, SYNOPSYS_UNCONNECTED_2}) );
  CSRFile_DW01_inc_J38_2 add_x_425 ( .A({io_pmp_5_addr[28:0], 
        io_pmp_5_cfg_a[0]}), .SUM({n_T_286, SYNOPSYS_UNCONNECTED_3}) );
  CSRFile_DW01_inc_J38_3 add_x_424 ( .A({io_pmp_4_addr[28:0], 
        io_pmp_4_cfg_a[0]}), .SUM({n_T_277, SYNOPSYS_UNCONNECTED_4}) );
  CSRFile_DW01_inc_J38_4 add_x_423 ( .A({io_pmp_3_addr[28:0], 
        io_pmp_3_cfg_a[0]}), .SUM({n_T_268, SYNOPSYS_UNCONNECTED_5}) );
  CSRFile_DW01_inc_J38_5 add_x_422 ( .A({io_pmp_2_addr[28:0], 
        io_pmp_2_cfg_a[0]}), .SUM({n_T_259, SYNOPSYS_UNCONNECTED_6}) );
  CSRFile_DW01_inc_J38_6 add_x_421 ( .A({io_pmp_1_addr[28:0], 
        io_pmp_1_cfg_a[0]}), .SUM({n_T_250, SYNOPSYS_UNCONNECTED_7}) );
  CSRFile_DW01_inc_J38_7 add_x_420 ( .A({io_pmp_0_addr[28:0], 
        io_pmp_0_cfg_a[0]}), .SUM({n_T_241, SYNOPSYS_UNCONNECTED_8}) );
  CSRFile_DW01_inc_J38_8 add_x_381 ( .A({n1936, n1937, n1938, n1939, n1940, 
        n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
        n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
        n1961, n1962, n1963, n1964, n1965, n1966, n1967, io_time[31:6]}), 
        .SUM({n_T_52, SYNOPSYS_UNCONNECTED_9}) );
  CSRFile_DW01_inc_J38_9 add_x_379 ( .A(n_T_45[63:6]), .SUM({n_T_44, 
        SYNOPSYS_UNCONNECTED_10}) );
  DFFX1_LVT reg_mip_seip_reg ( .D(n200), .CLK(n531), .Q(n_T_3694_9_) );
  DFFX1_LVT reg_mip_stip_reg ( .D(n199), .CLK(n531), .Q(n_T_61_5_) );
  DFFX1_LVT u_T_1579_reg ( .D(N1693), .CLK(net35147), .Q(n1918) );
  DFFX1_LVT u_T_47_reg_0_ ( .D(N1822), .CLK(n591), .Q(io_time[0]), .QN(n417)
         );
  DFFX1_LVT reg_stvec_reg_0_ ( .D(wdata[0]), .CLK(n568), .Q(n428), .QN(n658)
         );
  DFFX1_LVT reg_scounteren_reg_0_ ( .D(wdata[0]), .CLK(net34940), .Q(
        read_scounteren[0]) );
  DFFX1_LVT reg_mcounteren_reg_0_ ( .D(wdata[0]), .CLK(net34945), .Q(
        read_mcounteren[0]), .QN(n470) );
  DFFX1_LVT reg_medeleg_reg_0_ ( .D(wdata[0]), .CLK(net35172), .Q(
        read_medeleg_0) );
  DFFX1_LVT reg_dscratch_reg_0_ ( .D(wdata[0]), .CLK(n527), .Q(reg_dscratch[0]) );
  DFFX1_LVT reg_mscratch_reg_0_ ( .D(wdata[0]), .CLK(n553), .Q(reg_mscratch[0]) );
  DFFX1_LVT reg_sscratch_reg_0_ ( .D(wdata[0]), .CLK(n567), .Q(reg_sscratch[0]) );
  DFFX1_LVT u_T_39_reg_0_ ( .D(N1428), .CLK(n594), .Q(n_T_45[0]) );
  DFFX1_LVT reg_fflags_reg_0_ ( .D(n_GEN_345[0]), .CLK(n594), .Q(read_fcsr[0])
         );
  DFFX1_LVT reg_dcsr_prv_reg_0_ ( .D(n2156), .CLK(n594), .Q(n_T_389_0) );
  DFFX1_LVT reg_mstatus_mpp_reg_1_ ( .D(N334), .CLK(net35147), .Q(n[1929]) );
  DFFX1_LVT reg_stvec_reg_12_ ( .D(n367), .CLK(n568), .QN(reg_stvec[12]) );
  DFFSSRX1_LVT reg_mtvec_reg_12_ ( .D(n378), .SETB(wdata[12]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[12]) );
  DFFSSRX1_LVT reg_dcsr_ebreaku_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[12]), 
        .CLK(net35162), .Q(n_T_1155[0]) );
  DFFX1_LVT u_T_41_reg_6_ ( .D(N1503), .CLK(n579), .Q(n_T_45[12]) );
  DFFX1_LVT u_T_49_reg_6_ ( .D(N1897), .CLK(n521), .Q(io_time[12]) );
  DFFSSRX1_LVT reg_pmp_1_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[12]), .CLK(net35132), .Q(io_pmp_1_cfg_a[1]), .QN(n462) );
  DFFX1_LVT reg_pmp_0_addr_reg_0_ ( .D(n_GEN_258[0]), .CLK(n531), .Q(
        io_pmp_0_addr[0]) );
  DFFX1_LVT reg_pmp_0_addr_reg_9_ ( .D(n_GEN_258[9]), .CLK(n534), .Q(
        io_pmp_0_addr[9]), .QN(n419) );
  DFFX1_LVT reg_stvec_reg_9_ ( .D(wdata[9]), .CLK(n568), .Q(reg_stvec[9]) );
  DFFX1_LVT reg_mideleg_reg_9_ ( .D(wdata[9]), .CLK(net35167), .Q(
        read_mideleg_9_), .QN(n446) );
  DFFX1_LVT reg_mstatus_mpie_reg ( .D(N360), .CLK(net35147), .Q(n1932) );
  DFFX1_LVT reg_stvec_reg_7_ ( .D(wdata[7]), .CLK(n568), .Q(reg_stvec[7]) );
  DFFX1_LVT reg_dscratch_reg_7_ ( .D(wdata[7]), .CLK(n527), .Q(reg_dscratch[7]) );
  DFFX1_LVT reg_mscratch_reg_7_ ( .D(wdata[7]), .CLK(n553), .Q(reg_mscratch[7]) );
  DFFX1_LVT reg_sscratch_reg_7_ ( .D(wdata[7]), .CLK(n567), .Q(reg_sscratch[7]) );
  DFFSSRX1_LVT reg_mtvec_reg_7_ ( .D(n376), .SETB(wdata[7]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[7]) );
  DFFSSRX1_LVT reg_pmp_0_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[7]), 
        .CLK(net34905), .Q(io_pmp_0_cfg_l), .QN(n453) );
  DFFX1_LVT reg_pmp_0_cfg_r_reg ( .D(wdata[0]), .CLK(net34733), .Q(
        io_pmp_0_cfg_r) );
  DFFX1_LVT u_T_41_reg_1_ ( .D(N1498), .CLK(n579), .Q(n_T_45[7]) );
  DFFX1_LVT u_T_49_reg_1_ ( .D(N1892), .CLK(n521), .Q(io_time[7]) );
  DFFX1_LVT reg_mie_reg_7_ ( .D(N613), .CLK(net34728), .Q(reg_mie[7]) );
  DFFX1_LVT reg_frm_reg_2_ ( .D(n_GEN_155[2]), .CLK(net34900), .Q(
        io_fcsr_rm[2]) );
  DFFX1_LVT reg_stvec_reg_2_ ( .D(n1483), .CLK(n568), .QN(reg_stvec[2]) );
  DFFSSRX1_LVT reg_mtvec_reg_2_ ( .D(n376), .SETB(wdata[2]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[2]) );
  DFFSSRX1_LVT reg_dcsr_step_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[2]), 
        .CLK(net35162), .Q(n_T_389_2), .QN(n452) );
  DFFX1_LVT u_T_39_reg_2_ ( .D(N1430), .CLK(n594), .Q(n_T_45[2]) );
  DFFX1_LVT u_T_47_reg_2_ ( .D(N1824), .CLK(n591), .Q(io_time[2]) );
  DFFX1_LVT reg_pmp_0_addr_reg_2_ ( .D(n_GEN_258[2]), .CLK(n533), .Q(
        io_pmp_0_addr[2]) );
  DFFX1_LVT reg_fflags_reg_2_ ( .D(n_GEN_345[2]), .CLK(n594), .Q(read_fcsr[2]), 
        .QN(n477) );
  DFFX1_LVT reg_misa_reg_63_ ( .D(N1622), .CLK(net35137), .Q(n_T_3678_63_) );
  DFFX1_LVT reg_misa_reg_23_ ( .D(N1582), .CLK(net35137), .Q(n1919) );
  DFFX1_LVT reg_misa_reg_20_ ( .D(N1579), .CLK(net35137), .Q(n1920) );
  DFFX1_LVT reg_misa_reg_18_ ( .D(N1577), .CLK(net35137), .Q(n1921) );
  DFFX1_LVT reg_misa_reg_8_ ( .D(N1567), .CLK(net35137), .Q(n1922) );
  DFFX1_LVT reg_stvec_reg_8_ ( .D(wdata[8]), .CLK(n568), .Q(reg_stvec[8]) );
  DFFX1_LVT reg_medeleg_reg_8_ ( .D(wdata[8]), .CLK(net35172), .Q(
        read_medeleg_8) );
  DFFX1_LVT reg_dscratch_reg_8_ ( .D(wdata[8]), .CLK(n526), .Q(reg_dscratch[8]) );
  DFFX1_LVT reg_mscratch_reg_8_ ( .D(wdata[8]), .CLK(n552), .Q(reg_mscratch[8]) );
  DFFX1_LVT reg_sscratch_reg_8_ ( .D(wdata[8]), .CLK(n566), .Q(reg_sscratch[8]) );
  DFFSSRX1_LVT reg_mtvec_reg_8_ ( .D(n376), .SETB(wdata[8]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[8]) );
  DFFX1_LVT u_T_41_reg_2_ ( .D(N1499), .CLK(n579), .Q(n_T_45[8]) );
  DFFX1_LVT u_T_49_reg_2_ ( .D(N1893), .CLK(n521), .Q(io_time[8]) );
  DFFX1_LVT reg_mstatus_spp_reg ( .D(n1913), .CLK(n1915), .Q(n1931) );
  DFFX1_LVT reg_scause_reg_2_ ( .D(N1272), .CLK(n557), .Q(reg_scause[2]) );
  DFFX1_LVT reg_scause_reg_0_ ( .D(N1270), .CLK(n557), .Q(reg_scause[0]) );
  DFFX1_LVT reg_stval_reg_12_ ( .D(N1394), .CLK(n559), .Q(n_T_444[12]) );
  DFFX1_LVT reg_stval_reg_8_ ( .D(N1390), .CLK(n559), .Q(n_T_444[8]) );
  DFFX1_LVT reg_stval_reg_7_ ( .D(N1389), .CLK(n559), .Q(n_T_444[7]) );
  DFFX1_LVT reg_stval_reg_2_ ( .D(N1384), .CLK(n559), .Q(n_T_444[2]) );
  DFFX1_LVT reg_stval_reg_0_ ( .D(N1382), .CLK(n559), .Q(n_T_444[0]) );
  DFFX1_LVT reg_mtval_reg_12_ ( .D(N1005), .CLK(n572), .Q(n_T_383[12]) );
  DFFX1_LVT reg_mtval_reg_8_ ( .D(N1001), .CLK(n572), .Q(n_T_383[8]) );
  DFFX1_LVT reg_mtval_reg_7_ ( .D(N1000), .CLK(n572), .Q(n_T_383[7]) );
  DFFX1_LVT reg_mtval_reg_2_ ( .D(N995), .CLK(n572), .Q(n_T_383[2]) );
  DFFX1_LVT reg_mtval_reg_0_ ( .D(N993), .CLK(n572), .Q(n_T_383[0]) );
  DFFX1_LVT reg_mcause_reg_2_ ( .D(N883), .CLK(net34885), .Q(reg_mcause[2]) );
  DFFX1_LVT reg_mcause_reg_0_ ( .D(N881), .CLK(n580), .Q(reg_mcause[0]) );
  DFFX1_LVT reg_mepc_reg_2_ ( .D(net35076), .CLK(n545), .Q(reg_mepc[2]) );
  DFFX1_LVT reg_sepc_reg_2_ ( .D(net34874), .CLK(n581), .Q(reg_sepc[2]) );
  DFFX1_LVT reg_debug_reg ( .D(n2161), .CLK(n594), .Q(io_status_debug), .QN(
        io_status_debug_BAR) );
  DFFX1_LVT reg_singleStepped_reg ( .D(N435), .CLK(n594), .Q(n426), .QN(n860)
         );
  DFFX1_LVT reg_dpc_reg_2_ ( .D(net35298), .CLK(n528), .Q(reg_dpc[2]) );
  DFFX1_LVT reg_dcsr_cause_reg_1_ ( .D(N469), .CLK(net35177), .Q(n_T_389[7])
         );
  DFFX1_LVT reg_bp_0_control_tmatch_reg_1_ ( .D(wdata[8]), .CLK(net35319), .Q(
        io_bp_0_control_tmatch[1]) );
  DFFX1_LVT reg_bp_0_control_tmatch_reg_0_ ( .D(wdata[7]), .CLK(net35319), .Q(
        io_bp_0_control_tmatch[0]) );
  DFFX1_LVT reg_bp_0_control_dmode_reg ( .D(n1482), .CLK(net35314), .Q(
        n_T_366_59_), .QN(n457) );
  DFFX1_LVT reg_bp_0_control_action_reg ( .D(N485), .CLK(net35314), .Q(
        io_bp_0_control_action) );
  DFFSSRX1_LVT reg_bp_0_control_x_reg ( .D(n503), .SETB(1'b1), .RSTB(wdata[2]), 
        .CLK(net35314), .Q(io_bp_0_control_x) );
  DFFSSRX1_LVT reg_bp_0_control_r_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[0]), 
        .CLK(net35314), .Q(io_bp_0_control_r) );
  DFFX1_LVT reg_bp_0_address_reg_38_ ( .D(wdata[38]), .CLK(n584), .Q(
        io_bp_0_address[38]) );
  DFFX1_LVT reg_dscratch_reg_54_ ( .D(wdata[54]), .CLK(n526), .Q(
        reg_dscratch[54]) );
  DFFX1_LVT reg_mscratch_reg_54_ ( .D(wdata[54]), .CLK(n552), .Q(
        reg_mscratch[54]) );
  DFFX1_LVT reg_sscratch_reg_54_ ( .D(wdata[54]), .CLK(n566), .Q(
        reg_sscratch[54]) );
  DFFX1_LVT u_T_49_reg_48_ ( .D(N1939), .CLK(n521), .Q(n1945) );
  DFFX1_LVT reg_dscratch_reg_53_ ( .D(wdata[53]), .CLK(n526), .Q(
        reg_dscratch[53]) );
  DFFX1_LVT reg_mscratch_reg_53_ ( .D(wdata[53]), .CLK(n552), .Q(
        reg_mscratch[53]) );
  DFFX1_LVT reg_sscratch_reg_53_ ( .D(wdata[53]), .CLK(n566), .Q(
        reg_sscratch[53]) );
  DFFX1_LVT u_T_41_reg_47_ ( .D(N1544), .CLK(n579), .Q(n_T_45[53]) );
  DFFX1_LVT u_T_49_reg_47_ ( .D(N1938), .CLK(n521), .Q(n1946) );
  DFFX1_LVT reg_dscratch_reg_47_ ( .D(wdata[47]), .CLK(n526), .Q(
        reg_dscratch[47]) );
  DFFX1_LVT reg_mscratch_reg_47_ ( .D(wdata[47]), .CLK(n552), .Q(
        reg_mscratch[47]) );
  DFFX1_LVT reg_sscratch_reg_47_ ( .D(wdata[47]), .CLK(n566), .Q(
        reg_sscratch[47]) );
  DFFSSRX1_LVT reg_pmp_5_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[47]), 
        .CLK(net35112), .Q(io_pmp_5_cfg_l), .QN(n437) );
  DFFX1_LVT u_T_41_reg_41_ ( .D(N1538), .CLK(n579), .Q(n_T_45[47]) );
  DFFX1_LVT u_T_49_reg_41_ ( .D(N1932), .CLK(n521), .Q(n1952) );
  DFFX1_LVT reg_dscratch_reg_46_ ( .D(wdata[46]), .CLK(n526), .Q(
        reg_dscratch[46]) );
  DFFX1_LVT reg_mscratch_reg_46_ ( .D(wdata[46]), .CLK(n552), .Q(
        reg_mscratch[46]) );
  DFFX1_LVT reg_sscratch_reg_46_ ( .D(wdata[46]), .CLK(n566), .Q(
        reg_sscratch[46]) );
  DFFX1_LVT u_T_41_reg_40_ ( .D(N1537), .CLK(n579), .Q(n_T_45[46]) );
  DFFX1_LVT u_T_49_reg_40_ ( .D(N1931), .CLK(n521), .Q(n1953) );
  DFFX1_LVT reg_dscratch_reg_45_ ( .D(wdata[45]), .CLK(n526), .Q(
        reg_dscratch[45]) );
  DFFX1_LVT reg_mscratch_reg_45_ ( .D(wdata[45]), .CLK(n552), .Q(
        reg_mscratch[45]) );
  DFFX1_LVT reg_sscratch_reg_45_ ( .D(wdata[45]), .CLK(n566), .Q(
        reg_sscratch[45]) );
  DFFX1_LVT u_T_41_reg_39_ ( .D(N1536), .CLK(n579), .Q(n_T_45[45]) );
  DFFX1_LVT u_T_49_reg_39_ ( .D(N1930), .CLK(n521), .Q(n1954) );
  DFFX1_LVT reg_dscratch_reg_44_ ( .D(wdata[44]), .CLK(n526), .Q(
        reg_dscratch[44]) );
  DFFX1_LVT reg_mscratch_reg_44_ ( .D(wdata[44]), .CLK(n552), .Q(
        reg_mscratch[44]) );
  DFFX1_LVT reg_sscratch_reg_44_ ( .D(wdata[44]), .CLK(n566), .Q(
        reg_sscratch[44]) );
  DFFSSRX1_LVT reg_pmp_5_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[44]), .CLK(net35112), .Q(io_pmp_5_cfg_a[1]), .QN(n461) );
  DFFX1_LVT u_T_41_reg_38_ ( .D(N1535), .CLK(n579), .Q(n_T_45[44]) );
  DFFX1_LVT u_T_49_reg_38_ ( .D(N1929), .CLK(n521), .Q(n1955) );
  DFFX1_LVT reg_dscratch_reg_43_ ( .D(wdata[43]), .CLK(n526), .Q(
        reg_dscratch[43]) );
  DFFX1_LVT reg_mscratch_reg_43_ ( .D(wdata[43]), .CLK(n552), .Q(
        reg_mscratch[43]) );
  DFFX1_LVT reg_sscratch_reg_43_ ( .D(wdata[43]), .CLK(n566), .Q(
        reg_sscratch[43]) );
  DFFSSRX1_LVT reg_pmp_5_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[43]), .CLK(net35112), .Q(io_pmp_5_cfg_a[0]) );
  DFFX1_LVT u_T_41_reg_37_ ( .D(N1534), .CLK(n579), .Q(n_T_45[43]) );
  DFFX1_LVT u_T_49_reg_37_ ( .D(N1928), .CLK(n521), .Q(n1956) );
  DFFX1_LVT reg_dscratch_reg_42_ ( .D(wdata[42]), .CLK(n526), .Q(
        reg_dscratch[42]) );
  DFFX1_LVT reg_pmp_5_cfg_x_reg ( .D(wdata[42]), .CLK(net35097), .Q(
        io_pmp_5_cfg_x) );
  DFFX1_LVT reg_mscratch_reg_42_ ( .D(wdata[42]), .CLK(n552), .Q(
        reg_mscratch[42]) );
  DFFX1_LVT reg_sscratch_reg_42_ ( .D(wdata[42]), .CLK(n566), .Q(
        reg_sscratch[42]) );
  DFFX1_LVT u_T_41_reg_36_ ( .D(N1533), .CLK(n578), .Q(n_T_45[42]) );
  DFFX1_LVT u_T_49_reg_36_ ( .D(N1927), .CLK(n520), .Q(n1957) );
  DFFX1_LVT reg_dscratch_reg_40_ ( .D(wdata[40]), .CLK(n526), .Q(
        reg_dscratch[40]) );
  DFFX1_LVT reg_pmp_5_cfg_r_reg ( .D(wdata[40]), .CLK(net35097), .Q(
        io_pmp_5_cfg_r) );
  DFFX1_LVT reg_mscratch_reg_40_ ( .D(wdata[40]), .CLK(n552), .Q(
        reg_mscratch[40]) );
  DFFX1_LVT reg_sscratch_reg_40_ ( .D(wdata[40]), .CLK(n566), .Q(
        reg_sscratch[40]) );
  DFFX1_LVT u_T_41_reg_34_ ( .D(N1531), .CLK(n578), .Q(n_T_45[40]) );
  DFFX1_LVT u_T_49_reg_34_ ( .D(N1925), .CLK(n520), .Q(n1959) );
  DFFSSRX1_LVT reg_pmp_5_cfg_w_reg ( .D(wdata[40]), .SETB(1'b1), .RSTB(
        wdata[41]), .CLK(net35097), .Q(io_pmp_5_cfg_w) );
  DFFX1_LVT reg_dscratch_reg_41_ ( .D(wdata[41]), .CLK(n526), .Q(
        reg_dscratch[41]) );
  DFFX1_LVT reg_mscratch_reg_41_ ( .D(wdata[41]), .CLK(n552), .Q(
        reg_mscratch[41]) );
  DFFX1_LVT reg_sscratch_reg_41_ ( .D(wdata[41]), .CLK(n566), .Q(
        reg_sscratch[41]) );
  DFFX1_LVT u_T_41_reg_35_ ( .D(N1532), .CLK(n578), .Q(n_T_45[41]) );
  DFFX1_LVT u_T_49_reg_35_ ( .D(N1926), .CLK(n520), .Q(n1958) );
  DFFX1_LVT reg_dscratch_reg_62_ ( .D(wdata[62]), .CLK(n526), .Q(
        reg_dscratch[62]) );
  DFFX1_LVT reg_mscratch_reg_62_ ( .D(wdata[62]), .CLK(n552), .Q(
        reg_mscratch[62]) );
  DFFX1_LVT reg_sscratch_reg_62_ ( .D(wdata[62]), .CLK(n566), .Q(
        reg_sscratch[62]) );
  DFFX1_LVT u_T_41_reg_56_ ( .D(N1553), .CLK(n578), .Q(n_T_45[62]) );
  DFFX1_LVT u_T_49_reg_56_ ( .D(N1947), .CLK(n520), .Q(n1937) );
  DFFX1_LVT reg_dscratch_reg_39_ ( .D(wdata[39]), .CLK(n525), .Q(
        reg_dscratch[39]) );
  DFFX1_LVT reg_mscratch_reg_39_ ( .D(wdata[39]), .CLK(n551), .Q(
        reg_mscratch[39]) );
  DFFX1_LVT reg_sscratch_reg_39_ ( .D(wdata[39]), .CLK(n565), .Q(
        reg_sscratch[39]) );
  DFFX1_LVT reg_mtval_reg_39_ ( .D(N1032), .CLK(n572), .Q(n_T_383[39]) );
  DFFX1_LVT reg_stval_reg_39_ ( .D(N1421), .CLK(n559), .Q(n_T_444[39]) );
  DFFSSRX1_LVT reg_pmp_4_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[39]), 
        .CLK(net34910), .Q(io_pmp_4_cfg_l), .QN(n438) );
  DFFX1_LVT reg_pmp_4_addr_reg_0_ ( .D(n_GEN_286[0]), .CLK(n532), .Q(
        io_pmp_4_addr[0]) );
  DFFX1_LVT reg_pmp_4_addr_reg_2_ ( .D(n_GEN_286[2]), .CLK(n538), .Q(
        io_pmp_4_addr[2]) );
  DFFX1_LVT u_T_41_reg_33_ ( .D(N1530), .CLK(n578), .Q(n_T_45[39]) );
  DFFX1_LVT u_T_49_reg_33_ ( .D(N1924), .CLK(n520), .Q(n1960) );
  DFFX1_LVT reg_sepc_reg_39_ ( .D(net34763), .CLK(n581), .Q(reg_sepc[39]) );
  DFFX1_LVT reg_mepc_reg_39_ ( .D(net34965), .CLK(n545), .Q(reg_mepc[39]) );
  DFFX1_LVT reg_dpc_reg_39_ ( .D(net35187), .CLK(n528), .Q(reg_dpc[39]) );
  DFFX1_LVT reg_dscratch_reg_61_ ( .D(wdata[61]), .CLK(n525), .Q(
        reg_dscratch[61]) );
  DFFX1_LVT reg_mscratch_reg_61_ ( .D(wdata[61]), .CLK(n551), .Q(
        reg_mscratch[61]) );
  DFFX1_LVT reg_sscratch_reg_61_ ( .D(wdata[61]), .CLK(n565), .Q(
        reg_sscratch[61]) );
  DFFX1_LVT u_T_41_reg_55_ ( .D(N1552), .CLK(n578), .Q(n_T_45[61]) );
  DFFX1_LVT u_T_49_reg_55_ ( .D(N1946), .CLK(n520), .Q(n1938) );
  DFFX1_LVT reg_dscratch_reg_55_ ( .D(wdata[55]), .CLK(n525), .Q(
        reg_dscratch[55]) );
  DFFX1_LVT reg_mscratch_reg_55_ ( .D(wdata[55]), .CLK(n551), .Q(
        reg_mscratch[55]) );
  DFFX1_LVT reg_sscratch_reg_55_ ( .D(wdata[55]), .CLK(n565), .Q(
        reg_sscratch[55]) );
  DFFX1_LVT reg_pmp_6_cfg_r_reg ( .D(wdata[48]), .CLK(net35107), .Q(
        io_pmp_6_cfg_r) );
  DFFX1_LVT reg_dscratch_reg_48_ ( .D(wdata[48]), .CLK(n525), .Q(
        reg_dscratch[48]) );
  DFFX1_LVT reg_mscratch_reg_48_ ( .D(wdata[48]), .CLK(n551), .Q(
        reg_mscratch[48]) );
  DFFX1_LVT reg_sscratch_reg_48_ ( .D(wdata[48]), .CLK(n565), .Q(
        reg_sscratch[48]) );
  DFFX1_LVT u_T_41_reg_42_ ( .D(N1539), .CLK(n578), .Q(n_T_45[48]) );
  DFFX1_LVT u_T_49_reg_42_ ( .D(N1933), .CLK(n520), .Q(n1951) );
  DFFX1_LVT reg_dscratch_reg_49_ ( .D(wdata[49]), .CLK(n525), .Q(
        reg_dscratch[49]) );
  DFFX1_LVT reg_mscratch_reg_49_ ( .D(wdata[49]), .CLK(n551), .Q(
        reg_mscratch[49]) );
  DFFX1_LVT reg_sscratch_reg_49_ ( .D(wdata[49]), .CLK(n565), .Q(
        reg_sscratch[49]) );
  DFFX1_LVT u_T_41_reg_43_ ( .D(N1540), .CLK(n578), .Q(n_T_45[49]) );
  DFFX1_LVT u_T_49_reg_43_ ( .D(N1934), .CLK(n520), .Q(n1950) );
  DFFX1_LVT reg_pmp_6_cfg_x_reg ( .D(wdata[50]), .CLK(net35107), .Q(
        io_pmp_6_cfg_x) );
  DFFX1_LVT reg_dscratch_reg_50_ ( .D(wdata[50]), .CLK(n525), .Q(
        reg_dscratch[50]) );
  DFFX1_LVT reg_mscratch_reg_50_ ( .D(wdata[50]), .CLK(n551), .Q(
        reg_mscratch[50]) );
  DFFX1_LVT reg_sscratch_reg_50_ ( .D(wdata[50]), .CLK(n565), .Q(
        reg_sscratch[50]) );
  DFFX1_LVT u_T_41_reg_44_ ( .D(N1541), .CLK(n578), .Q(n_T_45[50]) );
  DFFX1_LVT u_T_49_reg_44_ ( .D(N1935), .CLK(n520), .Q(n1949) );
  DFFSSRX1_LVT reg_pmp_6_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[52]), .CLK(net35102), .Q(io_pmp_6_cfg_a[1]), .QN(n458) );
  DFFX1_LVT reg_dscratch_reg_52_ ( .D(wdata[52]), .CLK(n525), .Q(
        reg_dscratch[52]) );
  DFFX1_LVT reg_mscratch_reg_52_ ( .D(wdata[52]), .CLK(n551), .Q(
        reg_mscratch[52]) );
  DFFX1_LVT reg_sscratch_reg_52_ ( .D(wdata[52]), .CLK(n565), .Q(
        reg_sscratch[52]) );
  DFFX1_LVT u_T_41_reg_46_ ( .D(N1543), .CLK(n578), .Q(n_T_45[52]) );
  DFFX1_LVT u_T_49_reg_46_ ( .D(N1937), .CLK(n520), .Q(n1947) );
  DFFSSRX1_LVT reg_pmp_6_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[51]), .CLK(net35102), .Q(io_pmp_6_cfg_a[0]) );
  DFFX1_LVT reg_dscratch_reg_51_ ( .D(wdata[51]), .CLK(n525), .Q(
        reg_dscratch[51]) );
  DFFX1_LVT reg_mscratch_reg_51_ ( .D(wdata[51]), .CLK(n551), .Q(
        reg_mscratch[51]) );
  DFFX1_LVT reg_sscratch_reg_51_ ( .D(wdata[51]), .CLK(n565), .Q(
        reg_sscratch[51]) );
  DFFX1_LVT u_T_41_reg_45_ ( .D(N1542), .CLK(n578), .Q(n_T_45[51]) );
  DFFX1_LVT u_T_49_reg_45_ ( .D(N1936), .CLK(n520), .Q(n1948) );
  DFFX1_LVT reg_pmp_5_addr_reg_0_ ( .D(n_GEN_293[0]), .CLK(n540), .Q(
        io_pmp_5_addr[0]) );
  DFFX1_LVT reg_pmp_5_addr_reg_2_ ( .D(n_GEN_293[2]), .CLK(n539), .Q(
        io_pmp_5_addr[2]) );
  DFFX1_LVT u_T_41_reg_49_ ( .D(N1546), .CLK(n578), .Q(n_T_45[55]) );
  DFFX1_LVT u_T_49_reg_49_ ( .D(N1940), .CLK(n520), .Q(n1944) );
  DFFX1_LVT reg_stvec_reg_38_ ( .D(wdata[38]), .CLK(n568), .Q(reg_stvec[38]), 
        .QN(n465) );
  DFFX1_LVT reg_dscratch_reg_38_ ( .D(wdata[38]), .CLK(n525), .Q(
        reg_dscratch[38]) );
  DFFX1_LVT reg_mscratch_reg_38_ ( .D(wdata[38]), .CLK(n551), .Q(
        reg_mscratch[38]) );
  DFFX1_LVT reg_sscratch_reg_38_ ( .D(wdata[38]), .CLK(n565), .Q(
        reg_sscratch[38]) );
  DFFX1_LVT reg_mtval_reg_38_ ( .D(N1031), .CLK(n572), .Q(n_T_383[38]) );
  DFFX1_LVT reg_stval_reg_38_ ( .D(N1420), .CLK(n559), .Q(n_T_444[38]) );
  DFFX1_LVT u_T_41_reg_32_ ( .D(N1529), .CLK(n577), .Q(n_T_45[38]) );
  DFFX1_LVT u_T_49_reg_32_ ( .D(N1923), .CLK(n519), .Q(n1961) );
  DFFX1_LVT reg_sepc_reg_38_ ( .D(net34766), .CLK(n581), .Q(reg_sepc[38]) );
  DFFX1_LVT reg_mepc_reg_38_ ( .D(net34968), .CLK(n545), .Q(reg_mepc[38]) );
  DFFX1_LVT reg_dpc_reg_38_ ( .D(net35190), .CLK(n528), .Q(reg_dpc[38]) );
  DFFX1_LVT reg_bp_0_address_reg_37_ ( .D(wdata[37]), .CLK(n584), .Q(
        io_bp_0_address[37]) );
  DFFX1_LVT reg_stvec_reg_37_ ( .D(wdata[37]), .CLK(n568), .Q(reg_stvec[37])
         );
  DFFX1_LVT reg_dscratch_reg_37_ ( .D(wdata[37]), .CLK(n525), .Q(
        reg_dscratch[37]) );
  DFFX1_LVT reg_mscratch_reg_37_ ( .D(wdata[37]), .CLK(n551), .Q(
        reg_mscratch[37]) );
  DFFX1_LVT reg_sscratch_reg_37_ ( .D(wdata[37]), .CLK(n565), .Q(
        reg_sscratch[37]) );
  DFFX1_LVT reg_mtval_reg_37_ ( .D(N1030), .CLK(n572), .Q(n_T_383[37]) );
  DFFX1_LVT reg_stval_reg_37_ ( .D(N1419), .CLK(n559), .Q(n_T_444[37]) );
  DFFX1_LVT u_T_41_reg_31_ ( .D(N1528), .CLK(n577), .Q(n_T_45[37]) );
  DFFX1_LVT u_T_49_reg_31_ ( .D(N1922), .CLK(n519), .Q(n1962) );
  DFFX1_LVT reg_sepc_reg_37_ ( .D(net34769), .CLK(n581), .Q(reg_sepc[37]) );
  DFFX1_LVT reg_mepc_reg_37_ ( .D(net34971), .CLK(n545), .Q(reg_mepc[37]) );
  DFFX1_LVT reg_dpc_reg_37_ ( .D(net35193), .CLK(n528), .Q(reg_dpc[37]) );
  DFFX1_LVT reg_bp_0_address_reg_36_ ( .D(wdata[36]), .CLK(n584), .Q(
        io_bp_0_address[36]) );
  DFFX1_LVT reg_stvec_reg_36_ ( .D(wdata[36]), .CLK(n568), .Q(reg_stvec[36])
         );
  DFFX1_LVT reg_dscratch_reg_36_ ( .D(wdata[36]), .CLK(n525), .Q(
        reg_dscratch[36]) );
  DFFX1_LVT reg_mscratch_reg_36_ ( .D(wdata[36]), .CLK(n551), .Q(
        reg_mscratch[36]) );
  DFFX1_LVT reg_sscratch_reg_36_ ( .D(wdata[36]), .CLK(n565), .Q(
        reg_sscratch[36]) );
  DFFX1_LVT reg_mtval_reg_36_ ( .D(N1029), .CLK(n572), .Q(n_T_383[36]) );
  DFFX1_LVT reg_stval_reg_36_ ( .D(N1418), .CLK(n559), .Q(n_T_444[36]) );
  DFFSSRX1_LVT reg_pmp_4_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[36]), .CLK(net34910), .Q(io_pmp_4_cfg_a[1]), .QN(n464) );
  DFFX1_LVT u_T_41_reg_30_ ( .D(N1527), .CLK(n577), .Q(n_T_45[36]) );
  DFFX1_LVT u_T_49_reg_30_ ( .D(N1921), .CLK(n519), .Q(n1963) );
  DFFX1_LVT reg_sepc_reg_36_ ( .D(net34772), .CLK(n581), .Q(reg_sepc[36]) );
  DFFX1_LVT reg_mepc_reg_36_ ( .D(net34974), .CLK(n545), .Q(reg_mepc[36]) );
  DFFX1_LVT reg_dpc_reg_36_ ( .D(net35196), .CLK(n528), .Q(reg_dpc[36]) );
  DFFX1_LVT reg_bp_0_address_reg_35_ ( .D(wdata[35]), .CLK(n584), .Q(
        io_bp_0_address[35]) );
  DFFX1_LVT reg_stvec_reg_35_ ( .D(wdata[35]), .CLK(n568), .Q(reg_stvec[35])
         );
  DFFX1_LVT reg_dscratch_reg_35_ ( .D(wdata[35]), .CLK(n525), .Q(
        reg_dscratch[35]) );
  DFFX1_LVT reg_mscratch_reg_35_ ( .D(wdata[35]), .CLK(n551), .Q(
        reg_mscratch[35]) );
  DFFX1_LVT reg_sscratch_reg_35_ ( .D(wdata[35]), .CLK(n565), .Q(
        reg_sscratch[35]) );
  DFFX1_LVT reg_mtval_reg_35_ ( .D(N1028), .CLK(n572), .Q(n_T_383[35]) );
  DFFX1_LVT reg_stval_reg_35_ ( .D(N1417), .CLK(n559), .Q(n_T_444[35]) );
  DFFSSRX1_LVT reg_pmp_4_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[35]), .CLK(net34910), .Q(io_pmp_4_cfg_a[0]) );
  DFFX1_LVT u_T_41_reg_29_ ( .D(N1526), .CLK(n577), .Q(n_T_45[35]) );
  DFFX1_LVT u_T_49_reg_29_ ( .D(N1920), .CLK(n519), .Q(n1964) );
  DFFX1_LVT reg_sepc_reg_35_ ( .D(net34775), .CLK(n581), .Q(reg_sepc[35]) );
  DFFX1_LVT reg_mepc_reg_35_ ( .D(net34977), .CLK(n545), .Q(reg_mepc[35]) );
  DFFX1_LVT reg_dpc_reg_35_ ( .D(net35199), .CLK(n528), .Q(reg_dpc[35]) );
  DFFX1_LVT reg_bp_0_address_reg_34_ ( .D(wdata[34]), .CLK(n584), .Q(
        io_bp_0_address[34]) );
  DFFX1_LVT reg_stvec_reg_34_ ( .D(wdata[34]), .CLK(n568), .Q(reg_stvec[34])
         );
  DFFX1_LVT reg_dscratch_reg_34_ ( .D(wdata[34]), .CLK(n524), .Q(
        reg_dscratch[34]) );
  DFFX1_LVT reg_pmp_4_cfg_x_reg ( .D(wdata[34]), .CLK(net35117), .Q(
        io_pmp_4_cfg_x) );
  DFFX1_LVT reg_mscratch_reg_34_ ( .D(wdata[34]), .CLK(n550), .Q(
        reg_mscratch[34]) );
  DFFX1_LVT reg_sscratch_reg_34_ ( .D(wdata[34]), .CLK(n564), .Q(
        reg_sscratch[34]) );
  DFFX1_LVT reg_mtval_reg_34_ ( .D(N1027), .CLK(n572), .Q(n_T_383[34]) );
  DFFX1_LVT reg_stval_reg_34_ ( .D(N1416), .CLK(n559), .Q(n_T_444[34]) );
  DFFX1_LVT u_T_41_reg_28_ ( .D(N1525), .CLK(n577), .Q(n_T_45[34]) );
  DFFX1_LVT u_T_49_reg_28_ ( .D(N1919), .CLK(n519), .Q(n1965) );
  DFFX1_LVT reg_sepc_reg_34_ ( .D(net34778), .CLK(n581), .Q(reg_sepc[34]) );
  DFFX1_LVT reg_mepc_reg_34_ ( .D(net34980), .CLK(n545), .Q(reg_mepc[34]) );
  DFFX1_LVT reg_dpc_reg_34_ ( .D(net35202), .CLK(n528), .Q(reg_dpc[34]) );
  DFFX1_LVT reg_bp_0_address_reg_32_ ( .D(wdata[32]), .CLK(n584), .Q(
        io_bp_0_address[32]) );
  DFFX1_LVT reg_stvec_reg_32_ ( .D(wdata[32]), .CLK(n568), .Q(reg_stvec[32])
         );
  DFFX1_LVT reg_dscratch_reg_32_ ( .D(wdata[32]), .CLK(n524), .Q(
        reg_dscratch[32]) );
  DFFX1_LVT reg_pmp_4_cfg_r_reg ( .D(wdata[32]), .CLK(net35117), .Q(
        io_pmp_4_cfg_r) );
  DFFX1_LVT reg_mscratch_reg_32_ ( .D(wdata[32]), .CLK(n550), .Q(
        reg_mscratch[32]) );
  DFFX1_LVT reg_sscratch_reg_32_ ( .D(wdata[32]), .CLK(n564), .Q(
        reg_sscratch[32]) );
  DFFX1_LVT reg_mtval_reg_32_ ( .D(N1025), .CLK(n572), .Q(n_T_383[32]) );
  DFFX1_LVT reg_stval_reg_32_ ( .D(N1414), .CLK(n559), .Q(n_T_444[32]) );
  DFFX1_LVT u_T_41_reg_26_ ( .D(N1523), .CLK(n577), .Q(n_T_45[32]) );
  DFFX1_LVT u_T_49_reg_26_ ( .D(N1917), .CLK(n519), .Q(n1967) );
  DFFSSRX1_LVT reg_pmp_4_cfg_w_reg ( .D(wdata[32]), .SETB(1'b1), .RSTB(
        wdata[33]), .CLK(net35117), .Q(io_pmp_4_cfg_w) );
  DFFX1_LVT reg_stvec_reg_33_ ( .D(wdata[33]), .CLK(n569), .Q(reg_stvec[33])
         );
  DFFX1_LVT reg_dscratch_reg_33_ ( .D(wdata[33]), .CLK(n524), .Q(
        reg_dscratch[33]) );
  DFFX1_LVT reg_mscratch_reg_33_ ( .D(wdata[33]), .CLK(n550), .Q(
        reg_mscratch[33]) );
  DFFX1_LVT reg_sscratch_reg_33_ ( .D(wdata[33]), .CLK(n564), .Q(
        reg_sscratch[33]) );
  DFFX1_LVT reg_bp_0_address_reg_33_ ( .D(wdata[33]), .CLK(n584), .Q(
        io_bp_0_address[33]) );
  DFFX1_LVT reg_mtval_reg_33_ ( .D(N1026), .CLK(n573), .Q(n_T_383[33]) );
  DFFX1_LVT reg_stval_reg_33_ ( .D(N1415), .CLK(n560), .Q(n_T_444[33]) );
  DFFX1_LVT u_T_41_reg_27_ ( .D(N1524), .CLK(n577), .Q(n_T_45[33]) );
  DFFX1_LVT u_T_49_reg_27_ ( .D(N1918), .CLK(n519), .Q(n1966) );
  DFFX1_LVT reg_sepc_reg_33_ ( .D(net34781), .CLK(n581), .Q(reg_sepc[33]) );
  DFFX1_LVT reg_mepc_reg_33_ ( .D(net34983), .CLK(n545), .Q(reg_mepc[33]) );
  DFFX1_LVT reg_dpc_reg_33_ ( .D(net35205), .CLK(n528), .Q(reg_dpc[33]) );
  DFFX1_LVT reg_sepc_reg_32_ ( .D(net34784), .CLK(n581), .Q(reg_sepc[32]) );
  DFFX1_LVT reg_mepc_reg_32_ ( .D(net34986), .CLK(n545), .Q(reg_mepc[32]) );
  DFFX1_LVT reg_dpc_reg_32_ ( .D(net35208), .CLK(n528), .Q(reg_dpc[32]) );
  DFFX1_LVT reg_bp_0_address_reg_31_ ( .D(wdata[31]), .CLK(n584), .Q(
        io_bp_0_address[31]) );
  DFFX1_LVT reg_stvec_reg_31_ ( .D(wdata[31]), .CLK(n569), .Q(reg_stvec[31])
         );
  DFFX1_LVT reg_dscratch_reg_31_ ( .D(wdata[31]), .CLK(n524), .Q(
        reg_dscratch[31]) );
  DFFX1_LVT reg_mscratch_reg_31_ ( .D(wdata[31]), .CLK(n550), .Q(
        reg_mscratch[31]) );
  DFFX1_LVT reg_sscratch_reg_31_ ( .D(wdata[31]), .CLK(n564), .Q(
        reg_sscratch[31]) );
  DFFX1_LVT reg_mtval_reg_31_ ( .D(N1024), .CLK(n573), .Q(n_T_383[31]) );
  DFFX1_LVT reg_stval_reg_31_ ( .D(N1413), .CLK(n560), .Q(n_T_444[31]) );
  DFFSSRX1_LVT reg_pmp_3_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[31]), 
        .CLK(net35127), .Q(io_pmp_3_cfg_l), .QN(n443) );
  DFFX1_LVT reg_pmp_3_addr_reg_0_ ( .D(n_GEN_279[0]), .CLK(n537), .Q(
        io_pmp_3_addr[0]) );
  DFFX1_LVT reg_pmp_3_addr_reg_2_ ( .D(n_GEN_279[2]), .CLK(n536), .Q(
        io_pmp_3_addr[2]) );
  DFFX1_LVT u_T_41_reg_25_ ( .D(N1522), .CLK(n577), .Q(n_T_45[31]) );
  DFFX1_LVT u_T_49_reg_25_ ( .D(N1916), .CLK(n519), .Q(io_time[31]) );
  DFFX1_LVT reg_sepc_reg_31_ ( .D(net34787), .CLK(n581), .Q(reg_sepc[31]) );
  DFFX1_LVT reg_mepc_reg_31_ ( .D(net34989), .CLK(n545), .Q(reg_mepc[31]) );
  DFFX1_LVT reg_dpc_reg_31_ ( .D(net35211), .CLK(n528), .Q(reg_dpc[31]) );
  DFFX1_LVT reg_bp_0_address_reg_30_ ( .D(wdata[30]), .CLK(n584), .Q(
        io_bp_0_address[30]) );
  DFFX1_LVT reg_stvec_reg_30_ ( .D(wdata[30]), .CLK(n569), .Q(reg_stvec[30])
         );
  DFFX1_LVT reg_dscratch_reg_30_ ( .D(wdata[30]), .CLK(n524), .Q(
        reg_dscratch[30]) );
  DFFX1_LVT reg_mscratch_reg_30_ ( .D(wdata[30]), .CLK(n550), .Q(
        reg_mscratch[30]) );
  DFFX1_LVT reg_sscratch_reg_30_ ( .D(wdata[30]), .CLK(n564), .Q(
        reg_sscratch[30]) );
  DFFX1_LVT reg_mtval_reg_30_ ( .D(N1023), .CLK(n573), .Q(n_T_383[30]) );
  DFFSSRX1_LVT reg_mtvec_reg_30_ ( .D(n376), .SETB(wdata[30]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[30]) );
  DFFX1_LVT reg_stval_reg_30_ ( .D(N1412), .CLK(n560), .Q(n_T_444[30]) );
  DFFX1_LVT u_T_41_reg_24_ ( .D(N1521), .CLK(n577), .Q(n_T_45[30]) );
  DFFX1_LVT u_T_49_reg_24_ ( .D(N1915), .CLK(n519), .Q(io_time[30]) );
  DFFX1_LVT reg_sepc_reg_30_ ( .D(net34790), .CLK(n581), .Q(reg_sepc[30]) );
  DFFX1_LVT reg_mepc_reg_30_ ( .D(net34992), .CLK(n545), .Q(reg_mepc[30]) );
  DFFX1_LVT reg_dpc_reg_30_ ( .D(net35214), .CLK(n528), .Q(reg_dpc[30]) );
  DFFX1_LVT reg_bp_0_address_reg_13_ ( .D(wdata[13]), .CLK(n584), .Q(
        io_bp_0_address[13]) );
  DFFX1_LVT reg_stvec_reg_13_ ( .D(wdata[13]), .CLK(n569), .Q(reg_stvec[13])
         );
  DFFX1_LVT reg_medeleg_reg_13_ ( .D(wdata[13]), .CLK(net35172), .Q(
        read_medeleg_13) );
  DFFX1_LVT reg_dscratch_reg_13_ ( .D(wdata[13]), .CLK(n524), .Q(
        reg_dscratch[13]) );
  DFFX1_LVT reg_mscratch_reg_13_ ( .D(wdata[13]), .CLK(n550), .Q(
        reg_mscratch[13]) );
  DFFX1_LVT reg_sscratch_reg_13_ ( .D(wdata[13]), .CLK(n564), .Q(
        reg_sscratch[13]) );
  DFFX1_LVT reg_mtval_reg_13_ ( .D(N1006), .CLK(n573), .Q(n_T_383[13]) );
  DFFSSRX1_LVT reg_mtvec_reg_13_ ( .D(n376), .SETB(wdata[13]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[13]) );
  DFFX1_LVT reg_stval_reg_13_ ( .D(N1395), .CLK(n560), .Q(n_T_444[13]) );
  DFFSSRX1_LVT reg_dcsr_ebreaks_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[13]), 
        .CLK(net35162), .Q(n_T_1155[1]) );
  DFFX1_LVT u_T_41_reg_7_ ( .D(N1504), .CLK(n577), .Q(n_T_45[13]) );
  DFFX1_LVT u_T_49_reg_7_ ( .D(N1898), .CLK(n519), .Q(io_time[13]) );
  DFFSSRX1_LVT reg_mstatus_fs_reg_1_ ( .D(wdata[13]), .SETB(n51), .RSTB(n375), 
        .CLK(net35157), .Q(n1928) );
  DFFX1_LVT reg_dscratch_reg_63_ ( .D(wdata[63]), .CLK(n524), .Q(
        reg_dscratch[63]) );
  DFFX1_LVT reg_mscratch_reg_63_ ( .D(wdata[63]), .CLK(n550), .Q(
        reg_mscratch[63]) );
  DFFX1_LVT reg_sscratch_reg_63_ ( .D(wdata[63]), .CLK(n564), .Q(
        reg_sscratch[63]) );
  DFFX1_LVT reg_scause_reg_63_ ( .D(N1333), .CLK(n558), .Q(reg_scause[63]) );
  DFFSSRX1_LVT reg_pmp_7_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[63]), 
        .CLK(net34743), .Q(io_pmp_7_cfg_l), .QN(n442) );
  DFFX1_LVT reg_pmp_7_cfg_r_reg ( .D(wdata[56]), .CLK(net34738), .Q(
        io_pmp_7_cfg_r) );
  DFFX1_LVT reg_dscratch_reg_56_ ( .D(wdata[56]), .CLK(n524), .Q(
        reg_dscratch[56]) );
  DFFX1_LVT reg_mscratch_reg_56_ ( .D(wdata[56]), .CLK(n550), .Q(
        reg_mscratch[56]) );
  DFFX1_LVT reg_sscratch_reg_56_ ( .D(wdata[56]), .CLK(n564), .Q(
        reg_sscratch[56]) );
  DFFX1_LVT u_T_41_reg_50_ ( .D(N1547), .CLK(n577), .Q(n_T_45[56]) );
  DFFX1_LVT u_T_49_reg_50_ ( .D(N1941), .CLK(n519), .Q(n1943) );
  DFFSSRX1_LVT reg_pmp_7_cfg_w_reg ( .D(wdata[56]), .SETB(1'b1), .RSTB(
        wdata[57]), .CLK(net34738), .Q(io_pmp_7_cfg_w) );
  DFFX1_LVT reg_dscratch_reg_57_ ( .D(wdata[57]), .CLK(n524), .Q(
        reg_dscratch[57]) );
  DFFX1_LVT reg_mscratch_reg_57_ ( .D(wdata[57]), .CLK(n550), .Q(
        reg_mscratch[57]) );
  DFFX1_LVT reg_sscratch_reg_57_ ( .D(wdata[57]), .CLK(n564), .Q(
        reg_sscratch[57]) );
  DFFX1_LVT u_T_41_reg_51_ ( .D(N1548), .CLK(n577), .Q(n_T_45[57]) );
  DFFX1_LVT u_T_49_reg_51_ ( .D(N1942), .CLK(n519), .Q(n1942) );
  DFFX1_LVT reg_pmp_7_cfg_x_reg ( .D(wdata[58]), .CLK(net34738), .Q(
        io_pmp_7_cfg_x) );
  DFFX1_LVT reg_dscratch_reg_58_ ( .D(wdata[58]), .CLK(n524), .Q(
        reg_dscratch[58]) );
  DFFX1_LVT reg_mscratch_reg_58_ ( .D(wdata[58]), .CLK(n550), .Q(
        reg_mscratch[58]) );
  DFFX1_LVT reg_sscratch_reg_58_ ( .D(wdata[58]), .CLK(n564), .Q(
        reg_sscratch[58]) );
  DFFX1_LVT u_T_41_reg_52_ ( .D(N1549), .CLK(n576), .Q(n_T_45[58]) );
  DFFX1_LVT u_T_49_reg_52_ ( .D(N1943), .CLK(n518), .Q(n1941) );
  DFFSSRX1_LVT reg_pmp_7_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[60]), .CLK(net34743), .Q(io_pmp_7_cfg_a[1]), .QN(n459) );
  DFFX1_LVT reg_dscratch_reg_60_ ( .D(wdata[60]), .CLK(n524), .Q(
        reg_dscratch[60]) );
  DFFX1_LVT reg_mscratch_reg_60_ ( .D(wdata[60]), .CLK(n550), .Q(
        reg_mscratch[60]) );
  DFFX1_LVT reg_sscratch_reg_60_ ( .D(wdata[60]), .CLK(n564), .Q(
        reg_sscratch[60]) );
  DFFX1_LVT reg_satp_ppn_reg_13_ ( .D(wdata[13]), .CLK(net34915), .Q(
        io_ptbr_ppn[13]) );
  DFFX1_LVT reg_satp_ppn_reg_12_ ( .D(n367), .CLK(net34915), .QN(
        io_ptbr_ppn[12]) );
  DFFX1_LVT reg_satp_ppn_reg_8_ ( .D(wdata[8]), .CLK(net34915), .Q(
        io_ptbr_ppn[8]) );
  DFFX1_LVT reg_satp_ppn_reg_7_ ( .D(wdata[7]), .CLK(net34915), .Q(
        io_ptbr_ppn[7]) );
  DFFX1_LVT reg_satp_ppn_reg_2_ ( .D(n1483), .CLK(net34915), .QN(
        io_ptbr_ppn[2]) );
  DFFX1_LVT reg_satp_ppn_reg_0_ ( .D(wdata[0]), .CLK(net34915), .Q(
        io_ptbr_ppn[0]) );
  DFFX1_LVT reg_satp_mode_reg_3_ ( .D(wdata[63]), .CLK(net34915), .Q(
        io_ptbr_mode[3]) );
  DFFX1_LVT u_T_41_reg_54_ ( .D(N1551), .CLK(n576), .Q(n_T_45[60]) );
  DFFX1_LVT u_T_49_reg_54_ ( .D(N1945), .CLK(n518), .Q(n1939) );
  DFFSSRX1_LVT reg_pmp_7_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[59]), .CLK(net34743), .Q(io_pmp_7_cfg_a[0]) );
  DFFX1_LVT reg_dscratch_reg_59_ ( .D(wdata[59]), .CLK(n524), .Q(
        reg_dscratch[59]) );
  DFFX1_LVT reg_mscratch_reg_59_ ( .D(wdata[59]), .CLK(n550), .Q(
        reg_mscratch[59]) );
  DFFX1_LVT reg_sscratch_reg_59_ ( .D(wdata[59]), .CLK(n564), .Q(
        reg_sscratch[59]) );
  DFFX1_LVT u_T_41_reg_53_ ( .D(N1550), .CLK(n576), .Q(n_T_45[59]) );
  DFFX1_LVT u_T_49_reg_53_ ( .D(N1944), .CLK(n518), .Q(n1940) );
  DFFX1_LVT reg_pmp_6_addr_reg_0_ ( .D(n_GEN_300[0]), .CLK(n535), .Q(
        io_pmp_6_addr[0]) );
  DFFX1_LVT reg_pmp_6_addr_reg_2_ ( .D(n_GEN_300[2]), .CLK(n534), .Q(
        io_pmp_6_addr[2]) );
  DFFX1_LVT reg_pmp_7_addr_reg_0_ ( .D(n_GEN_307[0]), .CLK(n533), .Q(
        io_pmp_7_addr[0]) );
  DFFX1_LVT reg_pmp_7_addr_reg_28_ ( .D(n_GEN_307[28]), .CLK(n532), .Q(
        io_pmp_7_addr[28]) );
  DFFX1_LVT reg_stvec_reg_28_ ( .D(wdata[28]), .CLK(n569), .Q(reg_stvec[28])
         );
  DFFX1_LVT reg_dscratch_reg_28_ ( .D(wdata[28]), .CLK(n523), .Q(
        reg_dscratch[28]) );
  DFFX1_LVT reg_mscratch_reg_28_ ( .D(wdata[28]), .CLK(n549), .Q(
        reg_mscratch[28]) );
  DFFX1_LVT reg_sscratch_reg_28_ ( .D(wdata[28]), .CLK(n563), .Q(
        reg_sscratch[28]) );
  DFFX1_LVT reg_bp_0_address_reg_28_ ( .D(wdata[28]), .CLK(n584), .Q(
        io_bp_0_address[28]) );
  DFFX1_LVT reg_mtval_reg_28_ ( .D(N1021), .CLK(n573), .Q(n_T_383[28]) );
  DFFSSRX1_LVT reg_mtvec_reg_28_ ( .D(n376), .SETB(wdata[28]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[28]) );
  DFFX1_LVT reg_stval_reg_28_ ( .D(N1410), .CLK(n560), .Q(n_T_444[28]) );
  DFFSSRX1_LVT reg_pmp_3_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[28]), .CLK(net35127), .Q(io_pmp_3_cfg_a[1]), .QN(n460) );
  DFFX1_LVT reg_pmp_2_addr_reg_0_ ( .D(n_GEN_272[0]), .CLK(n538), .Q(
        io_pmp_2_addr[0]) );
  DFFX1_LVT reg_pmp_2_addr_reg_23_ ( .D(n_GEN_272[23]), .CLK(n540), .Q(
        io_pmp_2_addr[23]) );
  DFFX1_LVT reg_stvec_reg_23_ ( .D(wdata[23]), .CLK(n569), .Q(reg_stvec[23])
         );
  DFFX1_LVT reg_dscratch_reg_23_ ( .D(wdata[23]), .CLK(n523), .Q(
        reg_dscratch[23]) );
  DFFX1_LVT reg_mscratch_reg_23_ ( .D(wdata[23]), .CLK(n549), .Q(
        reg_mscratch[23]) );
  DFFX1_LVT reg_sscratch_reg_23_ ( .D(wdata[23]), .CLK(n563), .Q(
        reg_sscratch[23]) );
  DFFX1_LVT reg_bp_0_address_reg_23_ ( .D(wdata[23]), .CLK(n584), .Q(
        io_bp_0_address[23]) );
  DFFX1_LVT reg_mtval_reg_23_ ( .D(N1016), .CLK(n573), .Q(n_T_383[23]) );
  DFFSSRX1_LVT reg_mtvec_reg_23_ ( .D(n376), .SETB(wdata[23]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[23]) );
  DFFX1_LVT reg_stval_reg_23_ ( .D(N1405), .CLK(n560), .Q(n_T_444[23]) );
  DFFSSRX1_LVT reg_pmp_2_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[23]), 
        .CLK(net34753), .Q(io_pmp_2_cfg_l), .QN(n441) );
  DFFSSRX1_LVT reg_pmp_2_cfg_a_reg_0_ ( .D(n503), .SETB(1'b1), .RSTB(wdata[19]), .CLK(net34753), .Q(io_pmp_2_cfg_a[0]) );
  DFFX1_LVT reg_pmp_1_addr_reg_0_ ( .D(n_GEN_265[0]), .CLK(n539), .Q(
        io_pmp_1_addr[0]) );
  DFFX1_LVT reg_pmp_1_addr_reg_15_ ( .D(n_GEN_265[15]), .CLK(n537), .Q(
        io_pmp_1_addr[15]) );
  DFFX1_LVT reg_stvec_reg_15_ ( .D(wdata[15]), .CLK(n569), .Q(reg_stvec[15])
         );
  DFFX1_LVT reg_medeleg_reg_15_ ( .D(wdata[15]), .CLK(net35172), .Q(
        read_medeleg_15) );
  DFFX1_LVT reg_dscratch_reg_15_ ( .D(wdata[15]), .CLK(n523), .Q(
        reg_dscratch[15]) );
  DFFX1_LVT reg_mscratch_reg_15_ ( .D(wdata[15]), .CLK(n549), .Q(
        reg_mscratch[15]) );
  DFFX1_LVT reg_sscratch_reg_15_ ( .D(wdata[15]), .CLK(n563), .Q(
        reg_sscratch[15]) );
  DFFX1_LVT reg_bp_0_address_reg_15_ ( .D(wdata[15]), .CLK(n585), .Q(
        io_bp_0_address[15]) );
  DFFX1_LVT reg_satp_ppn_reg_15_ ( .D(wdata[15]), .CLK(net34915), .Q(
        io_ptbr_ppn[15]) );
  DFFX1_LVT reg_mtval_reg_15_ ( .D(N1008), .CLK(n573), .Q(n_T_383[15]) );
  DFFSSRX1_LVT reg_mtvec_reg_15_ ( .D(n376), .SETB(wdata[15]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[15]) );
  DFFX1_LVT reg_stval_reg_15_ ( .D(N1397), .CLK(n560), .Q(n_T_444[15]) );
  DFFSSRX1_LVT reg_pmp_1_cfg_l_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[15]), 
        .CLK(net35132), .Q(io_pmp_1_cfg_l), .QN(n440) );
  DFFX1_LVT reg_pmp_1_cfg_r_reg ( .D(wdata[8]), .CLK(net35087), .Q(
        io_pmp_1_cfg_r) );
  DFFX1_LVT u_T_49_reg_9_ ( .D(N1900), .CLK(n518), .Q(io_time[15]) );
  DFFX1_LVT u_T_41_reg_9_ ( .D(N1506), .CLK(n576), .Q(n_T_45[15]) );
  DFFSSRX1_LVT reg_dcsr_ebreakm_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[15]), 
        .CLK(net35162), .Q(n_T_1155_3) );
  DFFX1_LVT reg_pmp_0_addr_reg_15_ ( .D(n_GEN_258[15]), .CLK(n536), .Q(
        io_pmp_0_addr[15]) );
  DFFX1_LVT reg_pmp_2_addr_reg_15_ ( .D(n_GEN_272[15]), .CLK(n535), .Q(
        io_pmp_2_addr[15]) );
  DFFX1_LVT reg_pmp_3_addr_reg_15_ ( .D(n_GEN_279[15]), .CLK(n534), .Q(
        io_pmp_3_addr[15]) );
  DFFX1_LVT reg_pmp_4_addr_reg_15_ ( .D(n_GEN_286[15]), .CLK(n533), .Q(
        io_pmp_4_addr[15]) );
  DFFX1_LVT reg_pmp_5_addr_reg_15_ ( .D(n_GEN_293[15]), .CLK(n532), .Q(
        io_pmp_5_addr[15]) );
  DFFX1_LVT reg_pmp_6_addr_reg_15_ ( .D(n_GEN_300[15]), .CLK(n538), .Q(
        io_pmp_6_addr[15]) );
  DFFX1_LVT reg_pmp_7_addr_reg_15_ ( .D(n_GEN_307[15]), .CLK(n540), .Q(
        io_pmp_7_addr[15]) );
  DFFX1_LVT reg_sepc_reg_15_ ( .D(net34835), .CLK(n581), .Q(reg_sepc[15]) );
  DFFX1_LVT reg_mepc_reg_15_ ( .D(net35037), .CLK(n545), .Q(reg_mepc[15]) );
  DFFX1_LVT reg_dpc_reg_15_ ( .D(net35259), .CLK(n528), .Q(reg_dpc[15]) );
  DFFX1_LVT reg_pmp_1_addr_reg_16_ ( .D(n_GEN_265[16]), .CLK(n539), .Q(
        io_pmp_1_addr[16]) );
  DFFX1_LVT reg_stvec_reg_16_ ( .D(wdata[16]), .CLK(n569), .Q(reg_stvec[16])
         );
  DFFX1_LVT reg_dscratch_reg_16_ ( .D(wdata[16]), .CLK(n523), .Q(
        reg_dscratch[16]) );
  DFFX1_LVT reg_pmp_2_cfg_r_reg ( .D(wdata[16]), .CLK(net34748), .Q(
        io_pmp_2_cfg_r) );
  DFFX1_LVT reg_mscratch_reg_16_ ( .D(wdata[16]), .CLK(n549), .Q(
        reg_mscratch[16]) );
  DFFX1_LVT reg_sscratch_reg_16_ ( .D(wdata[16]), .CLK(n563), .Q(
        reg_sscratch[16]) );
  DFFX1_LVT reg_bp_0_address_reg_16_ ( .D(wdata[16]), .CLK(n585), .Q(
        io_bp_0_address[16]) );
  DFFX1_LVT reg_satp_ppn_reg_16_ ( .D(wdata[16]), .CLK(net34915), .Q(
        io_ptbr_ppn[16]) );
  DFFX1_LVT reg_mtval_reg_16_ ( .D(N1009), .CLK(n573), .Q(n_T_383[16]) );
  DFFSSRX1_LVT reg_mtvec_reg_16_ ( .D(n378), .SETB(wdata[16]), .RSTB(1'b1), 
        .CLK(n554), .QN(reg_mtvec[16]) );
  DFFX1_LVT reg_stval_reg_16_ ( .D(N1398), .CLK(n560), .Q(n_T_444[16]) );
  DFFX1_LVT u_T_41_reg_10_ ( .D(N1507), .CLK(n576), .Q(n_T_45[16]) );
  DFFX1_LVT u_T_49_reg_10_ ( .D(N1901), .CLK(n518), .Q(io_time[16]) );
  DFFX1_LVT reg_pmp_0_addr_reg_16_ ( .D(n_GEN_258[16]), .CLK(n537), .Q(
        io_pmp_0_addr[16]) );
  DFFX1_LVT reg_pmp_2_addr_reg_16_ ( .D(n_GEN_272[16]), .CLK(n536), .Q(
        io_pmp_2_addr[16]) );
  DFFX1_LVT reg_pmp_3_addr_reg_16_ ( .D(n_GEN_279[16]), .CLK(n535), .Q(
        io_pmp_3_addr[16]) );
  DFFX1_LVT reg_pmp_4_addr_reg_16_ ( .D(n_GEN_286[16]), .CLK(n534), .Q(
        io_pmp_4_addr[16]) );
  DFFX1_LVT reg_pmp_5_addr_reg_16_ ( .D(n_GEN_293[16]), .CLK(n533), .Q(
        io_pmp_5_addr[16]) );
  DFFX1_LVT reg_pmp_6_addr_reg_16_ ( .D(n_GEN_300[16]), .CLK(n532), .Q(
        io_pmp_6_addr[16]) );
  DFFX1_LVT reg_pmp_7_addr_reg_16_ ( .D(n_GEN_307[16]), .CLK(n538), .Q(
        io_pmp_7_addr[16]) );
  DFFX1_LVT reg_sepc_reg_16_ ( .D(net34832), .CLK(n582), .Q(reg_sepc[16]) );
  DFFX1_LVT reg_mepc_reg_16_ ( .D(net35034), .CLK(n546), .Q(reg_mepc[16]) );
  DFFX1_LVT reg_dpc_reg_16_ ( .D(net35256), .CLK(n529), .Q(reg_dpc[16]) );
  DFFX1_LVT reg_pmp_1_addr_reg_17_ ( .D(n_GEN_265[17]), .CLK(n540), .Q(
        io_pmp_1_addr[17]) );
  DFFX1_LVT reg_stvec_reg_17_ ( .D(wdata[17]), .CLK(n569), .Q(reg_stvec[17])
         );
  DFFX1_LVT reg_dscratch_reg_17_ ( .D(wdata[17]), .CLK(n523), .Q(
        reg_dscratch[17]) );
  DFFX1_LVT reg_mscratch_reg_17_ ( .D(wdata[17]), .CLK(n549), .Q(
        reg_mscratch[17]) );
  DFFX1_LVT reg_sscratch_reg_17_ ( .D(wdata[17]), .CLK(n563), .Q(
        reg_sscratch[17]) );
  DFFX1_LVT reg_bp_0_address_reg_17_ ( .D(wdata[17]), .CLK(n585), .Q(
        io_bp_0_address[17]) );
  DFFX1_LVT reg_satp_ppn_reg_17_ ( .D(wdata[17]), .CLK(net34915), .Q(
        io_ptbr_ppn[17]) );
  DFFX1_LVT reg_mtval_reg_17_ ( .D(N1010), .CLK(n573), .Q(n_T_383[17]) );
  DFFSSRX1_LVT reg_mtvec_reg_17_ ( .D(n378), .SETB(wdata[17]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[17]) );
  DFFX1_LVT reg_stval_reg_17_ ( .D(N1399), .CLK(n560), .Q(n_T_444[17]) );
  DFFSSRX1_LVT reg_mstatus_mprv_reg ( .D(n503), .SETB(1'b1), .RSTB(wdata[17]), 
        .CLK(net35152), .Q(n1927) );
  DFFX1_LVT u_T_41_reg_11_ ( .D(N1508), .CLK(n576), .Q(n_T_45[17]) );
  DFFX1_LVT u_T_49_reg_11_ ( .D(N1902), .CLK(n518), .Q(io_time[17]) );
  DFFX1_LVT reg_pmp_0_addr_reg_17_ ( .D(n_GEN_258[17]), .CLK(n539), .Q(
        io_pmp_0_addr[17]) );
  DFFX1_LVT reg_pmp_2_addr_reg_17_ ( .D(n_GEN_272[17]), .CLK(n537), .Q(
        io_pmp_2_addr[17]) );
  DFFX1_LVT reg_pmp_3_addr_reg_17_ ( .D(n_GEN_279[17]), .CLK(n536), .Q(
        io_pmp_3_addr[17]) );
  DFFX1_LVT reg_pmp_4_addr_reg_17_ ( .D(n_GEN_286[17]), .CLK(n535), .Q(
        io_pmp_4_addr[17]) );
  DFFX1_LVT reg_pmp_5_addr_reg_17_ ( .D(n_GEN_293[17]), .CLK(n531), .Q(
        io_pmp_5_addr[17]) );
  DFFX1_LVT reg_pmp_6_addr_reg_17_ ( .D(n_GEN_300[17]), .CLK(n531), .Q(
        io_pmp_6_addr[17]) );
  DFFX1_LVT reg_pmp_7_addr_reg_17_ ( .D(n_GEN_307[17]), .CLK(n531), .Q(
        io_pmp_7_addr[17]) );
  DFFSSRX1_LVT reg_pmp_2_cfg_w_reg ( .D(wdata[17]), .SETB(1'b1), .RSTB(
        wdata[16]), .CLK(net34748), .Q(io_pmp_2_cfg_w) );
  DFFX1_LVT reg_sepc_reg_17_ ( .D(net34829), .CLK(n582), .Q(reg_sepc[17]) );
  DFFX1_LVT reg_mepc_reg_17_ ( .D(net35031), .CLK(n546), .Q(reg_mepc[17]) );
  DFFX1_LVT reg_dpc_reg_17_ ( .D(net35253), .CLK(n529), .Q(reg_dpc[17]) );
  DFFX1_LVT reg_pmp_1_addr_reg_18_ ( .D(n_GEN_265[18]), .CLK(n531), .Q(
        io_pmp_1_addr[18]) );
  DFFX1_LVT reg_stvec_reg_18_ ( .D(wdata[18]), .CLK(n569), .Q(reg_stvec[18])
         );
  DFFX1_LVT reg_dscratch_reg_18_ ( .D(wdata[18]), .CLK(n523), .Q(
        reg_dscratch[18]) );
  DFFX1_LVT reg_pmp_2_cfg_x_reg ( .D(wdata[18]), .CLK(net34748), .Q(
        io_pmp_2_cfg_x) );
  DFFX1_LVT reg_mscratch_reg_18_ ( .D(wdata[18]), .CLK(n549), .Q(
        reg_mscratch[18]) );
  DFFX1_LVT reg_sscratch_reg_18_ ( .D(wdata[18]), .CLK(n563), .Q(
        reg_sscratch[18]) );
  DFFX1_LVT reg_bp_0_address_reg_18_ ( .D(wdata[18]), .CLK(n585), .Q(
        io_bp_0_address[18]) );
  DFFX1_LVT reg_satp_ppn_reg_18_ ( .D(wdata[18]), .CLK(net34915), .Q(
        io_ptbr_ppn[18]) );
  DFFX1_LVT reg_mtval_reg_18_ ( .D(N1011), .CLK(n573), .Q(n_T_383[18]) );
  DFFSSRX1_LVT reg_mtvec_reg_18_ ( .D(n378), .SETB(wdata[18]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[18]) );
  DFFX1_LVT reg_stval_reg_18_ ( .D(N1400), .CLK(n560), .Q(n_T_444[18]) );
  DFFSSRX1_LVT reg_mstatus_sum_reg ( .D(n503), .SETB(1'b1), .RSTB(wdata[18]), 
        .CLK(net35157), .Q(io_status_sum) );
  DFFX1_LVT u_T_41_reg_12_ ( .D(N1509), .CLK(n576), .Q(n_T_45[18]) );
  DFFX1_LVT u_T_49_reg_12_ ( .D(N1903), .CLK(n518), .Q(io_time[18]) );
  DFFX1_LVT reg_pmp_0_addr_reg_18_ ( .D(n_GEN_258[18]), .CLK(n531), .Q(
        io_pmp_0_addr[18]) );
  DFFX1_LVT reg_pmp_2_addr_reg_18_ ( .D(n_GEN_272[18]), .CLK(n531), .Q(
        io_pmp_2_addr[18]) );
  DFFX1_LVT reg_pmp_3_addr_reg_18_ ( .D(n_GEN_279[18]), .CLK(n531), .Q(
        io_pmp_3_addr[18]) );
  DFFX1_LVT reg_pmp_4_addr_reg_18_ ( .D(n_GEN_286[18]), .CLK(n531), .Q(
        io_pmp_4_addr[18]) );
  DFFX1_LVT reg_pmp_5_addr_reg_18_ ( .D(n_GEN_293[18]), .CLK(n531), .Q(
        io_pmp_5_addr[18]) );
  DFFX1_LVT reg_pmp_6_addr_reg_18_ ( .D(n_GEN_300[18]), .CLK(n531), .Q(
        io_pmp_6_addr[18]) );
  DFFX1_LVT reg_pmp_7_addr_reg_18_ ( .D(n_GEN_307[18]), .CLK(n531), .Q(
        io_pmp_7_addr[18]) );
  DFFX1_LVT reg_sepc_reg_18_ ( .D(net34826), .CLK(n582), .Q(reg_sepc[18]) );
  DFFX1_LVT reg_mepc_reg_18_ ( .D(net35028), .CLK(n546), .Q(reg_mepc[18]) );
  DFFX1_LVT reg_dpc_reg_18_ ( .D(net35250), .CLK(n529), .Q(reg_dpc[18]) );
  DFFX1_LVT reg_pmp_1_addr_reg_19_ ( .D(n_GEN_265[19]), .CLK(n531), .Q(
        io_pmp_1_addr[19]) );
  DFFX1_LVT reg_stvec_reg_19_ ( .D(wdata[19]), .CLK(n569), .Q(reg_stvec[19])
         );
  DFFX1_LVT reg_dscratch_reg_19_ ( .D(wdata[19]), .CLK(n523), .Q(
        reg_dscratch[19]) );
  DFFX1_LVT reg_mscratch_reg_19_ ( .D(wdata[19]), .CLK(n549), .Q(
        reg_mscratch[19]) );
  DFFX1_LVT reg_sscratch_reg_19_ ( .D(wdata[19]), .CLK(n563), .Q(
        reg_sscratch[19]) );
  DFFX1_LVT reg_bp_0_address_reg_19_ ( .D(wdata[19]), .CLK(n585), .Q(
        io_bp_0_address[19]) );
  DFFX1_LVT reg_satp_ppn_reg_19_ ( .D(wdata[19]), .CLK(net34915), .Q(
        io_ptbr_ppn[19]) );
  DFFX1_LVT reg_mtval_reg_19_ ( .D(N1012), .CLK(n573), .Q(n_T_383[19]) );
  DFFSSRX1_LVT reg_mtvec_reg_19_ ( .D(n378), .SETB(wdata[19]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[19]) );
  DFFX1_LVT reg_stval_reg_19_ ( .D(N1401), .CLK(n560), .Q(n_T_444[19]) );
  DFFX1_LVT u_T_49_reg_13_ ( .D(N1904), .CLK(n518), .Q(io_time[19]) );
  DFFX1_LVT u_T_41_reg_13_ ( .D(N1510), .CLK(n576), .Q(n_T_45[19]) );
  DFFSSRX1_LVT reg_mstatus_mxr_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[19]), 
        .CLK(net35157), .Q(io_status_mxr) );
  DFFX1_LVT reg_pmp_0_addr_reg_19_ ( .D(n_GEN_258[19]), .CLK(n544), .Q(
        io_pmp_0_addr[19]) );
  DFFX1_LVT reg_pmp_2_addr_reg_19_ ( .D(n_GEN_272[19]), .CLK(n544), .Q(
        io_pmp_2_addr[19]) );
  DFFX1_LVT reg_pmp_3_addr_reg_19_ ( .D(n_GEN_279[19]), .CLK(n544), .Q(
        io_pmp_3_addr[19]) );
  DFFX1_LVT reg_pmp_4_addr_reg_19_ ( .D(n_GEN_286[19]), .CLK(n544), .Q(
        io_pmp_4_addr[19]) );
  DFFX1_LVT reg_pmp_5_addr_reg_19_ ( .D(n_GEN_293[19]), .CLK(n544), .Q(
        io_pmp_5_addr[19]) );
  DFFX1_LVT reg_pmp_6_addr_reg_19_ ( .D(n_GEN_300[19]), .CLK(n544), .Q(
        io_pmp_6_addr[19]) );
  DFFX1_LVT reg_pmp_7_addr_reg_19_ ( .D(n_GEN_307[19]), .CLK(n544), .Q(
        io_pmp_7_addr[19]) );
  DFFX1_LVT reg_sepc_reg_19_ ( .D(net34823), .CLK(n582), .Q(reg_sepc[19]) );
  DFFX1_LVT reg_mepc_reg_19_ ( .D(net35025), .CLK(n546), .Q(reg_mepc[19]) );
  DFFX1_LVT reg_dpc_reg_19_ ( .D(net35247), .CLK(n529), .Q(reg_dpc[19]) );
  DFFX1_LVT reg_pmp_1_addr_reg_20_ ( .D(n_GEN_265[20]), .CLK(n544), .Q(
        io_pmp_1_addr[20]) );
  DFFX1_LVT reg_stvec_reg_20_ ( .D(wdata[20]), .CLK(n569), .Q(reg_stvec[20])
         );
  DFFX1_LVT reg_dscratch_reg_20_ ( .D(wdata[20]), .CLK(n523), .Q(
        reg_dscratch[20]) );
  DFFX1_LVT reg_mscratch_reg_20_ ( .D(wdata[20]), .CLK(n549), .Q(
        reg_mscratch[20]) );
  DFFX1_LVT reg_sscratch_reg_20_ ( .D(wdata[20]), .CLK(n563), .Q(
        reg_sscratch[20]) );
  DFFX1_LVT reg_bp_0_address_reg_20_ ( .D(wdata[20]), .CLK(n585), .Q(
        io_bp_0_address[20]) );
  DFFX1_LVT reg_mtval_reg_20_ ( .D(N1013), .CLK(n573), .Q(n_T_383[20]) );
  DFFSSRX1_LVT reg_mtvec_reg_20_ ( .D(n378), .SETB(wdata[20]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[20]) );
  DFFX1_LVT reg_stval_reg_20_ ( .D(N1402), .CLK(n560), .Q(n_T_444[20]) );
  DFFSSRX1_LVT reg_pmp_2_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[20]), .CLK(net34753), .Q(io_pmp_2_cfg_a[1]), .QN(n463) );
  DFFX1_LVT u_T_49_reg_14_ ( .D(N1905), .CLK(n518), .Q(io_time[20]) );
  DFFX1_LVT u_T_41_reg_14_ ( .D(N1511), .CLK(n576), .Q(n_T_45[20]) );
  DFFSSRX1_LVT reg_mstatus_tvm_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[20]), 
        .CLK(net35152), .Q(n1926), .QN(n447) );
  DFFX1_LVT reg_pmp_0_addr_reg_20_ ( .D(n_GEN_258[20]), .CLK(n544), .Q(
        io_pmp_0_addr[20]) );
  DFFX1_LVT reg_pmp_2_addr_reg_20_ ( .D(n_GEN_272[20]), .CLK(n544), .Q(
        io_pmp_2_addr[20]) );
  DFFX1_LVT reg_pmp_3_addr_reg_20_ ( .D(n_GEN_279[20]), .CLK(n544), .Q(
        io_pmp_3_addr[20]) );
  DFFX1_LVT reg_pmp_4_addr_reg_20_ ( .D(n_GEN_286[20]), .CLK(n544), .Q(
        io_pmp_4_addr[20]) );
  DFFX1_LVT reg_pmp_5_addr_reg_20_ ( .D(n_GEN_293[20]), .CLK(n543), .Q(
        io_pmp_5_addr[20]) );
  DFFX1_LVT reg_pmp_6_addr_reg_20_ ( .D(n_GEN_300[20]), .CLK(n543), .Q(
        io_pmp_6_addr[20]) );
  DFFX1_LVT reg_pmp_7_addr_reg_20_ ( .D(n_GEN_307[20]), .CLK(n543), .Q(
        io_pmp_7_addr[20]) );
  DFFX1_LVT reg_sepc_reg_20_ ( .D(net34820), .CLK(n582), .Q(reg_sepc[20]) );
  DFFX1_LVT reg_mepc_reg_20_ ( .D(net35022), .CLK(n546), .Q(reg_mepc[20]) );
  DFFX1_LVT reg_dpc_reg_20_ ( .D(net35244), .CLK(n529), .Q(reg_dpc[20]) );
  DFFX1_LVT reg_pmp_1_addr_reg_21_ ( .D(n_GEN_265[21]), .CLK(n543), .Q(
        io_pmp_1_addr[21]) );
  DFFX1_LVT reg_stvec_reg_21_ ( .D(wdata[21]), .CLK(n570), .Q(reg_stvec[21])
         );
  DFFX1_LVT reg_dscratch_reg_21_ ( .D(wdata[21]), .CLK(n523), .Q(
        reg_dscratch[21]) );
  DFFX1_LVT reg_mscratch_reg_21_ ( .D(wdata[21]), .CLK(n549), .Q(
        reg_mscratch[21]) );
  DFFX1_LVT reg_sscratch_reg_21_ ( .D(wdata[21]), .CLK(n563), .Q(
        reg_sscratch[21]) );
  DFFX1_LVT reg_bp_0_address_reg_21_ ( .D(wdata[21]), .CLK(n585), .Q(
        io_bp_0_address[21]) );
  DFFX1_LVT reg_mtval_reg_21_ ( .D(N1014), .CLK(n574), .Q(n_T_383[21]) );
  DFFSSRX1_LVT reg_mtvec_reg_21_ ( .D(n378), .SETB(wdata[21]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[21]) );
  DFFX1_LVT reg_stval_reg_21_ ( .D(N1403), .CLK(n561), .Q(n_T_444[21]) );
  DFFSSRX1_LVT reg_mstatus_tw_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[21]), 
        .CLK(net35152), .Q(n1925) );
  DFFX1_LVT u_T_41_reg_15_ ( .D(N1512), .CLK(n576), .Q(n_T_45[21]) );
  DFFX1_LVT u_T_49_reg_15_ ( .D(N1906), .CLK(n518), .Q(io_time[21]) );
  DFFX1_LVT reg_pmp_0_addr_reg_21_ ( .D(n_GEN_258[21]), .CLK(n543), .Q(
        io_pmp_0_addr[21]) );
  DFFX1_LVT reg_pmp_2_addr_reg_21_ ( .D(n_GEN_272[21]), .CLK(n543), .Q(
        io_pmp_2_addr[21]) );
  DFFX1_LVT reg_pmp_3_addr_reg_21_ ( .D(n_GEN_279[21]), .CLK(n543), .Q(
        io_pmp_3_addr[21]) );
  DFFX1_LVT reg_pmp_4_addr_reg_21_ ( .D(n_GEN_286[21]), .CLK(n543), .Q(
        io_pmp_4_addr[21]) );
  DFFX1_LVT reg_pmp_5_addr_reg_21_ ( .D(n_GEN_293[21]), .CLK(n543), .Q(
        io_pmp_5_addr[21]) );
  DFFX1_LVT reg_pmp_6_addr_reg_21_ ( .D(n_GEN_300[21]), .CLK(n543), .Q(
        io_pmp_6_addr[21]) );
  DFFX1_LVT reg_pmp_7_addr_reg_21_ ( .D(n_GEN_307[21]), .CLK(n543), .Q(
        io_pmp_7_addr[21]) );
  DFFX1_LVT reg_sepc_reg_21_ ( .D(net34817), .CLK(n582), .Q(reg_sepc[21]) );
  DFFX1_LVT reg_mepc_reg_21_ ( .D(net35019), .CLK(n546), .Q(reg_mepc[21]) );
  DFFX1_LVT reg_dpc_reg_21_ ( .D(net35241), .CLK(n529), .Q(reg_dpc[21]) );
  DFFX1_LVT reg_pmp_1_addr_reg_22_ ( .D(n_GEN_265[22]), .CLK(n543), .Q(
        io_pmp_1_addr[22]) );
  DFFX1_LVT reg_stvec_reg_22_ ( .D(wdata[22]), .CLK(n570), .Q(reg_stvec[22])
         );
  DFFX1_LVT reg_dscratch_reg_22_ ( .D(wdata[22]), .CLK(n523), .Q(
        reg_dscratch[22]) );
  DFFX1_LVT reg_mscratch_reg_22_ ( .D(wdata[22]), .CLK(n549), .Q(
        reg_mscratch[22]) );
  DFFX1_LVT reg_sscratch_reg_22_ ( .D(wdata[22]), .CLK(n563), .Q(
        reg_sscratch[22]) );
  DFFX1_LVT reg_bp_0_address_reg_22_ ( .D(wdata[22]), .CLK(n585), .Q(
        io_bp_0_address[22]) );
  DFFX1_LVT reg_mtval_reg_22_ ( .D(N1015), .CLK(n574), .Q(n_T_383[22]) );
  DFFSSRX1_LVT reg_mtvec_reg_22_ ( .D(n378), .SETB(wdata[22]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[22]) );
  DFFX1_LVT reg_stval_reg_22_ ( .D(N1404), .CLK(n561), .Q(n_T_444[22]) );
  DFFSSRX1_LVT reg_mstatus_tsr_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[22]), 
        .CLK(net35152), .Q(n1924) );
  DFFX1_LVT u_T_41_reg_16_ ( .D(N1513), .CLK(n576), .Q(n_T_45[22]) );
  DFFX1_LVT u_T_49_reg_16_ ( .D(N1907), .CLK(n518), .Q(io_time[22]) );
  DFFX1_LVT reg_pmp_0_addr_reg_22_ ( .D(n_GEN_258[22]), .CLK(n534), .Q(
        io_pmp_0_addr[22]) );
  DFFX1_LVT reg_pmp_2_addr_reg_22_ ( .D(n_GEN_272[22]), .CLK(n533), .Q(
        io_pmp_2_addr[22]) );
  DFFX1_LVT reg_pmp_3_addr_reg_22_ ( .D(n_GEN_279[22]), .CLK(n532), .Q(
        io_pmp_3_addr[22]) );
  DFFX1_LVT reg_pmp_4_addr_reg_22_ ( .D(n_GEN_286[22]), .CLK(n538), .Q(
        io_pmp_4_addr[22]) );
  DFFX1_LVT reg_pmp_5_addr_reg_22_ ( .D(n_GEN_293[22]), .CLK(n540), .Q(
        io_pmp_5_addr[22]) );
  DFFX1_LVT reg_pmp_6_addr_reg_22_ ( .D(n_GEN_300[22]), .CLK(n539), .Q(
        io_pmp_6_addr[22]) );
  DFFX1_LVT reg_pmp_7_addr_reg_22_ ( .D(n_GEN_307[22]), .CLK(n537), .Q(
        io_pmp_7_addr[22]) );
  DFFX1_LVT reg_sepc_reg_22_ ( .D(net34814), .CLK(n582), .Q(reg_sepc[22]) );
  DFFX1_LVT reg_mepc_reg_22_ ( .D(net35016), .CLK(n546), .Q(reg_mepc[22]) );
  DFFX1_LVT reg_dpc_reg_22_ ( .D(net35238), .CLK(n529), .Q(reg_dpc[22]) );
  DFFX1_LVT reg_pmp_1_addr_reg_2_ ( .D(n_GEN_265[2]), .CLK(n536), .Q(
        io_pmp_1_addr[2]) );
  DFFX1_LVT u_T_41_reg_17_ ( .D(N1514), .CLK(n576), .Q(n_T_45[23]) );
  DFFX1_LVT u_T_49_reg_17_ ( .D(N1908), .CLK(n518), .Q(io_time[23]) );
  DFFX1_LVT reg_pmp_0_addr_reg_23_ ( .D(n_GEN_258[23]), .CLK(n535), .Q(
        io_pmp_0_addr[23]) );
  DFFX1_LVT reg_pmp_1_addr_reg_23_ ( .D(n_GEN_265[23]), .CLK(n534), .Q(
        io_pmp_1_addr[23]) );
  DFFX1_LVT reg_pmp_3_addr_reg_23_ ( .D(n_GEN_279[23]), .CLK(n533), .Q(
        io_pmp_3_addr[23]) );
  DFFX1_LVT reg_pmp_4_addr_reg_23_ ( .D(n_GEN_286[23]), .CLK(n532), .Q(
        io_pmp_4_addr[23]) );
  DFFX1_LVT reg_pmp_5_addr_reg_23_ ( .D(n_GEN_293[23]), .CLK(n542), .Q(
        io_pmp_5_addr[23]) );
  DFFX1_LVT reg_pmp_6_addr_reg_23_ ( .D(n_GEN_300[23]), .CLK(n542), .Q(
        io_pmp_6_addr[23]) );
  DFFX1_LVT reg_pmp_7_addr_reg_23_ ( .D(n_GEN_307[23]), .CLK(n542), .Q(
        io_pmp_7_addr[23]) );
  DFFX1_LVT reg_sepc_reg_23_ ( .D(net34811), .CLK(n582), .Q(reg_sepc[23]) );
  DFFX1_LVT reg_mepc_reg_23_ ( .D(net35013), .CLK(n546), .Q(reg_mepc[23]) );
  DFFX1_LVT reg_dpc_reg_23_ ( .D(net35235), .CLK(n529), .Q(reg_dpc[23]) );
  DFFX1_LVT reg_pmp_2_addr_reg_24_ ( .D(n_GEN_272[24]), .CLK(n542), .Q(
        io_pmp_2_addr[24]) );
  DFFX1_LVT reg_stvec_reg_24_ ( .D(wdata[24]), .CLK(n570), .Q(reg_stvec[24])
         );
  DFFX1_LVT reg_dscratch_reg_24_ ( .D(wdata[24]), .CLK(n523), .Q(
        reg_dscratch[24]) );
  DFFX1_LVT reg_pmp_3_cfg_r_reg ( .D(wdata[24]), .CLK(net35122), .Q(
        io_pmp_3_cfg_r) );
  DFFX1_LVT reg_mscratch_reg_24_ ( .D(wdata[24]), .CLK(n549), .Q(
        reg_mscratch[24]) );
  DFFX1_LVT reg_sscratch_reg_24_ ( .D(wdata[24]), .CLK(n563), .Q(
        reg_sscratch[24]) );
  DFFX1_LVT reg_bp_0_address_reg_24_ ( .D(wdata[24]), .CLK(n585), .Q(
        io_bp_0_address[24]) );
  DFFX1_LVT reg_mtval_reg_24_ ( .D(N1017), .CLK(n574), .Q(n_T_383[24]) );
  DFFSSRX1_LVT reg_mtvec_reg_24_ ( .D(n378), .SETB(wdata[24]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[24]) );
  DFFX1_LVT reg_stval_reg_24_ ( .D(N1406), .CLK(n561), .Q(n_T_444[24]) );
  DFFX1_LVT u_T_41_reg_18_ ( .D(N1515), .CLK(n575), .Q(n_T_45[24]) );
  DFFX1_LVT u_T_49_reg_18_ ( .D(N1909), .CLK(n517), .Q(io_time[24]) );
  DFFX1_LVT reg_pmp_0_addr_reg_24_ ( .D(n_GEN_258[24]), .CLK(n542), .Q(
        io_pmp_0_addr[24]) );
  DFFX1_LVT reg_pmp_1_addr_reg_24_ ( .D(n_GEN_265[24]), .CLK(n542), .Q(
        io_pmp_1_addr[24]) );
  DFFX1_LVT reg_pmp_3_addr_reg_24_ ( .D(n_GEN_279[24]), .CLK(n542), .Q(
        io_pmp_3_addr[24]) );
  DFFX1_LVT reg_pmp_4_addr_reg_24_ ( .D(n_GEN_286[24]), .CLK(n542), .Q(
        io_pmp_4_addr[24]) );
  DFFX1_LVT reg_pmp_5_addr_reg_24_ ( .D(n_GEN_293[24]), .CLK(n542), .Q(
        io_pmp_5_addr[24]) );
  DFFX1_LVT reg_pmp_6_addr_reg_24_ ( .D(n_GEN_300[24]), .CLK(n542), .Q(
        io_pmp_6_addr[24]) );
  DFFX1_LVT reg_pmp_7_addr_reg_24_ ( .D(n_GEN_307[24]), .CLK(n542), .Q(
        io_pmp_7_addr[24]) );
  DFFX1_LVT reg_sepc_reg_24_ ( .D(net34808), .CLK(n582), .Q(reg_sepc[24]) );
  DFFX1_LVT reg_mepc_reg_24_ ( .D(net35010), .CLK(n546), .Q(reg_mepc[24]) );
  DFFX1_LVT reg_dpc_reg_24_ ( .D(net35232), .CLK(n529), .Q(reg_dpc[24]) );
  DFFX1_LVT reg_pmp_2_addr_reg_25_ ( .D(n_GEN_272[25]), .CLK(n542), .Q(
        io_pmp_2_addr[25]) );
  DFFX1_LVT reg_stvec_reg_25_ ( .D(wdata[25]), .CLK(n570), .Q(reg_stvec[25])
         );
  DFFX1_LVT reg_dscratch_reg_25_ ( .D(wdata[25]), .CLK(n523), .Q(
        reg_dscratch[25]) );
  DFFX1_LVT reg_mscratch_reg_25_ ( .D(wdata[25]), .CLK(n549), .Q(
        reg_mscratch[25]) );
  DFFX1_LVT reg_sscratch_reg_25_ ( .D(wdata[25]), .CLK(n563), .Q(
        reg_sscratch[25]) );
  DFFX1_LVT reg_bp_0_address_reg_25_ ( .D(wdata[25]), .CLK(n585), .Q(
        io_bp_0_address[25]) );
  DFFX1_LVT reg_mtval_reg_25_ ( .D(N1018), .CLK(n574), .Q(n_T_383[25]) );
  DFFSSRX1_LVT reg_mtvec_reg_25_ ( .D(n378), .SETB(wdata[25]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[25]) );
  DFFX1_LVT reg_stval_reg_25_ ( .D(N1407), .CLK(n561), .Q(n_T_444[25]) );
  DFFX1_LVT u_T_41_reg_19_ ( .D(N1516), .CLK(n575), .Q(n_T_45[25]) );
  DFFX1_LVT u_T_49_reg_19_ ( .D(N1910), .CLK(n517), .Q(io_time[25]) );
  DFFX1_LVT reg_pmp_0_addr_reg_25_ ( .D(n_GEN_258[25]), .CLK(n541), .Q(
        io_pmp_0_addr[25]) );
  DFFX1_LVT reg_pmp_1_addr_reg_25_ ( .D(n_GEN_265[25]), .CLK(n541), .Q(
        io_pmp_1_addr[25]) );
  DFFX1_LVT reg_pmp_3_addr_reg_25_ ( .D(n_GEN_279[25]), .CLK(n541), .Q(
        io_pmp_3_addr[25]) );
  DFFX1_LVT reg_pmp_4_addr_reg_25_ ( .D(n_GEN_286[25]), .CLK(n541), .Q(
        io_pmp_4_addr[25]) );
  DFFX1_LVT reg_pmp_5_addr_reg_25_ ( .D(n_GEN_293[25]), .CLK(n541), .Q(
        io_pmp_5_addr[25]) );
  DFFX1_LVT reg_pmp_6_addr_reg_25_ ( .D(n_GEN_300[25]), .CLK(n541), .Q(
        io_pmp_6_addr[25]) );
  DFFX1_LVT reg_pmp_7_addr_reg_25_ ( .D(n_GEN_307[25]), .CLK(n541), .Q(
        io_pmp_7_addr[25]) );
  DFFSSRX1_LVT reg_pmp_3_cfg_w_reg ( .D(wdata[24]), .SETB(1'b1), .RSTB(
        wdata[25]), .CLK(net35122), .Q(io_pmp_3_cfg_w) );
  DFFX1_LVT reg_sepc_reg_25_ ( .D(net34805), .CLK(n582), .Q(reg_sepc[25]) );
  DFFX1_LVT reg_mepc_reg_25_ ( .D(net35007), .CLK(n546), .Q(reg_mepc[25]) );
  DFFX1_LVT reg_dpc_reg_25_ ( .D(net35229), .CLK(n529), .Q(reg_dpc[25]) );
  DFFX1_LVT reg_pmp_2_addr_reg_26_ ( .D(n_GEN_272[26]), .CLK(n541), .Q(
        io_pmp_2_addr[26]) );
  DFFX1_LVT reg_stvec_reg_26_ ( .D(wdata[26]), .CLK(n570), .Q(reg_stvec[26])
         );
  DFFX1_LVT reg_dscratch_reg_26_ ( .D(wdata[26]), .CLK(n522), .Q(
        reg_dscratch[26]) );
  DFFX1_LVT reg_pmp_3_cfg_x_reg ( .D(wdata[26]), .CLK(net35122), .Q(
        io_pmp_3_cfg_x) );
  DFFX1_LVT reg_mscratch_reg_26_ ( .D(wdata[26]), .CLK(n548), .Q(
        reg_mscratch[26]) );
  DFFX1_LVT reg_sscratch_reg_26_ ( .D(wdata[26]), .CLK(n562), .Q(
        reg_sscratch[26]) );
  DFFX1_LVT reg_bp_0_address_reg_26_ ( .D(wdata[26]), .CLK(n585), .Q(
        io_bp_0_address[26]) );
  DFFX1_LVT reg_mtval_reg_26_ ( .D(N1019), .CLK(n574), .Q(n_T_383[26]) );
  DFFSSRX1_LVT reg_mtvec_reg_26_ ( .D(n378), .SETB(wdata[26]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[26]) );
  DFFX1_LVT reg_stval_reg_26_ ( .D(N1408), .CLK(n561), .Q(n_T_444[26]) );
  DFFX1_LVT u_T_41_reg_20_ ( .D(N1517), .CLK(n575), .Q(n_T_45[26]) );
  DFFX1_LVT u_T_49_reg_20_ ( .D(N1911), .CLK(n517), .Q(io_time[26]) );
  DFFX1_LVT reg_pmp_0_addr_reg_26_ ( .D(n_GEN_258[26]), .CLK(n541), .Q(
        io_pmp_0_addr[26]) );
  DFFX1_LVT reg_pmp_1_addr_reg_26_ ( .D(n_GEN_265[26]), .CLK(n541), .Q(
        io_pmp_1_addr[26]) );
  DFFX1_LVT reg_pmp_3_addr_reg_26_ ( .D(n_GEN_279[26]), .CLK(n541), .Q(
        io_pmp_3_addr[26]) );
  DFFX1_LVT reg_pmp_4_addr_reg_26_ ( .D(n_GEN_286[26]), .CLK(n541), .Q(
        io_pmp_4_addr[26]) );
  DFFX1_LVT reg_pmp_5_addr_reg_26_ ( .D(n_GEN_293[26]), .CLK(n538), .Q(
        io_pmp_5_addr[26]) );
  DFFX1_LVT reg_pmp_6_addr_reg_26_ ( .D(n_GEN_300[26]), .CLK(n540), .Q(
        io_pmp_6_addr[26]) );
  DFFX1_LVT reg_pmp_7_addr_reg_26_ ( .D(n_GEN_307[26]), .CLK(n540), .Q(
        io_pmp_7_addr[26]) );
  DFFX1_LVT reg_sepc_reg_26_ ( .D(net34802), .CLK(n582), .Q(reg_sepc[26]) );
  DFFX1_LVT reg_mepc_reg_26_ ( .D(net35004), .CLK(n546), .Q(reg_mepc[26]) );
  DFFX1_LVT reg_dpc_reg_26_ ( .D(net35226), .CLK(n529), .Q(reg_dpc[26]) );
  DFFX1_LVT reg_pmp_2_addr_reg_27_ ( .D(n_GEN_272[27]), .CLK(n539), .Q(
        io_pmp_2_addr[27]) );
  DFFX1_LVT reg_stvec_reg_27_ ( .D(wdata[27]), .CLK(n570), .Q(reg_stvec[27])
         );
  DFFX1_LVT reg_dscratch_reg_27_ ( .D(wdata[27]), .CLK(n522), .Q(
        reg_dscratch[27]) );
  DFFX1_LVT reg_mscratch_reg_27_ ( .D(wdata[27]), .CLK(n548), .Q(
        reg_mscratch[27]) );
  DFFX1_LVT reg_sscratch_reg_27_ ( .D(wdata[27]), .CLK(n562), .Q(
        reg_sscratch[27]) );
  DFFX1_LVT reg_bp_0_address_reg_27_ ( .D(wdata[27]), .CLK(n585), .Q(
        io_bp_0_address[27]) );
  DFFX1_LVT reg_mtval_reg_27_ ( .D(N1020), .CLK(n574), .Q(n_T_383[27]) );
  DFFSSRX1_LVT reg_mtvec_reg_27_ ( .D(n378), .SETB(wdata[27]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[27]) );
  DFFX1_LVT reg_stval_reg_27_ ( .D(N1409), .CLK(n561), .Q(n_T_444[27]) );
  DFFSSRX1_LVT reg_pmp_3_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[27]), .CLK(net35127), .Q(io_pmp_3_cfg_a[0]) );
  DFFX1_LVT u_T_41_reg_21_ ( .D(N1518), .CLK(n575), .Q(n_T_45[27]) );
  DFFX1_LVT u_T_49_reg_21_ ( .D(N1912), .CLK(n517), .Q(io_time[27]) );
  DFFX1_LVT reg_pmp_0_addr_reg_27_ ( .D(n_GEN_258[27]), .CLK(n537), .Q(
        io_pmp_0_addr[27]) );
  DFFX1_LVT reg_pmp_1_addr_reg_27_ ( .D(n_GEN_265[27]), .CLK(n536), .Q(
        io_pmp_1_addr[27]) );
  DFFX1_LVT reg_pmp_3_addr_reg_27_ ( .D(n_GEN_279[27]), .CLK(n535), .Q(
        io_pmp_3_addr[27]) );
  DFFX1_LVT reg_pmp_4_addr_reg_27_ ( .D(n_GEN_286[27]), .CLK(n534), .Q(
        io_pmp_4_addr[27]) );
  DFFX1_LVT reg_pmp_5_addr_reg_27_ ( .D(n_GEN_293[27]), .CLK(n533), .Q(
        io_pmp_5_addr[27]) );
  DFFX1_LVT reg_pmp_6_addr_reg_27_ ( .D(n_GEN_300[27]), .CLK(n532), .Q(
        io_pmp_6_addr[27]) );
  DFFX1_LVT reg_pmp_7_addr_reg_27_ ( .D(n_GEN_307[27]), .CLK(n538), .Q(
        io_pmp_7_addr[27]) );
  DFFX1_LVT reg_sepc_reg_27_ ( .D(net34799), .CLK(n582), .Q(reg_sepc[27]) );
  DFFX1_LVT reg_mepc_reg_27_ ( .D(net35001), .CLK(n546), .Q(reg_mepc[27]) );
  DFFX1_LVT reg_dpc_reg_27_ ( .D(net35223), .CLK(n529), .Q(reg_dpc[27]) );
  DFFX1_LVT reg_pmp_2_addr_reg_2_ ( .D(n_GEN_272[2]), .CLK(n539), .Q(
        io_pmp_2_addr[2]) );
  DFFX1_LVT u_T_41_reg_22_ ( .D(N1519), .CLK(n575), .Q(n_T_45[28]) );
  DFFX1_LVT u_T_49_reg_22_ ( .D(N1913), .CLK(n517), .Q(io_time[28]) );
  DFFX1_LVT reg_pmp_0_addr_reg_28_ ( .D(n_GEN_258[28]), .CLK(n537), .Q(
        io_pmp_0_addr[28]) );
  DFFX1_LVT reg_pmp_1_addr_reg_28_ ( .D(n_GEN_265[28]), .CLK(n536), .Q(
        io_pmp_1_addr[28]) );
  DFFX1_LVT reg_pmp_2_addr_reg_28_ ( .D(n_GEN_272[28]), .CLK(n535), .Q(
        io_pmp_2_addr[28]) );
  DFFX1_LVT reg_pmp_3_addr_reg_28_ ( .D(n_GEN_279[28]), .CLK(n534), .Q(
        io_pmp_3_addr[28]) );
  DFFX1_LVT reg_pmp_4_addr_reg_28_ ( .D(n_GEN_286[28]), .CLK(n533), .Q(
        io_pmp_4_addr[28]) );
  DFFX1_LVT reg_pmp_5_addr_reg_28_ ( .D(n_GEN_293[28]), .CLK(n532), .Q(
        io_pmp_5_addr[28]) );
  DFFX1_LVT reg_pmp_6_addr_reg_28_ ( .D(n_GEN_300[28]), .CLK(n538), .Q(
        io_pmp_6_addr[28]) );
  DFFX1_LVT reg_sepc_reg_28_ ( .D(net34796), .CLK(n583), .Q(reg_sepc[28]) );
  DFFX1_LVT reg_mepc_reg_28_ ( .D(net34998), .CLK(n547), .Q(reg_mepc[28]) );
  DFFX1_LVT reg_dpc_reg_28_ ( .D(net35220), .CLK(n530), .Q(reg_dpc[28]) );
  DFFX1_LVT reg_pmp_7_addr_reg_29_ ( .D(n_GEN_307[29]), .CLK(n540), .Q(
        io_pmp_7_addr[29]) );
  DFFX1_LVT reg_stvec_reg_29_ ( .D(wdata[29]), .CLK(n570), .Q(reg_stvec[29])
         );
  DFFX1_LVT reg_dscratch_reg_29_ ( .D(wdata[29]), .CLK(n522), .Q(
        reg_dscratch[29]) );
  DFFX1_LVT reg_mscratch_reg_29_ ( .D(wdata[29]), .CLK(n548), .Q(
        reg_mscratch[29]) );
  DFFX1_LVT reg_sscratch_reg_29_ ( .D(wdata[29]), .CLK(n562), .Q(
        reg_sscratch[29]) );
  DFFX1_LVT reg_bp_0_address_reg_29_ ( .D(wdata[29]), .CLK(n586), .Q(
        io_bp_0_address[29]) );
  DFFX1_LVT reg_mtval_reg_29_ ( .D(N1022), .CLK(n574), .Q(n_T_383[29]) );
  DFFSSRX1_LVT reg_mtvec_reg_29_ ( .D(n378), .SETB(wdata[29]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[29]) );
  DFFX1_LVT reg_stval_reg_29_ ( .D(N1411), .CLK(n561), .Q(n_T_444[29]) );
  DFFX1_LVT u_T_41_reg_23_ ( .D(N1520), .CLK(n575), .Q(n_T_45[29]) );
  DFFX1_LVT u_T_49_reg_23_ ( .D(N1914), .CLK(n517), .Q(io_time[29]) );
  DFFX1_LVT reg_pmp_0_addr_reg_29_ ( .D(n_GEN_258[29]), .CLK(n539), .Q(
        io_pmp_0_addr[29]) );
  DFFX1_LVT reg_pmp_1_addr_reg_29_ ( .D(n_GEN_265[29]), .CLK(n537), .Q(
        io_pmp_1_addr[29]) );
  DFFX1_LVT reg_pmp_2_addr_reg_29_ ( .D(n_GEN_272[29]), .CLK(n536), .Q(
        io_pmp_2_addr[29]) );
  DFFX1_LVT reg_pmp_3_addr_reg_29_ ( .D(n_GEN_279[29]), .CLK(n535), .Q(
        io_pmp_3_addr[29]) );
  DFFX1_LVT reg_pmp_4_addr_reg_29_ ( .D(n_GEN_286[29]), .CLK(n540), .Q(
        io_pmp_4_addr[29]) );
  DFFX1_LVT reg_pmp_5_addr_reg_29_ ( .D(n_GEN_293[29]), .CLK(n540), .Q(
        io_pmp_5_addr[29]) );
  DFFX1_LVT reg_pmp_6_addr_reg_29_ ( .D(n_GEN_300[29]), .CLK(n540), .Q(
        io_pmp_6_addr[29]) );
  DFFX1_LVT reg_sepc_reg_29_ ( .D(net34793), .CLK(n583), .Q(reg_sepc[29]) );
  DFFX1_LVT reg_mepc_reg_29_ ( .D(net34995), .CLK(n547), .Q(reg_mepc[29]) );
  DFFX1_LVT reg_dpc_reg_29_ ( .D(net35217), .CLK(n530), .Q(reg_dpc[29]) );
  DFFX1_LVT reg_pmp_7_addr_reg_2_ ( .D(n_GEN_307[2]), .CLK(n540), .Q(
        io_pmp_7_addr[2]) );
  DFFX1_LVT u_T_41_reg_57_ ( .D(N1554), .CLK(n575), .Q(n_T_45[63]) );
  DFFX1_LVT u_T_49_reg_57_ ( .D(N1948), .CLK(n517), .Q(n1936) );
  DFFX1_LVT reg_mcause_reg_63_ ( .D(N944), .CLK(n580), .Q(reg_mcause[63]) );
  DFFX1_LVT reg_stvec_reg_14_ ( .D(n51), .CLK(n570), .QN(reg_stvec[14]) );
  DFFX1_LVT reg_dscratch_reg_14_ ( .D(n51), .CLK(n522), .QN(reg_dscratch[14])
         );
  DFFX1_LVT reg_mscratch_reg_14_ ( .D(n51), .CLK(n548), .QN(reg_mscratch[14])
         );
  DFFX1_LVT reg_sscratch_reg_14_ ( .D(n51), .CLK(n562), .QN(reg_sscratch[14])
         );
  DFFX1_LVT reg_satp_ppn_reg_14_ ( .D(n51), .CLK(net34915), .QN(
        io_ptbr_ppn[14]) );
  DFFX1_LVT reg_mtval_reg_14_ ( .D(N1007), .CLK(n574), .Q(n_T_383[14]) );
  DFFSSRX1_LVT reg_mtvec_reg_14_ ( .D(n378), .SETB(wdata[14]), .RSTB(1'b1), 
        .CLK(n555), .QN(reg_mtvec[14]) );
  DFFX1_LVT reg_stval_reg_14_ ( .D(N1396), .CLK(n561), .Q(n_T_444[14]) );
  DFFX1_LVT u_T_41_reg_8_ ( .D(N1505), .CLK(n575), .Q(n_T_45[14]) );
  DFFX1_LVT u_T_49_reg_8_ ( .D(N1899), .CLK(n517), .Q(io_time[14]) );
  DFFX1_LVT reg_pmp_0_addr_reg_14_ ( .D(n_GEN_258[14]), .CLK(n540), .Q(
        io_pmp_0_addr[14]) );
  DFFX1_LVT reg_pmp_1_addr_reg_14_ ( .D(n_GEN_265[14]), .CLK(n540), .Q(
        io_pmp_1_addr[14]) );
  DFFX1_LVT reg_pmp_2_addr_reg_14_ ( .D(n_GEN_272[14]), .CLK(n540), .Q(
        io_pmp_2_addr[14]) );
  DFFX1_LVT reg_pmp_3_addr_reg_14_ ( .D(n_GEN_279[14]), .CLK(n540), .Q(
        io_pmp_3_addr[14]) );
  DFFX1_LVT reg_pmp_4_addr_reg_14_ ( .D(n_GEN_286[14]), .CLK(n540), .Q(
        io_pmp_4_addr[14]) );
  DFFX1_LVT reg_pmp_5_addr_reg_14_ ( .D(n_GEN_293[14]), .CLK(n540), .Q(
        io_pmp_5_addr[14]) );
  DFFX1_LVT reg_pmp_6_addr_reg_14_ ( .D(n_GEN_300[14]), .CLK(n540), .Q(
        io_pmp_6_addr[14]) );
  DFFX1_LVT reg_pmp_7_addr_reg_14_ ( .D(n_GEN_307[14]), .CLK(n540), .Q(
        io_pmp_7_addr[14]) );
  DFFX1_LVT reg_sepc_reg_14_ ( .D(net34838), .CLK(n583), .Q(reg_sepc[14]) );
  DFFX1_LVT reg_mepc_reg_14_ ( .D(net35040), .CLK(n547), .Q(reg_mepc[14]) );
  DFFX1_LVT reg_dpc_reg_14_ ( .D(net35262), .CLK(n530), .Q(reg_dpc[14]) );
  DFFX1_LVT reg_pmp_0_addr_reg_13_ ( .D(n_GEN_258[13]), .CLK(n539), .Q(
        io_pmp_0_addr[13]) );
  DFFX1_LVT reg_pmp_1_addr_reg_13_ ( .D(n_GEN_265[13]), .CLK(n539), .Q(
        io_pmp_1_addr[13]) );
  DFFX1_LVT reg_pmp_2_addr_reg_13_ ( .D(n_GEN_272[13]), .CLK(n539), .Q(
        io_pmp_2_addr[13]) );
  DFFX1_LVT reg_pmp_3_addr_reg_13_ ( .D(n_GEN_279[13]), .CLK(n539), .Q(
        io_pmp_3_addr[13]) );
  DFFX1_LVT reg_pmp_4_addr_reg_13_ ( .D(n_GEN_286[13]), .CLK(n539), .Q(
        io_pmp_4_addr[13]) );
  DFFX1_LVT reg_pmp_5_addr_reg_13_ ( .D(n_GEN_293[13]), .CLK(n539), .Q(
        io_pmp_5_addr[13]) );
  DFFX1_LVT reg_pmp_6_addr_reg_13_ ( .D(n_GEN_300[13]), .CLK(n539), .Q(
        io_pmp_6_addr[13]) );
  DFFX1_LVT reg_pmp_7_addr_reg_13_ ( .D(n_GEN_307[13]), .CLK(n539), .Q(
        io_pmp_7_addr[13]) );
  DFFX1_LVT reg_sepc_reg_13_ ( .D(net34841), .CLK(n583), .Q(reg_sepc[13]) );
  DFFX1_LVT reg_mepc_reg_13_ ( .D(net35043), .CLK(n547), .Q(reg_mepc[13]) );
  DFFX1_LVT reg_dpc_reg_13_ ( .D(net35265), .CLK(n530), .Q(reg_dpc[13]) );
  DFFX1_LVT reg_bp_0_address_reg_10_ ( .D(wdata[10]), .CLK(n586), .Q(
        io_bp_0_address[10]) );
  DFFX1_LVT reg_stvec_reg_10_ ( .D(wdata[10]), .CLK(n570), .Q(reg_stvec[10])
         );
  DFFX1_LVT reg_dscratch_reg_10_ ( .D(wdata[10]), .CLK(n522), .Q(
        reg_dscratch[10]) );
  DFFX1_LVT reg_pmp_1_cfg_x_reg ( .D(wdata[10]), .CLK(net35087), .Q(
        io_pmp_1_cfg_x) );
  DFFX1_LVT reg_mscratch_reg_10_ ( .D(wdata[10]), .CLK(n548), .Q(
        reg_mscratch[10]) );
  DFFX1_LVT reg_sscratch_reg_10_ ( .D(wdata[10]), .CLK(n562), .Q(
        reg_sscratch[10]) );
  DFFX1_LVT reg_satp_ppn_reg_10_ ( .D(wdata[10]), .CLK(net34915), .Q(
        io_ptbr_ppn[10]) );
  DFFX1_LVT reg_mtval_reg_10_ ( .D(N1003), .CLK(n574), .Q(n_T_383[10]) );
  DFFSSRX1_LVT reg_mtvec_reg_10_ ( .D(n378), .SETB(wdata[10]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[10]) );
  DFFX1_LVT reg_stval_reg_10_ ( .D(N1392), .CLK(n561), .Q(n_T_444[10]) );
  DFFX1_LVT u_T_41_reg_4_ ( .D(N1501), .CLK(n575), .Q(n_T_45[10]) );
  DFFX1_LVT u_T_49_reg_4_ ( .D(N1895), .CLK(n517), .Q(io_time[10]) );
  DFFX1_LVT reg_pmp_0_addr_reg_10_ ( .D(n_GEN_258[10]), .CLK(n539), .Q(
        io_pmp_0_addr[10]) );
  DFFX1_LVT reg_pmp_1_addr_reg_10_ ( .D(n_GEN_265[10]), .CLK(n539), .Q(
        io_pmp_1_addr[10]) );
  DFFX1_LVT reg_pmp_2_addr_reg_10_ ( .D(n_GEN_272[10]), .CLK(n539), .Q(
        io_pmp_2_addr[10]) );
  DFFX1_LVT reg_pmp_3_addr_reg_10_ ( .D(n_GEN_279[10]), .CLK(n539), .Q(
        io_pmp_3_addr[10]) );
  DFFX1_LVT reg_pmp_4_addr_reg_10_ ( .D(n_GEN_286[10]), .CLK(n538), .Q(
        io_pmp_4_addr[10]) );
  DFFX1_LVT reg_pmp_5_addr_reg_10_ ( .D(n_GEN_293[10]), .CLK(n538), .Q(
        io_pmp_5_addr[10]) );
  DFFX1_LVT reg_pmp_6_addr_reg_10_ ( .D(n_GEN_300[10]), .CLK(n538), .Q(
        io_pmp_6_addr[10]) );
  DFFX1_LVT reg_pmp_7_addr_reg_10_ ( .D(n_GEN_307[10]), .CLK(n538), .Q(
        io_pmp_7_addr[10]) );
  DFFX1_LVT reg_sepc_reg_10_ ( .D(net34850), .CLK(n583), .Q(reg_sepc[10]) );
  DFFX1_LVT reg_mepc_reg_10_ ( .D(net35052), .CLK(n547), .Q(reg_mepc[10]) );
  DFFX1_LVT reg_dpc_reg_10_ ( .D(net35274), .CLK(n530), .Q(reg_dpc[10]) );
  DFFX1_LVT reg_bp_0_address_reg_8_ ( .D(wdata[8]), .CLK(n586), .Q(
        io_bp_0_address[8]) );
  DFFX1_LVT reg_bp_0_address_reg_7_ ( .D(wdata[7]), .CLK(n586), .Q(
        io_bp_0_address[7]) );
  DFFX1_LVT reg_bp_0_address_reg_0_ ( .D(wdata[0]), .CLK(n586), .Q(
        io_bp_0_address[0]) );
  DFFX1_LVT reg_mstatus_mpp_reg_0_ ( .D(N333), .CLK(net35147), .Q(n[1930]) );
  DFFX1_LVT reg_stvec_reg_11_ ( .D(wdata[11]), .CLK(n570), .Q(reg_stvec[11])
         );
  DFFX1_LVT reg_dscratch_reg_11_ ( .D(wdata[11]), .CLK(n522), .Q(
        reg_dscratch[11]) );
  DFFX1_LVT reg_mscratch_reg_11_ ( .D(wdata[11]), .CLK(n548), .Q(
        reg_mscratch[11]) );
  DFFX1_LVT reg_sscratch_reg_11_ ( .D(wdata[11]), .CLK(n562), .Q(
        reg_sscratch[11]) );
  DFFX1_LVT reg_bp_0_address_reg_11_ ( .D(wdata[11]), .CLK(n586), .Q(
        io_bp_0_address[11]) );
  DFFX1_LVT reg_satp_ppn_reg_11_ ( .D(wdata[11]), .CLK(net34915), .Q(
        io_ptbr_ppn[11]) );
  DFFX1_LVT reg_mtval_reg_11_ ( .D(N1004), .CLK(n574), .Q(n_T_383[11]) );
  DFFSSRX1_LVT reg_mtvec_reg_11_ ( .D(n378), .SETB(wdata[11]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[11]) );
  DFFX1_LVT reg_stval_reg_11_ ( .D(N1393), .CLK(n561), .Q(n_T_444[11]) );
  DFFSSRX1_LVT reg_pmp_1_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[11]), .CLK(net35132), .Q(io_pmp_1_cfg_a[0]) );
  DFFX1_LVT u_T_41_reg_5_ ( .D(N1502), .CLK(n575), .Q(n_T_45[11]) );
  DFFX1_LVT u_T_49_reg_5_ ( .D(N1896), .CLK(n517), .Q(io_time[11]) );
  DFFX1_LVT reg_mie_reg_11_ ( .D(N617), .CLK(net34728), .Q(reg_mie[11]) );
  DFFX1_LVT reg_pmp_0_addr_reg_11_ ( .D(n_GEN_258[11]), .CLK(n538), .Q(
        io_pmp_0_addr[11]), .QN(n406) );
  DFFX1_LVT reg_pmp_1_addr_reg_11_ ( .D(n_GEN_265[11]), .CLK(n538), .Q(
        io_pmp_1_addr[11]), .QN(n402) );
  DFFX1_LVT reg_pmp_2_addr_reg_11_ ( .D(n_GEN_272[11]), .CLK(n538), .Q(
        io_pmp_2_addr[11]), .QN(n405) );
  DFFX1_LVT reg_pmp_3_addr_reg_11_ ( .D(n_GEN_279[11]), .CLK(n538), .Q(
        io_pmp_3_addr[11]), .QN(n401) );
  DFFX1_LVT reg_pmp_4_addr_reg_11_ ( .D(n_GEN_286[11]), .CLK(n538), .Q(
        io_pmp_4_addr[11]), .QN(n400) );
  DFFX1_LVT reg_pmp_5_addr_reg_11_ ( .D(n_GEN_293[11]), .CLK(n538), .Q(
        io_pmp_5_addr[11]), .QN(n399) );
  DFFX1_LVT reg_pmp_6_addr_reg_11_ ( .D(n_GEN_300[11]), .CLK(n538), .Q(
        io_pmp_6_addr[11]), .QN(n404) );
  DFFX1_LVT reg_pmp_7_addr_reg_11_ ( .D(n_GEN_307[11]), .CLK(n538), .Q(
        io_pmp_7_addr[11]), .QN(n403) );
  DFFX1_LVT reg_sepc_reg_11_ ( .D(net34847), .CLK(n583), .Q(reg_sepc[11]) );
  DFFX1_LVT reg_mepc_reg_11_ ( .D(net35049), .CLK(n547), .Q(reg_mepc[11]) );
  DFFX1_LVT reg_dpc_reg_11_ ( .D(net35271), .CLK(n530), .Q(reg_dpc[11]) );
  DFFX1_LVT u_T_1196_reg_0_ ( .D(N1691), .CLK(n594), .Q(io_status_dprv[0]) );
  DFFX1_LVT reg_pmp_0_addr_reg_8_ ( .D(n_GEN_258[8]), .CLK(n537), .Q(
        io_pmp_0_addr[8]) );
  DFFX1_LVT reg_pmp_1_addr_reg_8_ ( .D(n_GEN_265[8]), .CLK(n537), .Q(
        io_pmp_1_addr[8]) );
  DFFX1_LVT reg_pmp_2_addr_reg_8_ ( .D(n_GEN_272[8]), .CLK(n537), .Q(
        io_pmp_2_addr[8]) );
  DFFX1_LVT reg_pmp_3_addr_reg_8_ ( .D(n_GEN_279[8]), .CLK(n537), .Q(
        io_pmp_3_addr[8]) );
  DFFX1_LVT reg_pmp_4_addr_reg_8_ ( .D(n_GEN_286[8]), .CLK(n537), .Q(
        io_pmp_4_addr[8]) );
  DFFX1_LVT reg_pmp_5_addr_reg_8_ ( .D(n_GEN_293[8]), .CLK(n537), .Q(
        io_pmp_5_addr[8]) );
  DFFX1_LVT reg_pmp_6_addr_reg_8_ ( .D(n_GEN_300[8]), .CLK(n537), .Q(
        io_pmp_6_addr[8]) );
  DFFX1_LVT reg_pmp_7_addr_reg_8_ ( .D(n_GEN_307[8]), .CLK(n537), .Q(
        io_pmp_7_addr[8]) );
  DFFX1_LVT reg_sepc_reg_8_ ( .D(net34856), .CLK(n583), .Q(reg_sepc[8]) );
  DFFX1_LVT reg_mepc_reg_8_ ( .D(net35058), .CLK(n547), .Q(reg_mepc[8]) );
  DFFX1_LVT reg_dpc_reg_8_ ( .D(net35280), .CLK(n530), .Q(reg_dpc[8]) );
  DFFX1_LVT reg_stvec_reg_4_ ( .D(wdata[4]), .CLK(n570), .Q(reg_stvec[4]) );
  DFFX1_LVT reg_medeleg_reg_4_ ( .D(wdata[4]), .CLK(net35172), .Q(
        read_medeleg[4]) );
  DFFX1_LVT reg_dscratch_reg_4_ ( .D(wdata[4]), .CLK(n522), .Q(reg_dscratch[4]) );
  DFFX1_LVT reg_mscratch_reg_4_ ( .D(wdata[4]), .CLK(n548), .Q(reg_mscratch[4]) );
  DFFX1_LVT reg_sscratch_reg_4_ ( .D(wdata[4]), .CLK(n562), .Q(reg_sscratch[4]) );
  DFFX1_LVT reg_bp_0_address_reg_4_ ( .D(wdata[4]), .CLK(n586), .Q(
        io_bp_0_address[4]) );
  DFFX1_LVT reg_bp_0_control_s_reg ( .D(wdata[4]), .CLK(net35319), .Q(
        io_bp_0_control_s) );
  DFFX1_LVT reg_satp_ppn_reg_4_ ( .D(wdata[4]), .CLK(net34915), .Q(
        io_ptbr_ppn[4]) );
  DFFSSRX1_LVT reg_mtvec_reg_4_ ( .D(n378), .SETB(wdata[4]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[4]) );
  DFFX1_LVT reg_scause_reg_4_ ( .D(N1274), .CLK(n558), .Q(reg_scause[4]) );
  DFFX1_LVT reg_stval_reg_4_ ( .D(N1386), .CLK(n561), .Q(n_T_444[4]) );
  DFFSSRX1_LVT reg_pmp_0_cfg_a_reg_1_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[4]), 
        .CLK(net34905), .Q(io_pmp_0_cfg_a[1]) );
  DFFX1_LVT u_T_39_reg_4_ ( .D(N1432), .CLK(n594), .Q(n_T_45[4]) );
  DFFX1_LVT u_T_47_reg_4_ ( .D(N1826), .CLK(n591), .Q(io_time[4]), .QN(n454)
         );
  DFFX1_LVT reg_mtval_reg_4_ ( .D(N997), .CLK(n574), .Q(n_T_383[4]) );
  DFFX1_LVT reg_pmp_0_addr_reg_4_ ( .D(n_GEN_258[4]), .CLK(n537), .Q(
        io_pmp_0_addr[4]) );
  DFFX1_LVT reg_pmp_1_addr_reg_4_ ( .D(n_GEN_265[4]), .CLK(n537), .Q(
        io_pmp_1_addr[4]) );
  DFFX1_LVT reg_pmp_2_addr_reg_4_ ( .D(n_GEN_272[4]), .CLK(n537), .Q(
        io_pmp_2_addr[4]) );
  DFFX1_LVT reg_pmp_3_addr_reg_4_ ( .D(n_GEN_279[4]), .CLK(n537), .Q(
        io_pmp_3_addr[4]) );
  DFFX1_LVT reg_pmp_4_addr_reg_4_ ( .D(n_GEN_286[4]), .CLK(n536), .Q(
        io_pmp_4_addr[4]) );
  DFFX1_LVT reg_pmp_5_addr_reg_4_ ( .D(n_GEN_293[4]), .CLK(n536), .Q(
        io_pmp_5_addr[4]) );
  DFFX1_LVT reg_pmp_6_addr_reg_4_ ( .D(n_GEN_300[4]), .CLK(n536), .Q(
        io_pmp_6_addr[4]) );
  DFFX1_LVT reg_pmp_7_addr_reg_4_ ( .D(n_GEN_307[4]), .CLK(n536), .Q(
        io_pmp_7_addr[4]) );
  DFFX1_LVT reg_fflags_reg_4_ ( .D(n_GEN_345[4]), .CLK(n594), .Q(read_fcsr[4])
         );
  DFFX1_LVT reg_sepc_reg_4_ ( .D(net34868), .CLK(n583), .Q(reg_sepc[4]) );
  DFFX1_LVT reg_mepc_reg_4_ ( .D(net35070), .CLK(n547), .Q(reg_mepc[4]) );
  DFFX1_LVT reg_dpc_reg_4_ ( .D(net35292), .CLK(n530), .Q(reg_dpc[4]) );
  DFFSSRX1_LVT reg_misa_reg_2_ ( .D(n387), .SETB(wdata[2]), .RSTB(n590), .CLK(
        net35137), .QN(io_status_isa_2_) );
  DFFX1_LVT reg_scounteren_reg_1_ ( .D(wdata[1]), .CLK(net34940), .Q(
        read_scounteren[1]) );
  DFFX1_LVT reg_mcounteren_reg_1_ ( .D(wdata[1]), .CLK(net34945), .Q(
        read_mcounteren[1]) );
  DFFX1_LVT reg_mideleg_reg_1_ ( .D(wdata[1]), .CLK(net35167), .Q(
        read_mideleg_1), .QN(n407) );
  DFFX1_LVT reg_dscratch_reg_1_ ( .D(wdata[1]), .CLK(n522), .Q(reg_dscratch[1]) );
  DFFX1_LVT reg_mscratch_reg_1_ ( .D(wdata[1]), .CLK(n548), .Q(reg_mscratch[1]) );
  DFFX1_LVT reg_sscratch_reg_1_ ( .D(wdata[1]), .CLK(n562), .Q(reg_sscratch[1]) );
  DFFX1_LVT reg_bp_0_address_reg_1_ ( .D(wdata[1]), .CLK(n586), .Q(
        io_bp_0_address[1]) );
  DFFX1_LVT reg_satp_ppn_reg_1_ ( .D(wdata[1]), .CLK(net34915), .Q(
        io_ptbr_ppn[1]) );
  DFFX1_LVT reg_scause_reg_1_ ( .D(N1271), .CLK(n558), .Q(reg_scause[1]) );
  DFFX1_LVT reg_stval_reg_1_ ( .D(N1383), .CLK(n561), .Q(n_T_444[1]) );
  DFFSSRX1_LVT reg_bp_0_control_w_reg ( .D(n375), .SETB(1'b1), .RSTB(wdata[1]), 
        .CLK(net35314), .Q(io_bp_0_control_w) );
  DFFX1_LVT u_T_39_reg_1_ ( .D(N1429), .CLK(n593), .Q(n_T_45[1]) );
  DFFX1_LVT u_T_47_reg_1_ ( .D(N1823), .CLK(n591), .Q(io_time[1]) );
  DFFX1_LVT reg_mcause_reg_1_ ( .D(N882), .CLK(n580), .Q(reg_mcause[1]) );
  DFFX1_LVT reg_mstatus_sie_reg ( .D(n1062), .CLK(n1915), .Q(n1935) );
  DFFX1_LVT reg_mstatus_spie_reg ( .D(n1914), .CLK(n1915), .Q(n1933) );
  DFFX1_LVT reg_stvec_reg_5_ ( .D(wdata[5]), .CLK(n570), .Q(reg_stvec[5]) );
  DFFX1_LVT reg_mideleg_reg_5_ ( .D(wdata[5]), .CLK(net35167), .Q(
        read_mideleg_5), .QN(n427) );
  DFFX1_LVT reg_dscratch_reg_5_ ( .D(wdata[5]), .CLK(n522), .Q(reg_dscratch[5]) );
  DFFX1_LVT reg_mscratch_reg_5_ ( .D(wdata[5]), .CLK(n548), .Q(reg_mscratch[5]) );
  DFFX1_LVT reg_sscratch_reg_5_ ( .D(wdata[5]), .CLK(n562), .Q(reg_sscratch[5]) );
  DFFX1_LVT reg_bp_0_address_reg_5_ ( .D(wdata[5]), .CLK(n586), .Q(
        io_bp_0_address[5]) );
  DFFX1_LVT reg_satp_ppn_reg_5_ ( .D(wdata[5]), .CLK(net34915), .Q(
        io_ptbr_ppn[5]) );
  DFFSSRX1_LVT reg_mtvec_reg_5_ ( .D(n378), .SETB(wdata[5]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[5]) );
  DFFX1_LVT reg_stval_reg_5_ ( .D(N1387), .CLK(net34930), .Q(n_T_444[5]) );
  DFFX1_LVT u_T_39_reg_5_ ( .D(N1433), .CLK(n593), .Q(n_T_45[5]) );
  DFFSSRX1_LVT reg_misa_reg_3_ ( .D(n1346), .SETB(wdata[5]), .RSTB(n590), 
        .CLK(net35137), .QN(io_status_isa_3_) );
  DFFX1_LVT reg_stvec_reg_3_ ( .D(wdata[3]), .CLK(n571), .Q(reg_stvec[3]) );
  DFFX1_LVT reg_medeleg_reg_3_ ( .D(wdata[3]), .CLK(net35172), .Q(
        read_medeleg[3]) );
  DFFX1_LVT reg_dscratch_reg_3_ ( .D(wdata[3]), .CLK(n522), .Q(reg_dscratch[3]) );
  DFFX1_LVT reg_mscratch_reg_3_ ( .D(wdata[3]), .CLK(n548), .Q(reg_mscratch[3]) );
  DFFX1_LVT reg_sscratch_reg_3_ ( .D(wdata[3]), .CLK(n562), .Q(reg_sscratch[3]) );
  DFFX1_LVT reg_bp_0_address_reg_3_ ( .D(wdata[3]), .CLK(n587), .Q(
        io_bp_0_address[3]) );
  DFFX1_LVT reg_bp_0_control_u_reg ( .D(wdata[3]), .CLK(net35319), .Q(
        io_bp_0_control_u) );
  DFFX1_LVT reg_satp_ppn_reg_3_ ( .D(wdata[3]), .CLK(net34915), .Q(
        io_ptbr_ppn[3]) );
  DFFSSRX1_LVT reg_mtvec_reg_3_ ( .D(n378), .SETB(wdata[3]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[3]) );
  DFFX1_LVT reg_scause_reg_3_ ( .D(N1273), .CLK(n558), .Q(reg_scause[3]) );
  DFFX1_LVT reg_stval_reg_3_ ( .D(N1385), .CLK(net34930), .Q(n_T_444[3]) );
  DFFX1_LVT reg_mcause_reg_3_ ( .D(N884), .CLK(n580), .Q(reg_mcause[3]) );
  DFFX1_LVT u_T_47_reg_3_ ( .D(N1825), .CLK(n591), .Q(io_time[3]) );
  DFFX1_LVT u_T_39_reg_3_ ( .D(N1431), .CLK(n593), .Q(n_T_45[3]) );
  DFFSSRX1_LVT reg_pmp_0_cfg_a_reg_0_ ( .D(n375), .SETB(1'b1), .RSTB(wdata[3]), 
        .CLK(net34905), .Q(io_pmp_0_cfg_a[0]) );
  DFFX1_LVT reg_mie_reg_3_ ( .D(N609), .CLK(net34728), .Q(reg_mie[3]) );
  DFFX1_LVT reg_mtval_reg_3_ ( .D(N996), .CLK(n574), .Q(n_T_383[3]) );
  DFFX1_LVT reg_pmp_0_addr_reg_3_ ( .D(n_GEN_258[3]), .CLK(n536), .Q(
        io_pmp_0_addr[3]), .QN(n415) );
  DFFX1_LVT reg_pmp_1_addr_reg_3_ ( .D(n_GEN_265[3]), .CLK(n536), .Q(
        io_pmp_1_addr[3]), .QN(n411) );
  DFFX1_LVT reg_pmp_2_addr_reg_3_ ( .D(n_GEN_272[3]), .CLK(n536), .Q(
        io_pmp_2_addr[3]), .QN(n410) );
  DFFX1_LVT reg_pmp_3_addr_reg_3_ ( .D(n_GEN_279[3]), .CLK(n536), .Q(
        io_pmp_3_addr[3]), .QN(n409) );
  DFFX1_LVT reg_pmp_4_addr_reg_3_ ( .D(n_GEN_286[3]), .CLK(n536), .Q(
        io_pmp_4_addr[3]), .QN(n408) );
  DFFX1_LVT reg_pmp_5_addr_reg_3_ ( .D(n_GEN_293[3]), .CLK(n536), .Q(
        io_pmp_5_addr[3]), .QN(n414) );
  DFFX1_LVT reg_pmp_6_addr_reg_3_ ( .D(n_GEN_300[3]), .CLK(n536), .Q(
        io_pmp_6_addr[3]), .QN(n413) );
  DFFX1_LVT reg_pmp_7_addr_reg_3_ ( .D(n_GEN_307[3]), .CLK(n536), .Q(
        io_pmp_7_addr[3]), .QN(n412) );
  DFFX1_LVT reg_fflags_reg_3_ ( .D(n_GEN_345[3]), .CLK(n593), .Q(read_fcsr[3])
         );
  DFFX1_LVT reg_sepc_reg_3_ ( .D(net34871), .CLK(n583), .Q(reg_sepc[3]) );
  DFFX1_LVT reg_mepc_reg_3_ ( .D(net35073), .CLK(n547), .Q(reg_mepc[3]) );
  DFFX1_LVT reg_dpc_reg_3_ ( .D(net35295), .CLK(n530), .Q(reg_dpc[3]) );
  DFFSSRX1_LVT reg_misa_reg_5_ ( .D(n387), .SETB(wdata[5]), .RSTB(n590), .CLK(
        net35137), .QN(n1923) );
  DFFX1_LVT u_T_47_reg_5_ ( .D(N1827), .CLK(n591), .Q(io_time[5]) );
  DFFX1_LVT reg_mie_reg_5_ ( .D(N611), .CLK(net34728), .Q(reg_mie[5]) );
  DFFX1_LVT reg_mtval_reg_5_ ( .D(N998), .CLK(net34895), .Q(n_T_383[5]) );
  DFFX1_LVT reg_frm_reg_0_ ( .D(n_GEN_155[0]), .CLK(net34900), .Q(
        io_fcsr_rm[0]) );
  DFFX1_LVT reg_pmp_0_addr_reg_5_ ( .D(n_GEN_258[5]), .CLK(n535), .Q(
        io_pmp_0_addr[5]) );
  DFFX1_LVT reg_pmp_1_addr_reg_5_ ( .D(n_GEN_265[5]), .CLK(n535), .Q(
        io_pmp_1_addr[5]) );
  DFFX1_LVT reg_pmp_2_addr_reg_5_ ( .D(n_GEN_272[5]), .CLK(n535), .Q(
        io_pmp_2_addr[5]) );
  DFFX1_LVT reg_pmp_3_addr_reg_5_ ( .D(n_GEN_279[5]), .CLK(n535), .Q(
        io_pmp_3_addr[5]) );
  DFFX1_LVT reg_pmp_4_addr_reg_5_ ( .D(n_GEN_286[5]), .CLK(n535), .Q(
        io_pmp_4_addr[5]) );
  DFFX1_LVT reg_pmp_5_addr_reg_5_ ( .D(n_GEN_293[5]), .CLK(n535), .Q(
        io_pmp_5_addr[5]) );
  DFFX1_LVT reg_pmp_6_addr_reg_5_ ( .D(n_GEN_300[5]), .CLK(n535), .Q(
        io_pmp_6_addr[5]) );
  DFFX1_LVT reg_pmp_7_addr_reg_5_ ( .D(n_GEN_307[5]), .CLK(n535), .Q(
        io_pmp_7_addr[5]) );
  DFFX1_LVT reg_sepc_reg_5_ ( .D(net34865), .CLK(n583), .Q(reg_sepc[5]) );
  DFFX1_LVT reg_mepc_reg_5_ ( .D(net35067), .CLK(n547), .Q(reg_mepc[5]) );
  DFFX1_LVT reg_dpc_reg_5_ ( .D(net35289), .CLK(n530), .Q(reg_dpc[5]) );
  DFFX1_LVT reg_mie_reg_1_ ( .D(N607), .CLK(net34728), .Q(reg_mie[1]) );
  DFFX1_LVT reg_mtval_reg_1_ ( .D(N994), .CLK(net34895), .Q(n_T_383[1]) );
  DFFX1_LVT reg_frm_reg_1_ ( .D(n_GEN_155[1]), .CLK(net34900), .Q(
        io_fcsr_rm[1]) );
  DFFX1_LVT reg_stvec_reg_6_ ( .D(wdata[6]), .CLK(n571), .Q(reg_stvec[6]) );
  DFFX1_LVT reg_medeleg_reg_6_ ( .D(wdata[6]), .CLK(net35172), .Q(
        read_medeleg_6) );
  DFFX1_LVT reg_dscratch_reg_6_ ( .D(wdata[6]), .CLK(n522), .Q(reg_dscratch[6]) );
  DFFX1_LVT reg_mscratch_reg_6_ ( .D(wdata[6]), .CLK(n548), .Q(reg_mscratch[6]) );
  DFFX1_LVT reg_sscratch_reg_6_ ( .D(wdata[6]), .CLK(n562), .Q(reg_sscratch[6]) );
  DFFX1_LVT reg_bp_0_address_reg_6_ ( .D(wdata[6]), .CLK(n587), .Q(
        io_bp_0_address[6]) );
  DFFX1_LVT reg_bp_0_control_m_reg ( .D(wdata[6]), .CLK(net35319), .Q(
        io_bp_0_control_m) );
  DFFX1_LVT reg_satp_ppn_reg_6_ ( .D(wdata[6]), .CLK(net34915), .Q(
        io_ptbr_ppn[6]) );
  DFFSSRX1_LVT reg_mtvec_reg_6_ ( .D(n378), .SETB(wdata[6]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[6]) );
  DFFX1_LVT reg_stval_reg_6_ ( .D(N1388), .CLK(net34930), .Q(n_T_444[6]) );
  DFFX1_LVT u_T_41_reg_0_ ( .D(N1497), .CLK(n575), .Q(n_T_45[6]), .QN(n455) );
  DFFX1_LVT u_T_49_reg_0_ ( .D(N1891), .CLK(n517), .Q(io_time[6]), .QN(n456)
         );
  DFFX1_LVT reg_mtval_reg_6_ ( .D(N999), .CLK(net34895), .Q(n_T_383[6]) );
  DFFX1_LVT reg_pmp_0_addr_reg_6_ ( .D(n_GEN_258[6]), .CLK(n535), .Q(
        io_pmp_0_addr[6]) );
  DFFX1_LVT reg_pmp_1_addr_reg_6_ ( .D(n_GEN_265[6]), .CLK(n535), .Q(
        io_pmp_1_addr[6]) );
  DFFX1_LVT reg_pmp_2_addr_reg_6_ ( .D(n_GEN_272[6]), .CLK(n535), .Q(
        io_pmp_2_addr[6]) );
  DFFX1_LVT reg_pmp_3_addr_reg_6_ ( .D(n_GEN_279[6]), .CLK(n535), .Q(
        io_pmp_3_addr[6]) );
  DFFX1_LVT reg_pmp_4_addr_reg_6_ ( .D(n_GEN_286[6]), .CLK(n534), .Q(
        io_pmp_4_addr[6]) );
  DFFX1_LVT reg_pmp_5_addr_reg_6_ ( .D(n_GEN_293[6]), .CLK(n534), .Q(
        io_pmp_5_addr[6]) );
  DFFX1_LVT reg_pmp_6_addr_reg_6_ ( .D(n_GEN_300[6]), .CLK(n534), .Q(
        io_pmp_6_addr[6]) );
  DFFX1_LVT reg_pmp_7_addr_reg_6_ ( .D(n_GEN_307[6]), .CLK(n534), .Q(
        io_pmp_7_addr[6]) );
  DFFX1_LVT reg_sepc_reg_6_ ( .D(net34862), .CLK(n583), .Q(reg_sepc[6]) );
  DFFX1_LVT reg_mepc_reg_6_ ( .D(net35064), .CLK(n547), .Q(reg_mepc[6]) );
  DFFX1_LVT reg_dpc_reg_6_ ( .D(net35286), .CLK(n530), .Q(reg_dpc[6]) );
  DFFX1_LVT reg_pmp_0_addr_reg_1_ ( .D(n_GEN_258[1]), .CLK(n534), .Q(
        io_pmp_0_addr[1]) );
  DFFX1_LVT reg_pmp_1_addr_reg_1_ ( .D(n_GEN_265[1]), .CLK(n534), .Q(
        io_pmp_1_addr[1]) );
  DFFX1_LVT reg_pmp_2_addr_reg_1_ ( .D(n_GEN_272[1]), .CLK(n534), .Q(
        io_pmp_2_addr[1]) );
  DFFX1_LVT reg_pmp_3_addr_reg_1_ ( .D(n_GEN_279[1]), .CLK(n534), .Q(
        io_pmp_3_addr[1]) );
  DFFX1_LVT reg_pmp_4_addr_reg_1_ ( .D(n_GEN_286[1]), .CLK(n534), .Q(
        io_pmp_4_addr[1]) );
  DFFX1_LVT reg_pmp_5_addr_reg_1_ ( .D(n_GEN_293[1]), .CLK(n534), .Q(
        io_pmp_5_addr[1]) );
  DFFX1_LVT reg_pmp_6_addr_reg_1_ ( .D(n_GEN_300[1]), .CLK(n534), .Q(
        io_pmp_6_addr[1]) );
  DFFX1_LVT reg_pmp_7_addr_reg_1_ ( .D(n_GEN_307[1]), .CLK(n534), .Q(
        io_pmp_7_addr[1]) );
  DFFX1_LVT reg_fflags_reg_1_ ( .D(n_GEN_345[1]), .CLK(n594), .Q(read_fcsr[1])
         );
  DFFSSRX1_LVT reg_pmp_0_cfg_w_reg ( .D(wdata[1]), .SETB(1'b1), .RSTB(wdata[0]), .CLK(net34733), .Q(io_pmp_0_cfg_w) );
  DFFX1_LVT reg_dcsr_prv_reg_1_ ( .D(n2155), .CLK(n593), .Q(n_T_389_1) );
  DFFX1_LVT reg_sepc_reg_1_ ( .D(net34877), .CLK(n583), .Q(reg_sepc[1]) );
  DFFX1_LVT reg_mepc_reg_1_ ( .D(net35079), .CLK(n547), .Q(reg_mepc[1]) );
  DFFX1_LVT reg_dpc_reg_1_ ( .D(net35301), .CLK(n530), .Q(reg_dpc[1]) );
  DFFX1_LVT reg_mip_ssip_reg ( .D(n2162), .CLK(n533), .Q(n_T_61_1) );
  DFFSSRX1_LVT reg_misa_reg_0_ ( .D(n387), .SETB(wdata[0]), .RSTB(n590), .CLK(
        net35137), .Q(io_status_isa_0__BAR), .QN(io_status_isa_0_) );
  DFFX1_LVT reg_pmp_0_addr_reg_7_ ( .D(n_GEN_258[7]), .CLK(n533), .Q(
        io_pmp_0_addr[7]), .QN(n398) );
  DFFX1_LVT reg_pmp_1_addr_reg_7_ ( .D(n_GEN_265[7]), .CLK(n533), .Q(
        io_pmp_1_addr[7]), .QN(n397) );
  DFFX1_LVT reg_pmp_2_addr_reg_7_ ( .D(n_GEN_272[7]), .CLK(n533), .Q(
        io_pmp_2_addr[7]), .QN(n393) );
  DFFX1_LVT reg_pmp_3_addr_reg_7_ ( .D(n_GEN_279[7]), .CLK(n533), .Q(
        io_pmp_3_addr[7]), .QN(n396) );
  DFFX1_LVT reg_pmp_4_addr_reg_7_ ( .D(n_GEN_286[7]), .CLK(n533), .Q(
        io_pmp_4_addr[7]), .QN(n395) );
  DFFX1_LVT reg_pmp_5_addr_reg_7_ ( .D(n_GEN_293[7]), .CLK(n533), .Q(
        io_pmp_5_addr[7]), .QN(n392) );
  DFFX1_LVT reg_pmp_6_addr_reg_7_ ( .D(n_GEN_300[7]), .CLK(n533), .Q(
        io_pmp_6_addr[7]), .QN(n391) );
  DFFX1_LVT reg_pmp_7_addr_reg_7_ ( .D(n_GEN_307[7]), .CLK(n533), .Q(
        io_pmp_7_addr[7]), .QN(n394) );
  DFFX1_LVT reg_sepc_reg_7_ ( .D(net34859), .CLK(net34880), .Q(reg_sepc[7]) );
  DFFX1_LVT reg_mepc_reg_7_ ( .D(net35061), .CLK(net35082), .Q(reg_mepc[7]) );
  DFFX1_LVT reg_dpc_reg_7_ ( .D(net35283), .CLK(net35304), .Q(reg_dpc[7]) );
  DFFX1_LVT reg_dscratch_reg_9_ ( .D(wdata[9]), .CLK(n522), .Q(reg_dscratch[9]) );
  DFFX1_LVT reg_mscratch_reg_9_ ( .D(wdata[9]), .CLK(n548), .Q(reg_mscratch[9]) );
  DFFX1_LVT reg_sscratch_reg_9_ ( .D(wdata[9]), .CLK(n562), .Q(reg_sscratch[9]) );
  DFFX1_LVT reg_bp_0_address_reg_9_ ( .D(wdata[9]), .CLK(n587), .Q(
        io_bp_0_address[9]) );
  DFFX1_LVT reg_satp_ppn_reg_9_ ( .D(wdata[9]), .CLK(net34915), .Q(
        io_ptbr_ppn[9]) );
  DFFX1_LVT reg_mtval_reg_9_ ( .D(N1002), .CLK(net34895), .Q(n_T_383[9]) );
  DFFSSRX1_LVT reg_mtvec_reg_9_ ( .D(n376), .SETB(wdata[9]), .RSTB(1'b1), 
        .CLK(n556), .QN(reg_mtvec[9]) );
  DFFX1_LVT reg_stval_reg_9_ ( .D(N1391), .CLK(net34930), .Q(n_T_444[9]) );
  DFFX1_LVT u_T_41_reg_3_ ( .D(N1500), .CLK(n575), .Q(n_T_45[9]) );
  DFFX1_LVT u_T_49_reg_3_ ( .D(N1894), .CLK(n517), .Q(io_time[9]) );
  DFFX1_LVT reg_mie_reg_9_ ( .D(N615), .CLK(net34728), .Q(reg_mie[9]) );
  DFFX1_LVT reg_wfi_reg ( .D(N1821), .CLK(n591), .Q(io_status_wfi), .QN(n472)
         );
  DFFX1_LVT reg_pmp_1_addr_reg_9_ ( .D(n_GEN_265[9]), .CLK(n533), .Q(
        io_pmp_1_addr[9]), .QN(n425) );
  DFFX1_LVT reg_pmp_2_addr_reg_9_ ( .D(n_GEN_272[9]), .CLK(n533), .Q(
        io_pmp_2_addr[9]), .QN(n421) );
  DFFX1_LVT reg_pmp_3_addr_reg_9_ ( .D(n_GEN_279[9]), .CLK(n533), .Q(
        io_pmp_3_addr[9]), .QN(n418) );
  DFFX1_LVT reg_pmp_4_addr_reg_9_ ( .D(n_GEN_286[9]), .CLK(n532), .Q(
        io_pmp_4_addr[9]), .QN(n423) );
  DFFX1_LVT reg_pmp_5_addr_reg_9_ ( .D(n_GEN_293[9]), .CLK(n532), .Q(
        io_pmp_5_addr[9]), .QN(n422) );
  DFFX1_LVT reg_pmp_6_addr_reg_9_ ( .D(n_GEN_300[9]), .CLK(n532), .Q(
        io_pmp_6_addr[9]), .QN(n420) );
  DFFX1_LVT reg_pmp_7_addr_reg_9_ ( .D(n_GEN_307[9]), .CLK(n532), .Q(
        io_pmp_7_addr[9]), .QN(n424) );
  DFFSSRX1_LVT reg_pmp_1_cfg_w_reg ( .D(wdata[8]), .SETB(1'b1), .RSTB(wdata[9]), .CLK(net35087), .Q(io_pmp_1_cfg_w) );
  DFFX1_LVT reg_sepc_reg_9_ ( .D(net34853), .CLK(net34880), .Q(reg_sepc[9]) );
  DFFX1_LVT reg_mepc_reg_9_ ( .D(net35055), .CLK(net35082), .Q(reg_mepc[9]) );
  DFFX1_LVT reg_dpc_reg_9_ ( .D(net35277), .CLK(net35304), .Q(reg_dpc[9]) );
  DFFX1_LVT reg_pmp_0_addr_reg_12_ ( .D(n_GEN_258[12]), .CLK(n532), .Q(
        io_pmp_0_addr[12]) );
  DFFX1_LVT reg_pmp_1_addr_reg_12_ ( .D(n_GEN_265[12]), .CLK(n532), .Q(
        io_pmp_1_addr[12]) );
  DFFX1_LVT reg_pmp_2_addr_reg_12_ ( .D(n_GEN_272[12]), .CLK(n532), .Q(
        io_pmp_2_addr[12]) );
  DFFX1_LVT reg_pmp_3_addr_reg_12_ ( .D(n_GEN_279[12]), .CLK(n532), .Q(
        io_pmp_3_addr[12]) );
  DFFX1_LVT reg_pmp_4_addr_reg_12_ ( .D(n_GEN_286[12]), .CLK(n532), .Q(
        io_pmp_4_addr[12]) );
  DFFX1_LVT reg_pmp_5_addr_reg_12_ ( .D(n_GEN_293[12]), .CLK(n532), .Q(
        io_pmp_5_addr[12]) );
  DFFX1_LVT reg_pmp_6_addr_reg_12_ ( .D(n_GEN_300[12]), .CLK(n532), .Q(
        io_pmp_6_addr[12]) );
  DFFX1_LVT reg_pmp_7_addr_reg_12_ ( .D(n_GEN_307[12]), .CLK(n532), .Q(
        io_pmp_7_addr[12]) );
  DFFX1_LVT reg_sepc_reg_12_ ( .D(net34844), .CLK(net34880), .Q(reg_sepc[12])
         );
  DFFX1_LVT reg_mepc_reg_12_ ( .D(net35046), .CLK(net35082), .Q(reg_mepc[12])
         );
  DFFX1_LVT reg_dpc_reg_12_ ( .D(net35268), .CLK(net35304), .Q(reg_dpc[12]) );
  DFFX1_LVT u_T_1196_reg_1_ ( .D(N1692), .CLK(n593), .Q(io_status_dprv[1]) );
  SNPS_CLOCK_GATE_HIGH_CSRFile_0_5 clk_gate_reg_mstatus_spie_reg ( .CLK(n593), 
        .EN(n1917), .ENCLK(n1915), .TE(1'b0) );
  DFFX1_LVT reg_custom_0_reg_9_ ( .D(n1911), .CLK(n594), .Q(n1912), .QN(
        io_customCSRs_0_value[9]) );
  DFFX1_LVT reg_custom_0_reg_3_ ( .D(n1909), .CLK(n594), .Q(n1910), .QN(
        io_customCSRs_0_value[3]) );
  DFFX1_LVT reg_mstatus_prv_reg_0_ ( .D(n2157), .CLK(n594), .Q(
        io_status_prv[0]), .QN(n429) );
  DFFX1_LVT reg_mstatus_prv_reg_1_ ( .D(n2160), .CLK(n594), .Q(
        io_status_prv[1]), .QN(n381) );
  DFFX1_LVT reg_pmp_6_cfg_l_reg ( .D(n374), .CLK(net35102), .Q(io_pmp_6_cfg_l), 
        .QN(n439) );
  INVX0_LVT reg_dcsr_cause_reg_2__U4 ( .A(n1499), .Y(n372) );
  DFFX1_LVT reg_dcsr_cause_reg_2_ ( .D(n373), .CLK(net35177), .QN(n_T_389[8])
         );
  DFFX1_LVT u_T_41_reg_48_ ( .D(N1545), .CLK(net34890), .Q(n_T_45[54]) );
  DFFX1_LVT reg_mtvec_reg_0_ ( .D(n371), .CLK(net34950), .Q(n416), .QN(n659)
         );
  DFFX1_LVT reg_mtvec_reg_31_ ( .D(n370), .CLK(net34950), .QN(reg_mtvec[31])
         );
  DFFX1_LVT reg_pmp_6_cfg_w_reg ( .D(n369), .CLK(net35107), .Q(io_pmp_6_cfg_w)
         );
  INVX0_LVT reg_misa_reg_12__U4 ( .A(wdata[12]), .Y(n367) );
  OA21X1_LVT reg_misa_reg_12__U2 ( .A1(n367), .A2(n387), .A3(n590), .Y(n368)
         );
  DFFX1_LVT reg_misa_reg_12_ ( .D(n368), .CLK(net35137), .Q(
        io_status_isa_12__BAR), .QN(io_status_isa_12_) );
  DFFX1_LVT reg_pmp_0_cfg_x_reg ( .D(n1483), .CLK(net34733), .QN(
        io_pmp_0_cfg_x) );
  DFFX1_LVT reg_bp_0_address_reg_14_ ( .D(n51), .CLK(n586), .QN(
        io_bp_0_address[14]) );
  DFFX1_LVT reg_bp_0_address_reg_12_ ( .D(n367), .CLK(n586), .QN(
        io_bp_0_address[12]) );
  DFFX1_LVT reg_bp_0_address_reg_2_ ( .D(n1483), .CLK(n586), .QN(
        io_bp_0_address[2]) );
  DFFX1_LVT reg_scounteren_reg_2_ ( .D(n1483), .CLK(net34940), .QN(
        read_scounteren[2]) );
  DFFX1_LVT reg_mcounteren_reg_2_ ( .D(n1483), .CLK(net34945), .QN(
        read_mcounteren[2]) );
  DFFX1_LVT reg_medeleg_reg_12_ ( .D(n367), .CLK(net35172), .QN(
        read_medeleg_12) );
  DFFX1_LVT reg_medeleg_reg_2_ ( .D(n1483), .CLK(net35172), .QN(
        read_medeleg[2]) );
  DFFX1_LVT reg_sscratch_reg_12_ ( .D(n367), .CLK(n567), .QN(reg_sscratch[12])
         );
  DFFX1_LVT reg_sscratch_reg_2_ ( .D(n1483), .CLK(n567), .QN(reg_sscratch[2])
         );
  DFFX1_LVT reg_mscratch_reg_12_ ( .D(n367), .CLK(n553), .QN(reg_mscratch[12])
         );
  DFFX1_LVT reg_mscratch_reg_2_ ( .D(n1483), .CLK(n553), .QN(reg_mscratch[2])
         );
  DFFX1_LVT reg_dscratch_reg_12_ ( .D(n367), .CLK(n527), .QN(reg_dscratch[12])
         );
  DFFX1_LVT reg_dscratch_reg_2_ ( .D(n1483), .CLK(n527), .QN(reg_dscratch[2])
         );
  DFFX1_LVT reg_dcsr_cause_reg_0_ ( .D(n366), .CLK(net35177), .Q(n_T_389[6])
         );
  OA21X1_LVT reg_mstatus_mie_reg_U2 ( .A1(n1346), .A2(n1041), .A3(n194), .Y(
        n365) );
  DFFX1_LVT reg_mstatus_mie_reg ( .D(n365), .CLK(net35147), .Q(n383), .QN(
        n1934) );
  AO222X1_LVT U3 ( .A1(n323), .A2(n1185), .A3(io_interrupts_debug), .A4(1'b1), 
        .A5(n1183), .A6(n1184), .Y(io_interrupt_cause[2]) );
  AO221X1_LVT U4 ( .A1(1'b1), .A2(n333), .A3(n1153), .A4(n_T_383[21]), .A5(
        n334), .Y(n336) );
  AO221X1_LVT U5 ( .A1(1'b1), .A2(n1533), .A3(n_T_45[8]), .A4(n1689), .A5(n286), .Y(n288) );
  AO221X1_LVT U6 ( .A1(1'b1), .A2(n277), .A3(n1162), .A4(n1961), .A5(n278), 
        .Y(n280) );
  AO221X1_LVT U7 ( .A1(1'b1), .A2(n1650), .A3(n1485), .A4(reg_mscratch[38]), 
        .A5(n282), .Y(n283) );
  AO221X1_LVT U8 ( .A1(1'b1), .A2(n264), .A3(n1689), .A4(n_T_45[31]), .A5(n265), .Y(n267) );
  AO221X1_LVT U9 ( .A1(1'b1), .A2(n267), .A3(n1507), .A4(io_pmp_3_cfg_l), .A5(
        n268), .Y(n269) );
  AO221X1_LVT U10 ( .A1(1'b1), .A2(n263), .A3(n1510), .A4(reg_dscratch[31]), 
        .A5(n269), .Y(n270) );
  AO221X1_LVT U11 ( .A1(1'b1), .A2(n262), .A3(n1485), .A4(reg_mscratch[31]), 
        .A5(n270), .Y(io_rw_rdata[31]) );
  AO221X1_LVT U12 ( .A1(1'b1), .A2(n255), .A3(n1507), .A4(io_pmp_3_cfg_a[1]), 
        .A5(n256), .Y(n258) );
  AO221X1_LVT U13 ( .A1(1'b1), .A2(n258), .A3(n1153), .A4(n_T_383[28]), .A5(
        n259), .Y(n260) );
  AO221X1_LVT U14 ( .A1(1'b1), .A2(n241), .A3(n1510), .A4(reg_dscratch[26]), 
        .A5(n242), .Y(n244) );
  AO221X1_LVT U15 ( .A1(1'b1), .A2(n224), .A3(n1160), .A4(n_T_444[33]), .A5(
        n228), .Y(n230) );
  AO221X1_LVT U16 ( .A1(1'b1), .A2(n191), .A3(n1487), .A4(reg_stvec[35]), .A5(
        n196), .Y(n201) );
  AO221X1_LVT U17 ( .A1(1'b1), .A2(n1560), .A3(n_T_45[15]), .A4(n1689), .A5(
        n178), .Y(n180) );
  AO221X1_LVT U18 ( .A1(1'b1), .A2(n180), .A3(n1487), .A4(reg_stvec[15]), .A5(
        n181), .Y(n182) );
  AO221X1_LVT U19 ( .A1(1'b1), .A2(n163), .A3(n1153), .A4(n_T_383[25]), .A5(
        n164), .Y(n166) );
  AO221X1_LVT U20 ( .A1(1'b1), .A2(n142), .A3(n1167), .A4(read_fcsr[4]), .A5(
        n143), .Y(n145) );
  AO221X1_LVT U21 ( .A1(1'b1), .A2(n87), .A3(n1508), .A4(reg_sscratch[12]), 
        .A5(n88), .Y(n90) );
  AO221X1_LVT U22 ( .A1(1'b1), .A2(n669), .A3(io_pmp_1_cfg_a[1]), .A4(n1507), 
        .A5(n92), .Y(n93) );
  AO221X1_LVT U23 ( .A1(1'b1), .A2(n93), .A3(n1496), .A4(io_pmp_1_addr[12]), 
        .A5(n94), .Y(n95) );
  AO221X1_LVT U24 ( .A1(1'b1), .A2(n91), .A3(n1153), .A4(n_T_383[12]), .A5(n95), .Y(n96) );
  AO221X1_LVT U25 ( .A1(1'b1), .A2(n71), .A3(n1689), .A4(n_T_45[14]), .A5(n72), 
        .Y(n74) );
  AO221X1_LVT U26 ( .A1(1'b1), .A2(n75), .A3(n1160), .A4(n_T_444[14]), .A5(n76), .Y(n77) );
  AO221X1_LVT U27 ( .A1(1'b1), .A2(n32), .A3(n1160), .A4(n_T_444[22]), .A5(n33), .Y(n35) );
  AO221X1_LVT U28 ( .A1(1'b1), .A2(n37), .A3(n1157), .A4(n1924), .A5(n38), .Y(
        n39) );
  AO221X1_LVT U29 ( .A1(1'b1), .A2(n36), .A3(n1153), .A4(n_T_383[22]), .A5(n39), .Y(n40) );
  AO221X1_LVT U30 ( .A1(1'b1), .A2(n24), .A3(reg_mepc[39]), .A4(n502), .A5(n25), .Y(io_evec[39]) );
  AO221X1_LVT U31 ( .A1(1'b1), .A2(n14), .A3(n1493), .A4(reg_dpc[6]), .A5(n15), 
        .Y(n17) );
  AO221X1_LVT U32 ( .A1(1'b1), .A2(n20), .A3(n1491), .A4(io_pmp_4_addr[6]), 
        .A5(n21), .Y(n22) );
  AO221X1_LVT U33 ( .A1(1'b1), .A2(n2), .A3(n499), .A4(reg_stvec[30]), .A5(n3), 
        .Y(io_evec[30]) );
  IBUFFX2_LVT U34 ( .A(n1204), .Y(n1333) );
  NAND3X0_LVT U35 ( .A1(n1384), .A2(n489), .A3(n1386), .Y(n1) );
  NAND2X0_LVT U36 ( .A1(n1374), .A2(n1), .Y(n1416) );
  AO22X1_LVT U37 ( .A1(reg_sepc[30]), .A2(n500), .A3(reg_dpc[30]), .A4(n1356), 
        .Y(n2) );
  AO22X1_LVT U38 ( .A1(reg_mepc[30]), .A2(n502), .A3(reg_mtvec[30]), .A4(n1333), .Y(n3) );
  HADDX1_LVT U40 ( .A0(n1459), .B0(n_T_45[5]), .SO(n5) );
  AO22X1_LVT U41 ( .A1(n492), .A2(wdata[5]), .A3(n5), .A4(n961), .Y(N1433) );
  AOI22X1_LVT U42 ( .A1(n1495), .A2(n_T_389[6]), .A3(n1488), .A4(
        io_ptbr_ppn[6]), .Y(n6) );
  AOI22X1_LVT U43 ( .A1(n1510), .A2(reg_dscratch[6]), .A3(n1689), .A4(
        n_T_45[6]), .Y(n7) );
  NAND2X0_LVT U44 ( .A1(n1481), .A2(io_bp_0_control_m), .Y(n8) );
  NAND4X0_LVT U45 ( .A1(n6), .A2(n7), .A3(n924), .A4(n8), .Y(n9) );
  AO22X1_LVT U46 ( .A1(n1506), .A2(reg_sepc[6]), .A3(n1478), .A4(reg_stvec[6]), 
        .Y(n10) );
  AO22X1_LVT U47 ( .A1(n1508), .A2(reg_sscratch[6]), .A3(n1160), .A4(
        n_T_444[6]), .Y(n11) );
  AO22X1_LVT U48 ( .A1(n1480), .A2(io_pmp_0_addr[6]), .A3(n1479), .A4(
        io_pmp_7_addr[6]), .Y(n12) );
  NOR4X0_LVT U49 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .Y(n13) );
  AO22X1_LVT U50 ( .A1(n1162), .A2(io_time[6]), .A3(n1496), .A4(
        io_pmp_1_addr[6]), .Y(n14) );
  AO22X1_LVT U51 ( .A1(n1494), .A2(io_pmp_6_addr[6]), .A3(n1470), .A4(
        reg_mtvec[6]), .Y(n15) );
  AO22X1_LVT U53 ( .A1(n1492), .A2(io_pmp_2_addr[6]), .A3(n1469), .A4(
        read_medeleg_6), .Y(n18) );
  AO22X1_LVT U54 ( .A1(n1485), .A2(reg_mscratch[6]), .A3(n1473), .A4(
        io_pmp_3_addr[6]), .Y(n19) );
  AO22X1_LVT U55 ( .A1(n1489), .A2(reg_mepc[6]), .A3(n1490), .A4(
        io_bp_0_address[6]), .Y(n20) );
  AO22X1_LVT U56 ( .A1(n1472), .A2(io_pmp_5_addr[6]), .A3(n1477), .A4(
        io_fcsr_rm[1]), .Y(n21) );
  NOR4X0_LVT U57 ( .A1(n17), .A2(n18), .A3(n19), .A4(n22), .Y(n23) );
  NAND2X0_LVT U58 ( .A1(n13), .A2(n23), .Y(io_rw_rdata[6]) );
  AO22X1_LVT U59 ( .A1(reg_sepc[39]), .A2(n1355), .A3(n1356), .A4(reg_dpc[39]), 
        .Y(n24) );
  INVX0_LVT U60 ( .A(n1357), .Y(n25) );
  AO22X1_LVT U62 ( .A1(n1129), .A2(n_T_44[52]), .A3(wdata[58]), .A4(n1128), 
        .Y(N1549) );
  NAND4X0_LVT U63 ( .A1(n1390), .A2(n1379), .A3(n1417), .A4(io_decode_0_csr[7]), .Y(n27) );
  OR2X1_LVT U64 ( .A1(n1375), .A2(n27), .Y(n1396) );
  NAND3X0_LVT U65 ( .A1(io_pmp_6_cfg_l), .A2(n458), .A3(io_pmp_6_cfg_a[0]), 
        .Y(n28) );
  NAND3X0_LVT U66 ( .A1(n1472), .A2(n437), .A3(n28), .Y(n434) );
  AO222X1_LVT U67 ( .A1(reg_sepc[34]), .A2(n500), .A3(reg_dpc[34]), .A4(n1356), 
        .A5(reg_stvec[34]), .A6(n499), .Y(n29) );
  AO21X1_LVT U68 ( .A1(reg_mepc[34]), .A2(n502), .A3(n29), .Y(io_evec[34]) );
  INVX0_LVT U69 ( .A(io_rw_wdata[58]), .Y(n30) );
  OA222X1_LVT U70 ( .A1(io_rw_wdata[58]), .A2(io_rw_rdata[58]), .A3(
        io_rw_wdata[58]), .A4(n589), .A5(n516), .A6(n30), .Y(wdata[58]) );
  AND2X1_LVT U71 ( .A1(n1194), .A2(n1186), .Y(io_interrupt_cause[0]) );
  AO22X1_LVT U72 ( .A1(n1489), .A2(reg_mepc[22]), .A3(n1496), .A4(
        io_pmp_1_addr[22]), .Y(n31) );
  AO22X1_LVT U73 ( .A1(n1508), .A2(reg_sscratch[22]), .A3(n1473), .A4(
        io_pmp_3_addr[22]), .Y(n32) );
  AO22X1_LVT U74 ( .A1(n1162), .A2(io_time[22]), .A3(n1491), .A4(
        io_pmp_4_addr[22]), .Y(n33) );
  AO222X1_LVT U76 ( .A1(n1689), .A2(n_T_45[22]), .A3(n1487), .A4(reg_stvec[22]), .A5(n1493), .A6(reg_dpc[22]), .Y(n36) );
  AO22X1_LVT U77 ( .A1(n1494), .A2(io_pmp_6_addr[22]), .A3(n1479), .A4(
        io_pmp_7_addr[22]), .Y(n37) );
  AO22X1_LVT U78 ( .A1(n1485), .A2(reg_mscratch[22]), .A3(n1492), .A4(
        io_pmp_2_addr[22]), .Y(n38) );
  AO22X1_LVT U79 ( .A1(n1490), .A2(io_bp_0_address[22]), .A3(n1497), .A4(
        reg_mtvec[22]), .Y(n41) );
  AO22X1_LVT U80 ( .A1(n1510), .A2(reg_dscratch[22]), .A3(n1506), .A4(
        reg_sepc[22]), .Y(n42) );
  AO22X1_LVT U81 ( .A1(n1472), .A2(io_pmp_5_addr[22]), .A3(n1480), .A4(
        io_pmp_0_addr[22]), .Y(n43) );
  OR4X1_LVT U82 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .Y(n44) );
  OR3X1_LVT U83 ( .A1(n31), .A2(n35), .A3(n44), .Y(io_rw_rdata[22]) );
  AO22X1_LVT U84 ( .A1(n1487), .A2(reg_stvec[13]), .A3(n1496), .A4(
        io_pmp_1_addr[13]), .Y(n45) );
  AOI21X1_LVT U85 ( .A1(n_T_45[13]), .A2(n1689), .A3(n1559), .Y(n46) );
  AOI22X1_LVT U86 ( .A1(n1490), .A2(io_bp_0_address[13]), .A3(n1495), .A4(
        n_T_1155[1]), .Y(n47) );
  NAND4X0_LVT U87 ( .A1(n1155), .A2(n46), .A3(n758), .A4(n47), .Y(n48) );
  AO22X1_LVT U88 ( .A1(n1479), .A2(io_pmp_7_addr[13]), .A3(n1473), .A4(
        io_pmp_3_addr[13]), .Y(n49) );
  AO22X1_LVT U89 ( .A1(n1472), .A2(io_pmp_5_addr[13]), .A3(n1488), .A4(
        io_ptbr_ppn[13]), .Y(n50) );
  NOR4X0_LVT U90 ( .A1(n45), .A2(n48), .A3(n49), .A4(n50), .Y(n52) );
  AOI22X1_LVT U91 ( .A1(n1489), .A2(reg_mepc[13]), .A3(n1494), .A4(
        io_pmp_6_addr[13]), .Y(n53) );
  AOI22X1_LVT U92 ( .A1(n1480), .A2(io_pmp_0_addr[13]), .A3(n1469), .A4(
        read_medeleg_13), .Y(n54) );
  AO22X1_LVT U93 ( .A1(n1485), .A2(reg_mscratch[13]), .A3(n1497), .A4(
        reg_mtvec[13]), .Y(n55) );
  AO22X1_LVT U94 ( .A1(n1162), .A2(io_time[13]), .A3(n1491), .A4(
        io_pmp_4_addr[13]), .Y(n56) );
  AO22X1_LVT U95 ( .A1(n1160), .A2(n_T_444[13]), .A3(n1153), .A4(n_T_383[13]), 
        .Y(n57) );
  AO22X1_LVT U96 ( .A1(n1508), .A2(reg_sscratch[13]), .A3(n1492), .A4(
        io_pmp_2_addr[13]), .Y(n58) );
  NOR4X0_LVT U97 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .Y(n59) );
  NAND4X0_LVT U98 ( .A1(n52), .A2(n53), .A3(n54), .A4(n59), .Y(io_rw_rdata[13]) );
  OR3X1_LVT U99 ( .A1(n952), .A2(n950), .A3(n376), .Y(n60) );
  AO221X1_LVT U100 ( .A1(n951), .A2(io_rw_addr[9]), .A3(n951), .A4(n1931), 
        .A5(n60), .Y(n2157) );
  OA21X1_LVT U101 ( .A1(n960), .A2(n_T_45[4]), .A3(n961), .Y(n61) );
  INVX0_LVT U102 ( .A(n1459), .Y(n62) );
  AO22X1_LVT U103 ( .A1(n492), .A2(wdata[4]), .A3(n61), .A4(n62), .Y(N1432) );
  INVX0_LVT U104 ( .A(io_rw_wdata[57]), .Y(n63) );
  OA222X1_LVT U105 ( .A1(io_rw_wdata[57]), .A2(io_rw_rdata[57]), .A3(
        io_rw_wdata[57]), .A4(n589), .A5(n516), .A6(n63), .Y(wdata[57]) );
  AOI22X1_LVT U106 ( .A1(n1479), .A2(io_pmp_7_addr[14]), .A3(n1494), .A4(
        io_pmp_6_addr[14]), .Y(n64) );
  AOI22X1_LVT U107 ( .A1(n1485), .A2(reg_mscratch[14]), .A3(n1493), .A4(
        reg_dpc[14]), .Y(n65) );
  AOI22X1_LVT U108 ( .A1(n1508), .A2(reg_sscratch[14]), .A3(n1497), .A4(
        reg_mtvec[14]), .Y(n66) );
  AO22X1_LVT U109 ( .A1(n1490), .A2(io_bp_0_address[14]), .A3(n1480), .A4(
        io_pmp_0_addr[14]), .Y(n67) );
  AO22X1_LVT U110 ( .A1(n1496), .A2(io_pmp_1_addr[14]), .A3(n1473), .A4(
        io_pmp_3_addr[14]), .Y(n68) );
  AO222X1_LVT U111 ( .A1(n1162), .A2(io_time[14]), .A3(n1492), .A4(
        io_pmp_2_addr[14]), .A5(n1489), .A6(reg_mepc[14]), .Y(n69) );
  AO21X1_LVT U112 ( .A1(io_pmp_4_addr[14]), .A2(n1491), .A3(n1156), .Y(n70) );
  AO21X1_LVT U113 ( .A1(n1487), .A2(reg_stvec[14]), .A3(n70), .Y(n71) );
  AO22X1_LVT U114 ( .A1(n1153), .A2(n_T_383[14]), .A3(n1488), .A4(
        io_ptbr_ppn[14]), .Y(n72) );
  AO21X1_LVT U116 ( .A1(n1510), .A2(reg_dscratch[14]), .A3(n74), .Y(n75) );
  AO22X1_LVT U117 ( .A1(n1506), .A2(reg_sepc[14]), .A3(n1472), .A4(
        io_pmp_5_addr[14]), .Y(n76) );
  NOR4X0_LVT U118 ( .A1(n67), .A2(n68), .A3(n69), .A4(n77), .Y(n78) );
  NAND4X0_LVT U119 ( .A1(n64), .A2(n65), .A3(n66), .A4(n78), .Y(
        io_rw_rdata[14]) );
  HADDX1_LVT U120 ( .A0(n1144), .B0(io_time[3]), .SO(n79) );
  AO22X1_LVT U121 ( .A1(n1149), .A2(wdata[3]), .A3(n79), .A4(n1446), .Y(N1825)
         );
  AOI22X1_LVT U122 ( .A1(n[1930]), .A2(n930), .A3(io_status_prv[0]), .A4(n929), 
        .Y(n80) );
  NAND3X0_LVT U123 ( .A1(n931), .A2(n590), .A3(n80), .Y(N333) );
  INVX0_LVT U124 ( .A(io_rw_wdata[56]), .Y(n81) );
  OA222X1_LVT U125 ( .A1(io_rw_wdata[56]), .A2(io_rw_rdata[56]), .A3(
        io_rw_wdata[56]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n81), .Y(wdata[56]) );
  AND3X1_LVT U126 ( .A1(n1405), .A2(io_decode_0_csr[5]), .A3(n1368), .Y(n1384)
         );
  AND3X1_LVT U127 ( .A1(io_rw_addr[6]), .A2(io_rw_addr[9]), .A3(n1527), .Y(
        n620) );
  AO22X1_LVT U128 ( .A1(n1489), .A2(reg_mepc[12]), .A3(n1494), .A4(
        io_pmp_6_addr[12]), .Y(n82) );
  AO22X1_LVT U129 ( .A1(n1162), .A2(io_time[12]), .A3(n1479), .A4(
        io_pmp_7_addr[12]), .Y(n83) );
  AO22X1_LVT U130 ( .A1(n1480), .A2(io_pmp_0_addr[12]), .A3(n1492), .A4(
        io_pmp_2_addr[12]), .Y(n84) );
  AO22X1_LVT U131 ( .A1(n1493), .A2(reg_dpc[12]), .A3(n1472), .A4(
        io_pmp_5_addr[12]), .Y(n85) );
  AO22X1_LVT U132 ( .A1(n1160), .A2(n_T_444[12]), .A3(n1497), .A4(
        reg_mtvec[12]), .Y(n86) );
  AO22X1_LVT U133 ( .A1(n1490), .A2(io_bp_0_address[12]), .A3(n1491), .A4(
        io_pmp_4_addr[12]), .Y(n87) );
  AO22X1_LVT U134 ( .A1(n1510), .A2(reg_dscratch[12]), .A3(n1488), .A4(
        io_ptbr_ppn[12]), .Y(n88) );
  AO22X1_LVT U136 ( .A1(n1506), .A2(reg_sepc[12]), .A3(n1473), .A4(
        io_pmp_3_addr[12]), .Y(n91) );
  AO22X1_LVT U137 ( .A1(n1481), .A2(io_bp_0_control_action), .A3(n1452), .A4(
        io_status_isa_12_), .Y(n92) );
  AO22X1_LVT U138 ( .A1(n1485), .A2(reg_mscratch[12]), .A3(n1157), .A4(n[1929]), .Y(n94) );
  OR3X1_LVT U139 ( .A1(n86), .A2(n90), .A3(n96), .Y(n97) );
  OR3X1_LVT U140 ( .A1(n84), .A2(n85), .A3(n97), .Y(n98) );
  OR3X1_LVT U141 ( .A1(n82), .A2(n83), .A3(n98), .Y(io_rw_rdata[12]) );
  INVX0_LVT U142 ( .A(n879), .Y(n99) );
  INVX0_LVT U143 ( .A(wdata[9]), .Y(n100) );
  OA222X1_LVT U144 ( .A1(n99), .A2(n1912), .A3(n99), .A4(n590), .A5(n879), 
        .A6(n100), .Y(n1911) );
  INVX0_LVT U145 ( .A(io_rw_wdata[3]), .Y(n101) );
  OA222X1_LVT U146 ( .A1(io_rw_wdata[3]), .A2(n589), .A3(io_rw_wdata[3]), .A4(
        io_rw_rdata[3]), .A5(n516), .A6(n101), .Y(wdata[3]) );
  INVX0_LVT U147 ( .A(io_rw_wdata[59]), .Y(n102) );
  OA222X1_LVT U148 ( .A1(io_rw_wdata[59]), .A2(io_rw_rdata[59]), .A3(
        io_rw_wdata[59]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n102), .Y(
        wdata[59]) );
  INVX0_LVT U149 ( .A(io_rw_wdata[51]), .Y(n103) );
  OA222X1_LVT U150 ( .A1(io_rw_wdata[51]), .A2(io_rw_rdata[51]), .A3(
        io_rw_wdata[51]), .A4(n589), .A5(n516), .A6(n103), .Y(wdata[51]) );
  NAND2X0_LVT U151 ( .A1(n860), .A2(n1442), .Y(n104) );
  OA21X1_LVT U152 ( .A1(io_retire), .A2(n104), .A3(io_singleStep), .Y(N435) );
  INVX0_LVT U153 ( .A(n1378), .Y(n105) );
  NAND3X0_LVT U154 ( .A1(n1405), .A2(io_decode_0_csr[8]), .A3(n105), .Y(n1375)
         );
  AOI22X1_LVT U155 ( .A1(n1487), .A2(reg_stvec[12]), .A3(n1469), .A4(
        read_medeleg_12), .Y(n106) );
  AOI22X1_LVT U156 ( .A1(n1689), .A2(n_T_45[12]), .A3(n1495), .A4(n_T_1155[0]), 
        .Y(n107) );
  NAND3X0_LVT U157 ( .A1(n1083), .A2(n106), .A3(n107), .Y(n669) );
  NAND3X0_LVT U158 ( .A1(io_pmp_4_cfg_l), .A2(n464), .A3(io_pmp_4_cfg_a[0]), 
        .Y(n108) );
  NAND3X0_LVT U159 ( .A1(n1473), .A2(n443), .A3(n108), .Y(n436) );
  INVX0_LVT U160 ( .A(n1175), .Y(n109) );
  AO22X1_LVT U161 ( .A1(n1179), .A2(n1178), .A3(n1190), .A4(n109), .Y(n110) );
  NAND4X0_LVT U162 ( .A1(n1185), .A2(n1192), .A3(n1174), .A4(n110), .Y(n111)
         );
  OR2X1_LVT U163 ( .A1(n1191), .A2(n111), .Y(n1194) );
  INVX0_LVT U164 ( .A(io_rw_wdata[11]), .Y(n112) );
  OA222X1_LVT U165 ( .A1(io_rw_wdata[11]), .A2(n589), .A3(io_rw_wdata[11]), 
        .A4(io_rw_rdata[11]), .A5(n516), .A6(n112), .Y(wdata[11]) );
  INVX0_LVT U166 ( .A(io_rw_wdata[60]), .Y(n113) );
  OA222X1_LVT U167 ( .A1(io_rw_wdata[60]), .A2(n589), .A3(io_rw_wdata[60]), 
        .A4(io_rw_rdata[60]), .A5(n516), .A6(n113), .Y(wdata[60]) );
  INVX0_LVT U168 ( .A(io_rw_wdata[52]), .Y(n114) );
  OA222X1_LVT U169 ( .A1(io_rw_wdata[52]), .A2(io_rw_rdata[52]), .A3(
        io_rw_wdata[52]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n114), .Y(
        wdata[52]) );
  HADDX1_LVT U170 ( .A0(io_retire), .B0(n_T_45[0]), .SO(n115) );
  AO22X1_LVT U171 ( .A1(n492), .A2(wdata[0]), .A3(n115), .A4(n961), .Y(N1428)
         );
  INVX0_LVT U172 ( .A(n1375), .Y(n116) );
  NAND3X0_LVT U173 ( .A1(io_decode_0_csr[6]), .A2(n1386), .A3(n116), .Y(n1426)
         );
  NAND3X0_LVT U174 ( .A1(io_pmp_3_cfg_a[0]), .A2(n460), .A3(io_pmp_3_cfg_l), 
        .Y(n117) );
  NAND3X0_LVT U175 ( .A1(n1492), .A2(n441), .A3(n117), .Y(n432) );
  NAND3X0_LVT U176 ( .A1(io_pmp_7_cfg_l), .A2(n459), .A3(io_pmp_7_cfg_a[0]), 
        .Y(n118) );
  NAND3X0_LVT U177 ( .A1(n1494), .A2(n439), .A3(n118), .Y(n435) );
  NAND3X0_LVT U178 ( .A1(io_pmp_5_cfg_a[0]), .A2(n461), .A3(io_pmp_5_cfg_l), 
        .Y(n119) );
  NAND3X0_LVT U179 ( .A1(n1491), .A2(n438), .A3(n119), .Y(n433) );
  NAND3X0_LVT U180 ( .A1(io_pmp_1_cfg_a[0]), .A2(n462), .A3(io_pmp_1_cfg_l), 
        .Y(n120) );
  NAND3X0_LVT U181 ( .A1(n1480), .A2(n453), .A3(n120), .Y(n430) );
  AO222X1_LVT U182 ( .A1(n500), .A2(reg_sepc[36]), .A3(n499), .A4(
        reg_stvec[36]), .A5(n1356), .A6(reg_dpc[36]), .Y(n121) );
  AO21X1_LVT U183 ( .A1(n502), .A2(reg_mepc[36]), .A3(n121), .Y(io_evec[36])
         );
  AND3X1_LVT U184 ( .A1(n1516), .A2(n1505), .A3(n1527), .Y(n1504) );
  AO22X1_LVT U185 ( .A1(n497), .A2(n_T_52[32]), .A3(wdata[38]), .A4(n1149), 
        .Y(N1923) );
  AO22X1_LVT U186 ( .A1(n494), .A2(n_T_44[44]), .A3(wdata[50]), .A4(n1128), 
        .Y(N1541) );
  AND2X1_LVT U187 ( .A1(io_bp_0_control_action), .A2(n589), .Y(n122) );
  INVX0_LVT U188 ( .A(io_rw_wdata[12]), .Y(n123) );
  OA221X1_LVT U189 ( .A1(io_rw_wdata[12]), .A2(n122), .A3(n123), .A4(n516), 
        .A5(n1482), .Y(N485) );
  AND3X1_LVT U190 ( .A1(io_time[3]), .A2(io_time[4]), .A3(n1144), .Y(n1147) );
  AND3X1_LVT U191 ( .A1(n1516), .A2(n1512), .A3(n1527), .Y(n1154) );
  OA21X1_LVT U192 ( .A1(n959), .A2(n_T_45[3]), .A3(n961), .Y(n124) );
  INVX0_LVT U193 ( .A(n960), .Y(n125) );
  AO22X1_LVT U194 ( .A1(n492), .A2(wdata[3]), .A3(n124), .A4(n125), .Y(N1431)
         );
  INVX0_LVT U195 ( .A(io_rw_wdata[63]), .Y(n126) );
  OA222X1_LVT U196 ( .A1(io_rw_wdata[63]), .A2(io_rw_rdata[63]), .A3(
        io_rw_wdata[63]), .A4(n589), .A5(n516), .A6(n126), .Y(wdata[63]) );
  INVX0_LVT U197 ( .A(io_rw_wdata[50]), .Y(n127) );
  OA222X1_LVT U198 ( .A1(io_rw_wdata[50]), .A2(io_rw_rdata[50]), .A3(
        io_rw_wdata[50]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n127), .Y(
        wdata[50]) );
  INVX0_LVT U199 ( .A(n1500), .Y(n128) );
  INVX0_LVT U200 ( .A(wdata[0]), .Y(n129) );
  OAI222X1_LVT U201 ( .A1(n128), .A2(n954), .A3(n129), .A4(n1455), .A5(n953), 
        .A6(n1697), .Y(N1270) );
  INVX0_LVT U202 ( .A(n1907), .Y(n130) );
  OA222X1_LVT U203 ( .A1(n130), .A2(io_rw_rdata[9]), .A3(n130), .A4(n589), 
        .A5(n516), .A6(n1907), .Y(wdata[9]) );
  AOI22X1_LVT U204 ( .A1(n1492), .A2(io_pmp_2_addr[4]), .A3(n1494), .A4(
        io_pmp_6_addr[4]), .Y(n131) );
  AO22X1_LVT U205 ( .A1(n1168), .A2(reg_scause[4]), .A3(n1478), .A4(
        reg_stvec[4]), .Y(n132) );
  AO22X1_LVT U206 ( .A1(n1162), .A2(io_time[4]), .A3(n1491), .A4(
        io_pmp_4_addr[4]), .Y(n133) );
  AO22X1_LVT U207 ( .A1(n1493), .A2(reg_dpc[4]), .A3(n1480), .A4(
        io_pmp_0_addr[4]), .Y(n134) );
  AO22X1_LVT U208 ( .A1(n1485), .A2(reg_mscratch[4]), .A3(n1469), .A4(
        read_medeleg[4]), .Y(n135) );
  NOR4X0_LVT U209 ( .A1(n132), .A2(n133), .A3(n134), .A4(n135), .Y(n136) );
  AO22X1_LVT U210 ( .A1(n1473), .A2(io_pmp_3_addr[4]), .A3(n1488), .A4(
        io_ptbr_ppn[4]), .Y(n137) );
  AO22X1_LVT U211 ( .A1(n1490), .A2(io_bp_0_address[4]), .A3(n1479), .A4(
        io_pmp_7_addr[4]), .Y(n138) );
  AO22X1_LVT U212 ( .A1(n1508), .A2(reg_sscratch[4]), .A3(n1472), .A4(
        io_pmp_5_addr[4]), .Y(n139) );
  AO22X1_LVT U213 ( .A1(n1160), .A2(n_T_444[4]), .A3(n1153), .A4(n_T_383[4]), 
        .Y(n140) );
  AO22X1_LVT U214 ( .A1(n1489), .A2(reg_mepc[4]), .A3(n1496), .A4(
        io_pmp_1_addr[4]), .Y(n141) );
  AO222X1_LVT U215 ( .A1(n1510), .A2(reg_dscratch[4]), .A3(n1507), .A4(
        io_pmp_0_cfg_a[1]), .A5(n_T_45[4]), .A6(n1689), .Y(n142) );
  AO22X1_LVT U216 ( .A1(n1506), .A2(reg_sepc[4]), .A3(n1481), .A4(
        io_bp_0_control_s), .Y(n143) );
  OR3X1_LVT U218 ( .A1(n140), .A2(n141), .A3(n145), .Y(n146) );
  NOR4X0_LVT U219 ( .A1(n137), .A2(n138), .A3(n139), .A4(n146), .Y(n147) );
  NAND2X0_LVT U220 ( .A1(n1470), .A2(reg_mtvec[4]), .Y(n148) );
  NAND4X0_LVT U221 ( .A1(n131), .A2(n136), .A3(n147), .A4(n148), .Y(
        io_rw_rdata[4]) );
  INVX0_LVT U222 ( .A(n1183), .Y(n149) );
  AND2X1_LVT U223 ( .A1(n149), .A2(n1176), .Y(n1180) );
  AO21X1_LVT U224 ( .A1(read_mideleg_9_), .A2(n1504), .A3(n1502), .Y(n150) );
  INVX0_LVT U225 ( .A(n742), .Y(n151) );
  AO22X1_LVT U226 ( .A1(wdata[9]), .A2(n150), .A3(n446), .A4(n151), .Y(N615)
         );
  INVX0_LVT U227 ( .A(io_rw_wdata[49]), .Y(n152) );
  OA222X1_LVT U228 ( .A1(io_rw_wdata[49]), .A2(io_rw_rdata[49]), .A3(
        io_rw_wdata[49]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n152), .Y(
        wdata[49]) );
  INVX0_LVT U229 ( .A(io_rw_wdata[39]), .Y(n153) );
  OA222X1_LVT U230 ( .A1(io_rw_wdata[39]), .A2(io_rw_rdata[39]), .A3(
        io_rw_wdata[39]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n153), .Y(
        wdata[39]) );
  AND2X1_LVT U231 ( .A1(io_status_prv[0]), .A2(n501), .Y(n154) );
  AO22X1_LVT U232 ( .A1(n1443), .A2(n154), .A3(n949), .A4(wdata[8]), .Y(n1913)
         );
  AOI222X1_LVT U233 ( .A1(n1489), .A2(reg_mepc[25]), .A3(n1506), .A4(
        reg_sepc[25]), .A5(n1491), .A6(io_pmp_4_addr[25]), .Y(n155) );
  AOI22X1_LVT U234 ( .A1(n1162), .A2(io_time[25]), .A3(n1494), .A4(
        io_pmp_6_addr[25]), .Y(n156) );
  AOI22X1_LVT U235 ( .A1(n1508), .A2(reg_sscratch[25]), .A3(n1485), .A4(
        reg_mscratch[25]), .Y(n157) );
  AO22X1_LVT U236 ( .A1(n1492), .A2(io_pmp_2_addr[25]), .A3(n1480), .A4(
        io_pmp_0_addr[25]), .Y(n158) );
  AO22X1_LVT U237 ( .A1(n1490), .A2(io_bp_0_address[25]), .A3(n1479), .A4(
        io_pmp_7_addr[25]), .Y(n159) );
  AO222X1_LVT U238 ( .A1(n1507), .A2(io_pmp_3_cfg_w), .A3(n1496), .A4(
        io_pmp_1_addr[25]), .A5(n1160), .A6(n_T_444[25]), .Y(n160) );
  AO222X1_LVT U239 ( .A1(n1689), .A2(n_T_45[25]), .A3(n1497), .A4(
        reg_mtvec[25]), .A5(reg_dpc[25]), .A6(n1493), .Y(n161) );
  AO21X1_LVT U240 ( .A1(n1510), .A2(reg_dscratch[25]), .A3(n161), .Y(n162) );
  AO21X1_LVT U241 ( .A1(n1487), .A2(reg_stvec[25]), .A3(n162), .Y(n163) );
  AO22X1_LVT U242 ( .A1(n1472), .A2(io_pmp_5_addr[25]), .A3(n1473), .A4(
        io_pmp_3_addr[25]), .Y(n164) );
  NOR4X0_LVT U244 ( .A1(n158), .A2(n159), .A3(n160), .A4(n166), .Y(n167) );
  NAND4X0_LVT U245 ( .A1(n155), .A2(n156), .A3(n157), .A4(n167), .Y(
        io_rw_rdata[25]) );
  INVX0_LVT U246 ( .A(io_csr_stall), .Y(n168) );
  INVX0_LVT U247 ( .A(n1142), .Y(n169) );
  OA221X1_LVT U248 ( .A1(io_time[1]), .A2(io_time[0]), .A3(io_time[1]), .A4(
        n168), .A5(n169), .Y(n170) );
  AO22X1_LVT U249 ( .A1(n1446), .A2(n170), .A3(wdata[1]), .A4(n1149), .Y(N1823) );
  AO22X1_LVT U250 ( .A1(n494), .A2(n_T_44[32]), .A3(wdata[38]), .A4(n1128), 
        .Y(N1529) );
  INVX0_LVT U251 ( .A(io_rw_wdata[48]), .Y(n171) );
  OA222X1_LVT U252 ( .A1(io_rw_wdata[48]), .A2(io_rw_rdata[48]), .A3(
        io_rw_wdata[48]), .A4(n589), .A5(n516), .A6(n171), .Y(wdata[48]) );
  INVX0_LVT U253 ( .A(io_rw_wdata[62]), .Y(n172) );
  OA222X1_LVT U254 ( .A1(io_rw_wdata[62]), .A2(n589), .A3(io_rw_wdata[62]), 
        .A4(io_rw_rdata[62]), .A5(n516), .A6(n172), .Y(wdata[62]) );
  AOI22X1_LVT U255 ( .A1(n[1929]), .A2(n930), .A3(io_status_prv[1]), .A4(n929), 
        .Y(n173) );
  OR2X1_LVT U256 ( .A1(n931), .A2(n367), .Y(n174) );
  NAND3X0_LVT U257 ( .A1(n174), .A2(n590), .A3(n173), .Y(N334) );
  AO222X1_LVT U258 ( .A1(n1160), .A2(n_T_444[15]), .A3(n1480), .A4(
        io_pmp_0_addr[15]), .A5(io_pmp_5_addr[15]), .A6(n1472), .Y(n175) );
  AO22X1_LVT U259 ( .A1(n1491), .A2(io_pmp_4_addr[15]), .A3(n1492), .A4(
        io_pmp_2_addr[15]), .Y(n176) );
  AOI22X1_LVT U260 ( .A1(n1495), .A2(n_T_1155_3), .A3(n1488), .A4(
        io_ptbr_ppn[15]), .Y(n177) );
  NAND3X0_LVT U261 ( .A1(n177), .A2(n631), .A3(n632), .Y(n178) );
  AO22X1_LVT U263 ( .A1(n1162), .A2(io_time[15]), .A3(n1490), .A4(
        io_bp_0_address[15]), .Y(n181) );
  AO22X1_LVT U264 ( .A1(n1496), .A2(io_pmp_1_addr[15]), .A3(n1473), .A4(
        io_pmp_3_addr[15]), .Y(n183) );
  NOR4X0_LVT U265 ( .A1(n175), .A2(n176), .A3(n182), .A4(n183), .Y(n184) );
  AO22X1_LVT U266 ( .A1(n1153), .A2(n_T_383[15]), .A3(n1494), .A4(
        io_pmp_6_addr[15]), .Y(n185) );
  AO22X1_LVT U267 ( .A1(n1489), .A2(reg_mepc[15]), .A3(n1497), .A4(
        reg_mtvec[15]), .Y(n186) );
  AO22X1_LVT U268 ( .A1(n1508), .A2(reg_sscratch[15]), .A3(n1479), .A4(
        io_pmp_7_addr[15]), .Y(n187) );
  AO22X1_LVT U269 ( .A1(n1510), .A2(reg_dscratch[15]), .A3(n1485), .A4(
        reg_mscratch[15]), .Y(n188) );
  NOR4X0_LVT U270 ( .A1(n185), .A2(n186), .A3(n187), .A4(n188), .Y(n189) );
  NAND2X0_LVT U271 ( .A1(n184), .A2(n189), .Y(io_rw_rdata[15]) );
  AO222X1_LVT U272 ( .A1(n1485), .A2(reg_mscratch[35]), .A3(n1489), .A4(
        reg_mepc[35]), .A5(n_T_444[35]), .A6(n1160), .Y(n190) );
  AO22X1_LVT U273 ( .A1(n1162), .A2(n1964), .A3(n1153), .A4(n_T_383[35]), .Y(
        n191) );
  AOI22X1_LVT U274 ( .A1(n1510), .A2(reg_dscratch[35]), .A3(n1689), .A4(
        n_T_45[35]), .Y(n192) );
  AOI22X1_LVT U275 ( .A1(n1507), .A2(io_pmp_4_cfg_a[0]), .A3(n1490), .A4(
        io_bp_0_address[35]), .Y(n193) );
  NAND2X0_LVT U276 ( .A1(n1493), .A2(reg_dpc[35]), .Y(n195) );
  NAND4X0_LVT U277 ( .A1(n192), .A2(n1041), .A3(n193), .A4(n195), .Y(n196) );
  AO22X1_LVT U279 ( .A1(n1508), .A2(reg_sscratch[35]), .A3(n1506), .A4(
        reg_sepc[35]), .Y(n202) );
  OR3X1_LVT U280 ( .A1(n190), .A2(n201), .A3(n202), .Y(io_rw_rdata[35]) );
  AND3X1_LVT U281 ( .A1(io_rw_addr[6]), .A2(n1515), .A3(n1527), .Y(n1509) );
  INVX0_LVT U282 ( .A(io_rw_wdata[25]), .Y(n203) );
  OA222X1_LVT U283 ( .A1(io_rw_wdata[25]), .A2(io_rw_rdata[25]), .A3(
        io_rw_wdata[25]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n203), .Y(
        wdata[25]) );
  AO22X1_LVT U284 ( .A1(n497), .A2(n_T_52[44]), .A3(wdata[50]), .A4(n1149), 
        .Y(N1935) );
  INVX0_LVT U285 ( .A(io_rw_wdata[41]), .Y(n204) );
  OA222X1_LVT U286 ( .A1(io_rw_wdata[41]), .A2(io_rw_rdata[41]), .A3(
        io_rw_wdata[41]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n204), .Y(
        wdata[41]) );
  INVX0_LVT U287 ( .A(io_rw_wdata[44]), .Y(n205) );
  OA222X1_LVT U288 ( .A1(io_rw_wdata[44]), .A2(io_rw_rdata[44]), .A3(
        io_rw_wdata[44]), .A4(n589), .A5(n516), .A6(n205), .Y(wdata[44]) );
  INVX0_LVT U289 ( .A(n1498), .Y(n206) );
  OAI22X1_LVT U290 ( .A1(n701), .A2(n1483), .A3(n899), .A4(n206), .Y(N883) );
  AO21X1_LVT U291 ( .A1(n1191), .A2(n1190), .A3(n1189), .Y(n207) );
  NAND3X0_LVT U292 ( .A1(n1192), .A2(n1193), .A3(n207), .Y(n208) );
  OR2X1_LVT U293 ( .A1(n1187), .A2(n1188), .Y(n209) );
  NAND3X0_LVT U294 ( .A1(n209), .A2(n208), .A3(n1186), .Y(
        io_interrupt_cause[3]) );
  AO22X1_LVT U295 ( .A1(n1491), .A2(io_pmp_4_addr[10]), .A3(n1479), .A4(
        io_pmp_7_addr[10]), .Y(n210) );
  AO22X1_LVT U296 ( .A1(n1507), .A2(io_pmp_1_cfg_x), .A3(n1506), .A4(
        reg_sepc[10]), .Y(n211) );
  AO22X1_LVT U297 ( .A1(n1162), .A2(io_time[10]), .A3(n1472), .A4(
        io_pmp_5_addr[10]), .Y(n212) );
  AO22X1_LVT U298 ( .A1(n1510), .A2(reg_dscratch[10]), .A3(n1493), .A4(
        reg_dpc[10]), .Y(n213) );
  NOR4X0_LVT U299 ( .A1(n210), .A2(n211), .A3(n212), .A4(n213), .Y(n214) );
  AO22X1_LVT U300 ( .A1(n1689), .A2(n_T_45[10]), .A3(n1153), .A4(n_T_383[10]), 
        .Y(n215) );
  AO222X1_LVT U301 ( .A1(n1489), .A2(reg_mepc[10]), .A3(n1473), .A4(
        io_pmp_3_addr[10]), .A5(io_pmp_1_addr[10]), .A6(n1496), .Y(n216) );
  AO22X1_LVT U302 ( .A1(n1480), .A2(io_pmp_0_addr[10]), .A3(n1494), .A4(
        io_pmp_6_addr[10]), .Y(n217) );
  AO222X1_LVT U303 ( .A1(n1485), .A2(reg_mscratch[10]), .A3(n488), .A4(
        io_ptbr_ppn[10]), .A5(n1160), .A6(n_T_444[10]), .Y(n218) );
  NOR4X0_LVT U304 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .Y(n219) );
  AOI22X1_LVT U305 ( .A1(n1490), .A2(io_bp_0_address[10]), .A3(n1492), .A4(
        io_pmp_2_addr[10]), .Y(n220) );
  AO22X1_LVT U306 ( .A1(n1508), .A2(reg_sscratch[10]), .A3(n1497), .A4(
        reg_mtvec[10]), .Y(n221) );
  AOI21X1_LVT U307 ( .A1(n1487), .A2(reg_stvec[10]), .A3(n221), .Y(n222) );
  NAND4X0_LVT U308 ( .A1(n214), .A2(n219), .A3(n220), .A4(n222), .Y(
        io_rw_rdata[10]) );
  AO22X1_LVT U309 ( .A1(n1485), .A2(reg_mscratch[33]), .A3(n1489), .A4(
        reg_mepc[33]), .Y(n223) );
  AO22X1_LVT U310 ( .A1(n1162), .A2(n1966), .A3(n1506), .A4(reg_sepc[33]), .Y(
        n224) );
  AOI22X1_LVT U311 ( .A1(n1510), .A2(reg_dscratch[33]), .A3(n1689), .A4(
        n_T_45[33]), .Y(n225) );
  AOI22X1_LVT U312 ( .A1(n1493), .A2(reg_dpc[33]), .A3(n1490), .A4(
        io_bp_0_address[33]), .Y(n226) );
  AOI22X1_LVT U313 ( .A1(n1153), .A2(n_T_383[33]), .A3(n1487), .A4(
        reg_stvec[33]), .Y(n227) );
  NAND4X0_LVT U314 ( .A1(n1026), .A2(n225), .A3(n226), .A4(n227), .Y(n228) );
  AO22X1_LVT U316 ( .A1(n1508), .A2(reg_sscratch[33]), .A3(n1507), .A4(
        io_pmp_4_cfg_w), .Y(n231) );
  OR3X1_LVT U317 ( .A1(n223), .A2(n230), .A3(n231), .Y(io_rw_rdata[33]) );
  INVX0_LVT U318 ( .A(n1904), .Y(n232) );
  OA222X1_LVT U319 ( .A1(n232), .A2(io_rw_cmd[1]), .A3(n232), .A4(
        io_rw_rdata[5]), .A5(n516), .A6(n1904), .Y(wdata[5]) );
  INVX0_LVT U320 ( .A(io_rw_wdata[40]), .Y(n233) );
  OA222X1_LVT U321 ( .A1(io_rw_wdata[40]), .A2(io_rw_rdata[40]), .A3(
        io_rw_wdata[40]), .A4(n589), .A5(n516), .A6(n233), .Y(wdata[40]) );
  INVX0_LVT U322 ( .A(io_rw_wdata[45]), .Y(n234) );
  OA222X1_LVT U323 ( .A1(io_rw_wdata[45]), .A2(io_rw_rdata[45]), .A3(
        io_rw_wdata[45]), .A4(n589), .A5(n516), .A6(n234), .Y(wdata[45]) );
  AO222X1_LVT U324 ( .A1(n1508), .A2(reg_sscratch[26]), .A3(n1480), .A4(
        io_pmp_0_addr[26]), .A5(n1160), .A6(n_T_444[26]), .Y(n235) );
  AO22X1_LVT U325 ( .A1(n1485), .A2(reg_mscratch[26]), .A3(n1491), .A4(
        io_pmp_4_addr[26]), .Y(n236) );
  AO22X1_LVT U326 ( .A1(n1494), .A2(io_pmp_6_addr[26]), .A3(n1473), .A4(
        io_pmp_3_addr[26]), .Y(n237) );
  AO22X1_LVT U327 ( .A1(n1507), .A2(io_pmp_3_cfg_x), .A3(n1472), .A4(
        io_pmp_5_addr[26]), .Y(n238) );
  NOR4X0_LVT U328 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .Y(n239) );
  AO222X1_LVT U329 ( .A1(n1489), .A2(reg_mepc[26]), .A3(n1492), .A4(
        io_pmp_2_addr[26]), .A5(n1487), .A6(reg_stvec[26]), .Y(n240) );
  AO222X1_LVT U330 ( .A1(n1689), .A2(n_T_45[26]), .A3(n1497), .A4(
        reg_mtvec[26]), .A5(reg_dpc[26]), .A6(n1493), .Y(n241) );
  AO22X1_LVT U331 ( .A1(n1153), .A2(n_T_383[26]), .A3(n1479), .A4(
        io_pmp_7_addr[26]), .Y(n242) );
  AO22X1_LVT U333 ( .A1(n1162), .A2(io_time[26]), .A3(n1496), .A4(
        io_pmp_1_addr[26]), .Y(n245) );
  AO22X1_LVT U334 ( .A1(n1506), .A2(reg_sepc[26]), .A3(n1490), .A4(
        io_bp_0_address[26]), .Y(n246) );
  NOR4X0_LVT U335 ( .A1(n240), .A2(n244), .A3(n245), .A4(n246), .Y(n247) );
  NAND2X0_LVT U336 ( .A1(n239), .A2(n247), .Y(io_rw_rdata[26]) );
  AOI22X1_LVT U337 ( .A1(n1494), .A2(io_pmp_6_addr[28]), .A3(n1497), .A4(
        reg_mtvec[28]), .Y(n248) );
  AOI22X1_LVT U338 ( .A1(n1496), .A2(io_pmp_1_addr[28]), .A3(n1492), .A4(
        io_pmp_2_addr[28]), .Y(n249) );
  AOI22X1_LVT U339 ( .A1(n1485), .A2(reg_mscratch[28]), .A3(n1487), .A4(
        reg_stvec[28]), .Y(n250) );
  AO22X1_LVT U340 ( .A1(n1508), .A2(reg_sscratch[28]), .A3(n1480), .A4(
        io_pmp_0_addr[28]), .Y(n251) );
  AO22X1_LVT U341 ( .A1(n1510), .A2(reg_dscratch[28]), .A3(n1491), .A4(
        io_pmp_4_addr[28]), .Y(n252) );
  AO22X1_LVT U342 ( .A1(n1472), .A2(io_pmp_5_addr[28]), .A3(n1473), .A4(
        io_pmp_3_addr[28]), .Y(n253) );
  AO222X1_LVT U343 ( .A1(n1689), .A2(n_T_45[28]), .A3(n1506), .A4(reg_sepc[28]), .A5(n1489), .A6(reg_mepc[28]), .Y(n254) );
  AO21X1_LVT U344 ( .A1(n1493), .A2(reg_dpc[28]), .A3(n254), .Y(n255) );
  AO22X1_LVT U345 ( .A1(n1490), .A2(io_bp_0_address[28]), .A3(n1479), .A4(
        io_pmp_7_addr[28]), .Y(n256) );
  AO22X1_LVT U347 ( .A1(n1162), .A2(io_time[28]), .A3(n1160), .A4(n_T_444[28]), 
        .Y(n259) );
  NOR4X0_LVT U348 ( .A1(n251), .A2(n252), .A3(n253), .A4(n260), .Y(n261) );
  NAND4X0_LVT U349 ( .A1(n248), .A2(n249), .A3(n250), .A4(n261), .Y(
        io_rw_rdata[28]) );
  AO22X1_LVT U350 ( .A1(n1160), .A2(n_T_444[31]), .A3(n1153), .A4(n_T_383[31]), 
        .Y(n262) );
  AO22X1_LVT U351 ( .A1(n1490), .A2(io_bp_0_address[31]), .A3(n1487), .A4(
        reg_stvec[31]), .Y(n263) );
  AO22X1_LVT U352 ( .A1(n1489), .A2(reg_mepc[31]), .A3(n1506), .A4(
        reg_sepc[31]), .Y(n264) );
  AO22X1_LVT U353 ( .A1(n1493), .A2(reg_dpc[31]), .A3(n1497), .A4(
        reg_mtvec[31]), .Y(n265) );
  AO22X1_LVT U355 ( .A1(n1508), .A2(reg_sscratch[31]), .A3(n1162), .A4(
        io_time[31]), .Y(n268) );
  AND4X1_LVT U356 ( .A1(io_rw_addr[0]), .A2(io_rw_addr[1]), .A3(n616), .A4(
        io_rw_addr[2]), .Y(n1479) );
  NAND2X0_LVT U357 ( .A1(wdata[5]), .A2(n949), .Y(n271) );
  NAND2X0_LVT U358 ( .A1(n1935), .A2(n1443), .Y(n272) );
  NAND3X0_LVT U359 ( .A1(n271), .A2(n917), .A3(n272), .Y(n1914) );
  INVX0_LVT U360 ( .A(io_rw_wdata[17]), .Y(n273) );
  OA222X1_LVT U361 ( .A1(io_rw_wdata[17]), .A2(n589), .A3(io_rw_wdata[17]), 
        .A4(io_rw_rdata[17]), .A5(n516), .A6(n273), .Y(wdata[17]) );
  AO22X1_LVT U362 ( .A1(n497), .A2(n_T_52[52]), .A3(wdata[58]), .A4(n1149), 
        .Y(N1943) );
  INVX0_LVT U363 ( .A(io_rw_wdata[55]), .Y(n274) );
  OA222X1_LVT U364 ( .A1(io_rw_wdata[55]), .A2(io_rw_rdata[55]), .A3(
        io_rw_wdata[55]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n274), .Y(
        wdata[55]) );
  INVX0_LVT U365 ( .A(io_rw_wdata[42]), .Y(n275) );
  OA222X1_LVT U366 ( .A1(io_rw_wdata[42]), .A2(io_rw_rdata[42]), .A3(
        io_rw_wdata[42]), .A4(n589), .A5(n516), .A6(n275), .Y(wdata[42]) );
  INVX0_LVT U367 ( .A(io_rw_wdata[53]), .Y(n276) );
  OA222X1_LVT U368 ( .A1(io_rw_wdata[53]), .A2(io_rw_rdata[53]), .A3(
        io_rw_wdata[53]), .A4(n589), .A5(n516), .A6(n276), .Y(wdata[53]) );
  AO22X1_LVT U369 ( .A1(n1689), .A2(n_T_45[38]), .A3(n1493), .A4(reg_dpc[38]), 
        .Y(n277) );
  AO22X1_LVT U370 ( .A1(n1506), .A2(reg_sepc[38]), .A3(n1153), .A4(n_T_383[38]), .Y(n278) );
  AO22X1_LVT U372 ( .A1(n1510), .A2(reg_dscratch[38]), .A3(n1508), .A4(
        reg_sscratch[38]), .Y(n281) );
  AO22X1_LVT U373 ( .A1(n1160), .A2(n_T_444[38]), .A3(n1489), .A4(reg_mepc[38]), .Y(n282) );
  OR3X1_LVT U374 ( .A1(n280), .A2(n281), .A3(n283), .Y(io_rw_rdata[38]) );
  AOI22X1_LVT U375 ( .A1(n1473), .A2(io_pmp_3_addr[8]), .A3(n1481), .A4(
        io_bp_0_control_tmatch[1]), .Y(n284) );
  NAND2X0_LVT U376 ( .A1(io_ptbr_ppn[8]), .A2(n1488), .Y(n285) );
  NAND3X0_LVT U377 ( .A1(n285), .A2(n948), .A3(n947), .Y(n286) );
  AO22X1_LVT U379 ( .A1(n1487), .A2(reg_stvec[8]), .A3(n1154), .A4(n1931), .Y(
        n289) );
  AO22X1_LVT U380 ( .A1(n1153), .A2(n_T_383[8]), .A3(n1452), .A4(n1922), .Y(
        n290) );
  AO22X1_LVT U381 ( .A1(n1160), .A2(n_T_444[8]), .A3(n1469), .A4(
        read_medeleg_8), .Y(n291) );
  NOR4X0_LVT U382 ( .A1(n288), .A2(n289), .A3(n290), .A4(n291), .Y(n292) );
  AO22X1_LVT U383 ( .A1(n1496), .A2(io_pmp_1_addr[8]), .A3(n1491), .A4(
        io_pmp_4_addr[8]), .Y(n293) );
  AO22X1_LVT U384 ( .A1(n1162), .A2(io_time[8]), .A3(n1494), .A4(
        io_pmp_6_addr[8]), .Y(n294) );
  AO22X1_LVT U385 ( .A1(n1485), .A2(reg_mscratch[8]), .A3(n1489), .A4(
        reg_mepc[8]), .Y(n295) );
  NOR3X0_LVT U386 ( .A1(n293), .A2(n294), .A3(n295), .Y(n296) );
  AO22X1_LVT U387 ( .A1(n1479), .A2(io_pmp_7_addr[8]), .A3(n1492), .A4(
        io_pmp_2_addr[8]), .Y(n297) );
  AO22X1_LVT U388 ( .A1(n1472), .A2(io_pmp_5_addr[8]), .A3(n1480), .A4(
        io_pmp_0_addr[8]), .Y(n298) );
  AO22X1_LVT U389 ( .A1(n1508), .A2(reg_sscratch[8]), .A3(n1510), .A4(
        reg_dscratch[8]), .Y(n299) );
  AO22X1_LVT U390 ( .A1(n1507), .A2(io_pmp_1_cfg_r), .A3(n1506), .A4(
        reg_sepc[8]), .Y(n300) );
  NOR4X0_LVT U391 ( .A1(n297), .A2(n298), .A3(n299), .A4(n300), .Y(n301) );
  NAND4X0_LVT U392 ( .A1(n284), .A2(n292), .A3(n296), .A4(n301), .Y(
        io_rw_rdata[8]) );
  INVX0_LVT U393 ( .A(io_csr_stall), .Y(n302) );
  AND3X1_LVT U394 ( .A1(io_time[0]), .A2(io_time[1]), .A3(n302), .Y(n1142) );
  AND3X1_LVT U395 ( .A1(n1514), .A2(n1512), .A3(n1526), .Y(n1507) );
  INVX0_LVT U396 ( .A(n1467), .Y(n303) );
  OA21X1_LVT U397 ( .A1(n1201), .A2(n303), .A3(n1471), .Y(n366) );
  INVX0_LVT U398 ( .A(n376), .Y(n304) );
  NAND2X0_LVT U399 ( .A1(wdata[31]), .A2(n304), .Y(n370) );
  INVX0_LVT U400 ( .A(io_rw_wdata[10]), .Y(n305) );
  OA222X1_LVT U401 ( .A1(io_rw_wdata[10]), .A2(n589), .A3(io_rw_wdata[10]), 
        .A4(io_rw_rdata[10]), .A5(n516), .A6(n305), .Y(wdata[10]) );
  INVX0_LVT U402 ( .A(io_rw_wdata[26]), .Y(n306) );
  OA222X1_LVT U403 ( .A1(io_rw_wdata[26]), .A2(n589), .A3(io_rw_wdata[26]), 
        .A4(io_rw_rdata[26]), .A5(n516), .A6(n306), .Y(wdata[26]) );
  INVX0_LVT U404 ( .A(io_rw_wdata[24]), .Y(n307) );
  OA222X1_LVT U405 ( .A1(io_rw_wdata[24]), .A2(io_rw_rdata[24]), .A3(
        io_rw_wdata[24]), .A4(n589), .A5(n516), .A6(n307), .Y(wdata[24]) );
  INVX0_LVT U406 ( .A(io_rw_wdata[22]), .Y(n308) );
  OA222X1_LVT U407 ( .A1(io_rw_wdata[22]), .A2(n589), .A3(io_rw_wdata[22]), 
        .A4(io_rw_rdata[22]), .A5(n516), .A6(n308), .Y(wdata[22]) );
  INVX0_LVT U408 ( .A(io_rw_wdata[21]), .Y(n309) );
  OA222X1_LVT U409 ( .A1(io_rw_wdata[21]), .A2(io_rw_rdata[21]), .A3(
        io_rw_wdata[21]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n309), .Y(
        wdata[21]) );
  INVX0_LVT U410 ( .A(io_rw_wdata[20]), .Y(n310) );
  OA222X1_LVT U411 ( .A1(io_rw_wdata[20]), .A2(io_rw_rdata[20]), .A3(
        io_rw_wdata[20]), .A4(n589), .A5(n516), .A6(n310), .Y(wdata[20]) );
  INVX0_LVT U412 ( .A(io_rw_wdata[18]), .Y(n311) );
  OA222X1_LVT U413 ( .A1(io_rw_wdata[18]), .A2(n589), .A3(io_rw_wdata[18]), 
        .A4(io_rw_rdata[18]), .A5(n516), .A6(n311), .Y(wdata[18]) );
  INVX0_LVT U414 ( .A(io_rw_wdata[28]), .Y(n312) );
  OA222X1_LVT U415 ( .A1(io_rw_wdata[28]), .A2(n589), .A3(io_rw_wdata[28]), 
        .A4(io_rw_rdata[28]), .A5(n516), .A6(n312), .Y(wdata[28]) );
  INVX0_LVT U416 ( .A(io_rw_wdata[30]), .Y(n313) );
  OA222X1_LVT U417 ( .A1(io_rw_wdata[30]), .A2(n589), .A3(io_rw_wdata[30]), 
        .A4(io_rw_rdata[30]), .A5(n516), .A6(n313), .Y(wdata[30]) );
  INVX0_LVT U418 ( .A(io_rw_wdata[33]), .Y(n314) );
  OA222X1_LVT U419 ( .A1(io_rw_wdata[33]), .A2(n589), .A3(io_rw_wdata[33]), 
        .A4(io_rw_rdata[33]), .A5(n516), .A6(n314), .Y(wdata[33]) );
  INVX0_LVT U420 ( .A(io_rw_wdata[36]), .Y(n315) );
  OA222X1_LVT U421 ( .A1(io_rw_wdata[36]), .A2(io_rw_rdata[36]), .A3(
        io_rw_wdata[36]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n315), .Y(
        wdata[36]) );
  INVX0_LVT U422 ( .A(io_rw_wdata[37]), .Y(n316) );
  OA222X1_LVT U423 ( .A1(io_rw_wdata[37]), .A2(n589), .A3(io_rw_wdata[37]), 
        .A4(io_rw_rdata[37]), .A5(n516), .A6(n316), .Y(wdata[37]) );
  INVX0_LVT U424 ( .A(io_rw_wdata[43]), .Y(n317) );
  OA222X1_LVT U425 ( .A1(io_rw_wdata[43]), .A2(io_rw_rdata[43]), .A3(
        io_rw_wdata[43]), .A4(n589), .A5(n516), .A6(n317), .Y(wdata[43]) );
  AO22X1_LVT U426 ( .A1(n497), .A2(n_T_52[48]), .A3(wdata[54]), .A4(n1149), 
        .Y(N1939) );
  INVX0_LVT U427 ( .A(io_rw_wdata[59]), .Y(n318) );
  OA222X1_LVT U428 ( .A1(io_rw_wdata[59]), .A2(n_T_366_59_), .A3(
        io_rw_wdata[59]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n318), .Y(n319) );
  AND3X1_LVT U429 ( .A1(n503), .A2(n319), .A3(io_status_debug), .Y(n1482) );
  INVX0_LVT U430 ( .A(io_rw_wdata[7]), .Y(n320) );
  OA222X1_LVT U431 ( .A1(io_rw_wdata[7]), .A2(n589), .A3(io_rw_wdata[7]), .A4(
        io_rw_rdata[7]), .A5(n516), .A6(n320), .Y(wdata[7]) );
  INVX0_LVT U432 ( .A(io_rw_wdata[0]), .Y(n321) );
  OA222X1_LVT U433 ( .A1(io_rw_wdata[0]), .A2(n589), .A3(io_rw_wdata[0]), .A4(
        io_rw_rdata[0]), .A5(n516), .A6(n321), .Y(wdata[0]) );
  INVX0_LVT U434 ( .A(n1181), .Y(n322) );
  AO21X1_LVT U435 ( .A1(n1190), .A2(n322), .A3(n1182), .Y(n323) );
  OR3X1_LVT U436 ( .A1(n1392), .A2(n490), .A3(io_decode_0_csr[5]), .Y(n1378)
         );
  AO22X1_LVT U437 ( .A1(n1162), .A2(io_time[21]), .A3(n1472), .A4(
        io_pmp_5_addr[21]), .Y(n324) );
  AO22X1_LVT U438 ( .A1(n1480), .A2(io_pmp_0_addr[21]), .A3(n1492), .A4(
        io_pmp_2_addr[21]), .Y(n325) );
  AO22X1_LVT U439 ( .A1(n1496), .A2(io_pmp_1_addr[21]), .A3(n1494), .A4(
        io_pmp_6_addr[21]), .Y(n326) );
  AO22X1_LVT U440 ( .A1(n1510), .A2(reg_dscratch[21]), .A3(n1479), .A4(
        io_pmp_7_addr[21]), .Y(n327) );
  NOR4X0_LVT U441 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .Y(n328) );
  AOI22X1_LVT U442 ( .A1(n1506), .A2(reg_sepc[21]), .A3(n1490), .A4(
        io_bp_0_address[21]), .Y(n329) );
  AO22X1_LVT U443 ( .A1(n1485), .A2(reg_mscratch[21]), .A3(n1493), .A4(
        reg_dpc[21]), .Y(n330) );
  AO22X1_LVT U444 ( .A1(n1491), .A2(io_pmp_4_addr[21]), .A3(n1473), .A4(
        io_pmp_3_addr[21]), .Y(n331) );
  AO22X1_LVT U445 ( .A1(n1160), .A2(n_T_444[21]), .A3(n1489), .A4(reg_mepc[21]), .Y(n332) );
  AO222X1_LVT U446 ( .A1(n1689), .A2(n_T_45[21]), .A3(n1497), .A4(
        reg_mtvec[21]), .A5(n1487), .A6(reg_stvec[21]), .Y(n333) );
  AO22X1_LVT U447 ( .A1(n1508), .A2(reg_sscratch[21]), .A3(n1157), .A4(n1925), 
        .Y(n334) );
  NOR4X0_LVT U449 ( .A1(n330), .A2(n331), .A3(n332), .A4(n336), .Y(n337) );
  NAND3X0_LVT U450 ( .A1(n328), .A2(n329), .A3(n337), .Y(io_rw_rdata[21]) );
  AND4X1_LVT U451 ( .A1(io_rw_addr[0]), .A2(io_rw_addr[2]), .A3(n1519), .A4(
        n633), .Y(n338) );
  AND2X1_LVT U452 ( .A1(n1527), .A2(n338), .Y(n1487) );
  INVX0_LVT U453 ( .A(io_rw_wdata[6]), .Y(n339) );
  OA222X1_LVT U454 ( .A1(io_rw_wdata[6]), .A2(io_rw_rdata[6]), .A3(
        io_rw_wdata[6]), .A4(n589), .A5(n516), .A6(n339), .Y(wdata[6]) );
  INVX0_LVT U455 ( .A(io_rw_wdata[4]), .Y(n340) );
  OA222X1_LVT U456 ( .A1(io_rw_wdata[4]), .A2(n589), .A3(io_rw_wdata[4]), .A4(
        io_rw_rdata[4]), .A5(n516), .A6(n340), .Y(wdata[4]) );
  INVX0_LVT U457 ( .A(io_rw_wdata[14]), .Y(n341) );
  OA222X1_LVT U458 ( .A1(io_rw_wdata[14]), .A2(n589), .A3(io_rw_wdata[14]), 
        .A4(io_rw_rdata[14]), .A5(n516), .A6(n341), .Y(wdata[14]) );
  INVX0_LVT U459 ( .A(io_rw_wdata[29]), .Y(n342) );
  OA222X1_LVT U460 ( .A1(io_rw_wdata[29]), .A2(io_rw_rdata[29]), .A3(
        io_rw_wdata[29]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n342), .Y(
        wdata[29]) );
  INVX0_LVT U461 ( .A(io_rw_wdata[27]), .Y(n343) );
  OA222X1_LVT U462 ( .A1(io_rw_wdata[27]), .A2(io_rw_rdata[27]), .A3(
        io_rw_wdata[27]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n343), .Y(
        wdata[27]) );
  INVX0_LVT U463 ( .A(io_rw_wdata[16]), .Y(n344) );
  OA222X1_LVT U464 ( .A1(io_rw_wdata[16]), .A2(io_rw_rdata[16]), .A3(
        io_rw_wdata[16]), .A4(n589), .A5(n516), .A6(n344), .Y(wdata[16]) );
  INVX0_LVT U465 ( .A(io_rw_wdata[15]), .Y(n345) );
  OA222X1_LVT U466 ( .A1(io_rw_wdata[15]), .A2(io_rw_rdata[15]), .A3(
        io_rw_wdata[15]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n345), .Y(
        wdata[15]) );
  INVX0_LVT U467 ( .A(io_rw_wdata[19]), .Y(n346) );
  OA222X1_LVT U468 ( .A1(io_rw_wdata[19]), .A2(n589), .A3(io_rw_wdata[19]), 
        .A4(io_rw_rdata[19]), .A5(n516), .A6(n346), .Y(wdata[19]) );
  INVX0_LVT U469 ( .A(io_rw_wdata[23]), .Y(n347) );
  OA222X1_LVT U470 ( .A1(io_rw_wdata[23]), .A2(io_rw_rdata[23]), .A3(
        io_rw_wdata[23]), .A4(n589), .A5(n516), .A6(n347), .Y(wdata[23]) );
  INVX0_LVT U471 ( .A(io_rw_wdata[13]), .Y(n348) );
  OA222X1_LVT U472 ( .A1(io_rw_wdata[13]), .A2(n589), .A3(io_rw_wdata[13]), 
        .A4(io_rw_rdata[13]), .A5(n516), .A6(n348), .Y(wdata[13]) );
  INVX0_LVT U473 ( .A(io_rw_wdata[31]), .Y(n349) );
  OA222X1_LVT U474 ( .A1(io_rw_wdata[31]), .A2(io_rw_rdata[31]), .A3(
        io_rw_wdata[31]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n349), .Y(
        wdata[31]) );
  INVX0_LVT U475 ( .A(io_rw_wdata[32]), .Y(n350) );
  OA222X1_LVT U476 ( .A1(io_rw_wdata[32]), .A2(io_rw_rdata[32]), .A3(
        io_rw_wdata[32]), .A4(n589), .A5(n516), .A6(n350), .Y(wdata[32]) );
  INVX0_LVT U477 ( .A(io_rw_wdata[34]), .Y(n351) );
  OA222X1_LVT U478 ( .A1(io_rw_wdata[34]), .A2(io_rw_rdata[34]), .A3(
        io_rw_wdata[34]), .A4(n589), .A5(n516), .A6(n351), .Y(wdata[34]) );
  INVX0_LVT U479 ( .A(io_rw_wdata[35]), .Y(n352) );
  OA222X1_LVT U480 ( .A1(io_rw_wdata[35]), .A2(io_rw_rdata[35]), .A3(
        io_rw_wdata[35]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n352), .Y(
        wdata[35]) );
  INVX0_LVT U481 ( .A(io_rw_wdata[61]), .Y(n353) );
  OA222X1_LVT U482 ( .A1(io_rw_wdata[61]), .A2(io_rw_rdata[61]), .A3(
        io_rw_wdata[61]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n353), .Y(
        wdata[61]) );
  INVX0_LVT U483 ( .A(io_rw_wdata[46]), .Y(n354) );
  OA222X1_LVT U484 ( .A1(io_rw_wdata[46]), .A2(io_rw_rdata[46]), .A3(
        io_rw_wdata[46]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n354), .Y(
        wdata[46]) );
  INVX0_LVT U485 ( .A(io_rw_wdata[47]), .Y(n355) );
  OA222X1_LVT U486 ( .A1(io_rw_wdata[47]), .A2(io_rw_rdata[47]), .A3(
        io_rw_wdata[47]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n355), .Y(
        wdata[47]) );
  INVX0_LVT U487 ( .A(io_rw_wdata[54]), .Y(n356) );
  OA222X1_LVT U488 ( .A1(io_rw_wdata[54]), .A2(io_rw_rdata[54]), .A3(
        io_rw_wdata[54]), .A4(io_rw_cmd[1]), .A5(n516), .A6(n356), .Y(
        wdata[54]) );
  INVX0_LVT U489 ( .A(io_rw_wdata[38]), .Y(n357) );
  OA222X1_LVT U490 ( .A1(io_rw_wdata[38]), .A2(io_rw_rdata[38]), .A3(
        io_rw_wdata[38]), .A4(n589), .A5(n516), .A6(n357), .Y(wdata[38]) );
  INVX0_LVT U491 ( .A(n1501), .Y(n358) );
  OAI22X1_LVT U492 ( .A1(n1455), .A2(n1483), .A3(n899), .A4(n358), .Y(N1272)
         );
  INVX0_LVT U493 ( .A(io_rw_wdata[8]), .Y(n359) );
  OA222X1_LVT U494 ( .A1(io_rw_wdata[8]), .A2(n589), .A3(io_rw_wdata[8]), .A4(
        io_rw_rdata[8]), .A5(n516), .A6(n359), .Y(wdata[8]) );
  INVX0_LVT U495 ( .A(io_rw_wdata[12]), .Y(n360) );
  OA222X1_LVT U496 ( .A1(io_rw_wdata[12]), .A2(n589), .A3(io_rw_wdata[12]), 
        .A4(io_rw_rdata[12]), .A5(n516), .A6(n360), .Y(wdata[12]) );
  HADDX1_LVT U497 ( .A0(io_csr_stall), .B0(n417), .SO(n361) );
  AO22X1_LVT U498 ( .A1(n1149), .A2(wdata[0]), .A3(n361), .A4(n1446), .Y(N1822) );
  IBUFFX2_LVT U500 ( .A(wdata[3]), .Y(n588) );
  AND2X4_LVT U501 ( .A1(n1139), .A2(n1456), .Y(n1159) );
  IBUFFX8_LVT U502 ( .A(n629), .Y(n1149) );
  AND2X4_LVT U503 ( .A1(n1139), .A2(n1457), .Y(n1152) );
  AND2X1_LVT U504 ( .A1(wdata[48]), .A2(wdata[49]), .Y(n369) );
  AND2X1_LVT U505 ( .A1(n590), .A2(wdata[0]), .Y(n371) );
  OR2X1_LVT U506 ( .A1(n860), .A2(n372), .Y(n373) );
  AND2X1_LVT U507 ( .A1(n375), .A2(wdata[55]), .Y(n374) );
  AND2X1_LVT U508 ( .A1(n1459), .A2(n673), .Y(n1129) );
  AND2X1_LVT U509 ( .A1(n1446), .A2(n1445), .Y(n1150) );
  IBUFFX2_LVT U510 ( .A(n957), .Y(n1128) );
  INVX1_LVT U511 ( .A(n389), .Y(n503) );
  INVX2_LVT U512 ( .A(n389), .Y(n375) );
  INVX1_LVT U513 ( .A(io_cause[0]), .Y(n954) );
  INVX1_LVT U514 ( .A(io_cause[1]), .Y(n902) );
  INVX0_LVT U515 ( .A(io_decode_0_csr[5]), .Y(n1406) );
  INVX1_LVT U516 ( .A(io_decode_0_csr[6]), .Y(n1376) );
  INVX1_LVT U517 ( .A(io_decode_0_csr[11]), .Y(n1405) );
  INVX1_LVT U518 ( .A(io_decode_0_csr[2]), .Y(n1417) );
  INVX1_LVT U519 ( .A(io_decode_0_csr[3]), .Y(n1430) );
  INVX1_LVT U520 ( .A(io_rw_wdata[9]), .Y(n1907) );
  INVX1_LVT U521 ( .A(io_rw_wdata[5]), .Y(n1904) );
  INVX0_LVT U522 ( .A(io_rw_addr[2]), .Y(n1518) );
  INVX0_LVT U523 ( .A(io_rw_addr[7]), .Y(n1528) );
  NOR2X1_LVT U524 ( .A1(io_rw_addr[4]), .A2(io_rw_addr[3]), .Y(n1529) );
  INVX1_LVT U525 ( .A(io_rw_addr[1]), .Y(n1519) );
  INVX1_LVT U526 ( .A(io_rw_wdata[1]), .Y(n697) );
  INVX0_LVT U527 ( .A(io_rw_addr[9]), .Y(n1515) );
  NOR2X1_LVT U528 ( .A1(io_rw_addr[0]), .A2(io_rw_addr[1]), .Y(n630) );
  INVX1_LVT U529 ( .A(io_rw_addr[4]), .Y(n1521) );
  INVX1_LVT U530 ( .A(n590), .Y(n378) );
  INVX1_LVT U531 ( .A(io_interrupts_debug), .Y(n1186) );
  IBUFFX2_LVT U532 ( .A(n590), .Y(n376) );
  INVX0_LVT U533 ( .A(n1468), .Y(n1346) );
  INVX1_LVT U534 ( .A(n1352), .Y(n1348) );
  OR2X1_LVT U535 ( .A1(n1442), .A2(n1441), .Y(n1462) );
  INVX1_LVT U536 ( .A(n925), .Y(n1461) );
  OR2X1_LVT U537 ( .A1(n1199), .A2(n1441), .Y(n1352) );
  INVX0_LVT U538 ( .A(n908), .Y(n911) );
  INVX0_LVT U539 ( .A(n1416), .Y(n1436) );
  INVX0_LVT U540 ( .A(n1374), .Y(n1373) );
  NOR2X1_LVT U541 ( .A1(n1481), .A2(n1690), .Y(n968) );
  NOR2X1_LVT U542 ( .A1(n1458), .A2(n956), .Y(n712) );
  INVX0_LVT U543 ( .A(n1427), .Y(n1418) );
  NOR2X1_LVT U544 ( .A1(n1653), .A2(n1657), .Y(n650) );
  NOR2X1_LVT U545 ( .A1(n1140), .A2(n1139), .Y(N1821) );
  NOR2X1_LVT U546 ( .A1(n1590), .A2(n1589), .Y(n1094) );
  NOR2X1_LVT U547 ( .A1(n1585), .A2(n1586), .Y(n1107) );
  INVX0_LVT U548 ( .A(n1432), .Y(n1433) );
  NOR2X1_LVT U549 ( .A1(n1621), .A2(n1624), .Y(n1052) );
  OR2X1_LVT U550 ( .A1(n708), .A2(n1467), .Y(n1257) );
  INVX0_LVT U551 ( .A(n961), .Y(n1458) );
  INVX0_LVT U552 ( .A(n1495), .Y(n484) );
  INVX0_LVT U553 ( .A(n1381), .Y(n1367) );
  OA22X1_LVT U554 ( .A1(n490), .A2(n1419), .A3(io_decode_0_csr[7]), .A4(n1398), 
        .Y(n1404) );
  INVX0_LVT U555 ( .A(n1419), .Y(n1420) );
  INVX0_LVT U556 ( .A(n1375), .Y(n1377) );
  AND2X1_LVT U557 ( .A1(n629), .A2(n590), .Y(n1446) );
  NOR2X1_LVT U558 ( .A1(n1584), .A2(n1583), .Y(n1109) );
  INVX0_LVT U559 ( .A(n702), .Y(n949) );
  INVX0_LVT U560 ( .A(n1445), .Y(n1447) );
  NOR2X1_LVT U561 ( .A1(n1180), .A2(n1189), .Y(n1185) );
  INVX0_LVT U562 ( .A(n1455), .Y(n923) );
  INVX0_LVT U563 ( .A(n1139), .Y(n1442) );
  INVX0_LVT U564 ( .A(n1171), .Y(n1170) );
  NAND3X0_LVT U565 ( .A1(n503), .A2(n672), .A3(n671), .Y(n957) );
  INVX0_LVT U566 ( .A(n1209), .Y(n888) );
  INVX0_LVT U567 ( .A(n1226), .Y(n895) );
  INVX1_LVT U568 ( .A(n891), .Y(n1202) );
  INVX1_LVT U569 ( .A(n1041), .Y(n1157) );
  OR2X1_LVT U570 ( .A1(n699), .A2(io_exception), .Y(n1139) );
  INVX0_LVT U571 ( .A(n1378), .Y(n1380) );
  INVX0_LVT U572 ( .A(n1384), .Y(n1385) );
  INVX0_LVT U573 ( .A(n1155), .Y(n1156) );
  AND3X1_LVT U574 ( .A1(io_rw_addr[1]), .A2(n1520), .A3(n1531), .Y(n1689) );
  INVX0_LVT U575 ( .A(n1210), .Y(n1211) );
  INVX0_LVT U576 ( .A(n1154), .Y(n1026) );
  INVX0_LVT U577 ( .A(n1903), .Y(n1199) );
  MUX21X1_LVT U578 ( .A1(n700), .A2(io_cause[1]), .S0(n1697), .Y(n1209) );
  MUX21X1_LVT U579 ( .A1(n1520), .A2(io_cause[3]), .S0(n1697), .Y(n1226) );
  NOR2X1_LVT U580 ( .A1(io_rw_addr[9]), .A2(n1903), .Y(n1355) );
  MUX21X1_LVT U581 ( .A1(n953), .A2(n954), .S0(n1697), .Y(n891) );
  INVX0_LVT U582 ( .A(n1697), .Y(n699) );
  INVX0_LVT U583 ( .A(n1368), .Y(n1369) );
  NOR2X1_LVT U584 ( .A1(n1520), .A2(n1697), .Y(n1210) );
  INVX0_LVT U585 ( .A(n866), .Y(n743) );
  INVX0_LVT U586 ( .A(n1179), .Y(n1169) );
  AND2X1_LVT U587 ( .A1(n620), .A2(n1505), .Y(n1474) );
  INVX0_LVT U588 ( .A(n1144), .Y(n1141) );
  AND2X1_LVT U589 ( .A1(n620), .A2(n676), .Y(n1153) );
  NOR2X1_LVT U590 ( .A1(n605), .A2(n601), .Y(n488) );
  INVX0_LVT U591 ( .A(n1192), .Y(n1184) );
  AND2X1_LVT U592 ( .A1(n858), .A2(n857), .Y(n1469) );
  NOR2X1_LVT U593 ( .A1(n427), .A2(io_cause[3]), .Y(n901) );
  NAND2X0_LVT U594 ( .A1(n504), .A2(n590), .Y(n389) );
  INVX0_LVT U595 ( .A(n1134), .Y(n941) );
  OR2X1_LVT U596 ( .A1(io_interrupts_seip), .A2(n_T_3694_9_), .Y(n1136) );
  INVX0_LVT U597 ( .A(n1178), .Y(n1177) );
  NOR2X1_LVT U598 ( .A1(io_decode_0_csr[1]), .A2(io_decode_0_csr[0]), .Y(n1390) );
  INVX1_LVT U599 ( .A(n489), .Y(n490) );
  NOR2X1_LVT U600 ( .A1(io_decode_0_csr[9]), .A2(io_decode_0_csr[6]), .Y(n1379) );
  INVX0_LVT U601 ( .A(n1176), .Y(n1187) );
  INVX0_LVT U602 ( .A(n1172), .Y(n1173) );
  NOR4X0_LVT U603 ( .A1(io_rw_addr[4]), .A2(io_rw_addr[3]), .A3(n1525), .A4(
        n1524), .Y(n1526) );
  AND2X1_LVT U604 ( .A1(n630), .A2(n1518), .Y(n1512) );
  OR2X1_LVT U605 ( .A1(io_decode_0_csr[4]), .A2(io_decode_0_csr[3]), .Y(n1392)
         );
  INVX1_LVT U606 ( .A(io_decode_0_csr[10]), .Y(n489) );
  INVX0_LVT U607 ( .A(n605), .Y(n633) );
  INVX0_LVT U608 ( .A(io_decode_0_csr[8]), .Y(n1371) );
  INVX0_LVT U609 ( .A(n597), .Y(n598) );
  NOR2X1_LVT U610 ( .A1(io_status_prv[0]), .A2(io_rw_addr[0]), .Y(n953) );
  OR2X1_LVT U611 ( .A1(io_rw_addr[6]), .A2(io_rw_addr[9]), .Y(n605) );
  NBUFFX2_LVT U612 ( .A(net35092), .Y(n531) );
  IBUFFX4_LVT U613 ( .A(reset), .Y(n590) );
  MUX21X1_LVT U614 ( .A1(n588), .A2(n880), .S0(n879), .Y(n1909) );
  MUX21X1_LVT U615 ( .A1(io_pc[3]), .A2(wdata[3]), .S0(n515), .Y(net35295) );
  MUX21X1_LVT U616 ( .A1(io_pc[9]), .A2(wdata[9]), .S0(n514), .Y(net35055) );
  OAI21X1_LVT U617 ( .A1(n_T_45[2]), .A2(n956), .A3(n961), .Y(n958) );
  NBUFFX2_LVT U618 ( .A(clock), .Y(n594) );
  NBUFFX2_LVT U619 ( .A(net34722), .Y(n586) );
  NBUFFX2_LVT U620 ( .A(net34722), .Y(n585) );
  NBUFFX2_LVT U621 ( .A(net34722), .Y(n584) );
  NBUFFX2_LVT U622 ( .A(net34950), .Y(n556) );
  NBUFFX2_LVT U623 ( .A(net34925), .Y(n567) );
  NBUFFX2_LVT U624 ( .A(net34955), .Y(n553) );
  NBUFFX2_LVT U625 ( .A(net35309), .Y(n527) );
  NBUFFX2_LVT U626 ( .A(net34950), .Y(n554) );
  NBUFFX2_LVT U627 ( .A(net34950), .Y(n555) );
  NBUFFX2_LVT U628 ( .A(net34890), .Y(n579) );
  NBUFFX2_LVT U629 ( .A(net34920), .Y(n569) );
  NBUFFX2_LVT U630 ( .A(net34920), .Y(n570) );
  NBUFFX2_LVT U631 ( .A(net34920), .Y(n568) );
  NBUFFX2_LVT U632 ( .A(net34890), .Y(n576) );
  NBUFFX2_LVT U633 ( .A(net34890), .Y(n577) );
  NBUFFX2_LVT U634 ( .A(net34890), .Y(n575) );
  NBUFFX2_LVT U635 ( .A(net34890), .Y(n578) );
  NBUFFX2_LVT U636 ( .A(net35304), .Y(n529) );
  NBUFFX2_LVT U637 ( .A(net34880), .Y(n581) );
  NBUFFX2_LVT U638 ( .A(net35304), .Y(n530) );
  NBUFFX2_LVT U639 ( .A(net35082), .Y(n546) );
  NBUFFX2_LVT U640 ( .A(net35082), .Y(n545) );
  NBUFFX2_LVT U641 ( .A(net34880), .Y(n582) );
  NBUFFX2_LVT U642 ( .A(net35082), .Y(n547) );
  NBUFFX2_LVT U643 ( .A(net35304), .Y(n528) );
  NBUFFX2_LVT U644 ( .A(net34880), .Y(n583) );
  NBUFFX2_LVT U645 ( .A(net34955), .Y(n551) );
  NBUFFX2_LVT U646 ( .A(net34925), .Y(n565) );
  NBUFFX2_LVT U647 ( .A(net35309), .Y(n525) );
  NBUFFX2_LVT U648 ( .A(net34925), .Y(n563) );
  NBUFFX2_LVT U649 ( .A(net34955), .Y(n549) );
  NBUFFX2_LVT U650 ( .A(net35309), .Y(n522) );
  NBUFFX2_LVT U651 ( .A(net35309), .Y(n523) );
  NBUFFX2_LVT U652 ( .A(net35309), .Y(n524) );
  NBUFFX2_LVT U653 ( .A(net35309), .Y(n526) );
  NBUFFX2_LVT U654 ( .A(net34925), .Y(n566) );
  NBUFFX2_LVT U655 ( .A(net34955), .Y(n548) );
  NBUFFX2_LVT U656 ( .A(net34955), .Y(n552) );
  NBUFFX2_LVT U657 ( .A(net34955), .Y(n550) );
  NBUFFX2_LVT U658 ( .A(net34925), .Y(n562) );
  NBUFFX2_LVT U659 ( .A(net34925), .Y(n564) );
  NBUFFX2_LVT U660 ( .A(net34930), .Y(n560) );
  NBUFFX2_LVT U661 ( .A(net34930), .Y(n561) );
  NBUFFX2_LVT U662 ( .A(clock), .Y(n593) );
  NBUFFX2_LVT U663 ( .A(net34895), .Y(n573) );
  NBUFFX2_LVT U664 ( .A(net34895), .Y(n574) );
  NBUFFX2_LVT U665 ( .A(net34930), .Y(n559) );
  NBUFFX2_LVT U666 ( .A(net34895), .Y(n572) );
  NBUFFX2_LVT U667 ( .A(n1128), .Y(n491) );
  NBUFFX2_LVT U668 ( .A(net35092), .Y(n538) );
  NBUFFX2_LVT U669 ( .A(net35092), .Y(n540) );
  NBUFFX2_LVT U670 ( .A(net35092), .Y(n539) );
  NBUFFX2_LVT U671 ( .A(net35092), .Y(n537) );
  NBUFFX2_LVT U672 ( .A(net35092), .Y(n536) );
  NBUFFX2_LVT U673 ( .A(net35092), .Y(n535) );
  NBUFFX2_LVT U674 ( .A(net35092), .Y(n534) );
  NBUFFX2_LVT U675 ( .A(net35092), .Y(n533) );
  NBUFFX2_LVT U676 ( .A(net35092), .Y(n532) );
  NAND4X0_LVT U677 ( .A1(n940), .A2(n590), .A3(n939), .A4(n938), .Y(n2160) );
  NAND3X0_LVT U678 ( .A1(n1462), .A2(n1443), .A3(n501), .Y(n1917) );
  NBUFFX2_LVT U679 ( .A(n531), .Y(n544) );
  NBUFFX2_LVT U680 ( .A(n531), .Y(n542) );
  NBUFFX2_LVT U681 ( .A(n531), .Y(n541) );
  NBUFFX2_LVT U682 ( .A(n531), .Y(n543) );
  NBUFFX2_LVT U683 ( .A(clock), .Y(n592) );
  NAND4X0_LVT U684 ( .A1(n915), .A2(n590), .A3(n387), .A4(n501), .Y(n921) );
  MUX21X1_LVT U685 ( .A1(n927), .A2(n926), .S0(n387), .Y(n928) );
  NAND2X0_LVT U686 ( .A1(n906), .A2(n381), .Y(n1255) );
  MUX21X1_LVT U687 ( .A1(n905), .A2(n904), .S0(n1201), .Y(n906) );
  MUX21X1_LVT U688 ( .A1(n1411), .A2(n1410), .S0(io_decode_0_csr[0]), .Y(n1415) );
  OR2X1_LVT U689 ( .A1(n1370), .A2(n1369), .Y(n1419) );
  INVX1_LVT U690 ( .A(io_decode_0_csr[7]), .Y(n1386) );
  INVX1_LVT U691 ( .A(io_decode_0_csr[1]), .Y(n1407) );
  MUX21X1_LVT U692 ( .A1(io_pc[11]), .A2(wdata[11]), .S0(n513), .Y(net34847)
         );
  MUX21X1_LVT U693 ( .A1(io_pc[11]), .A2(wdata[11]), .S0(n515), .Y(net35271)
         );
  MUX21X1_LVT U694 ( .A1(io_pc[7]), .A2(wdata[7]), .S0(n513), .Y(net34859) );
  MUX21X1_LVT U695 ( .A1(io_pc[7]), .A2(wdata[7]), .S0(n515), .Y(net35283) );
  MUX21X1_LVT U696 ( .A1(io_pc[7]), .A2(wdata[7]), .S0(n514), .Y(net35061) );
  MUX21X1_LVT U697 ( .A1(io_pmp_1_addr[3]), .A2(wdata[3]), .S0(n506), .Y(
        n_GEN_265[3]) );
  MUX21X1_LVT U698 ( .A1(io_pmp_7_addr[9]), .A2(wdata[9]), .S0(n512), .Y(
        n_GEN_307[9]) );
  MUX21X1_LVT U699 ( .A1(io_pmp_2_addr[9]), .A2(wdata[9]), .S0(n507), .Y(
        n_GEN_272[9]) );
  MUX21X1_LVT U700 ( .A1(io_pmp_0_addr[9]), .A2(wdata[9]), .S0(n505), .Y(
        n_GEN_258[9]) );
  INVX1_LVT U701 ( .A(n436), .Y(n508) );
  INVX1_LVT U702 ( .A(n433), .Y(n509) );
  INVX1_LVT U703 ( .A(n432), .Y(n507) );
  INVX1_LVT U704 ( .A(n434), .Y(n510) );
  INVX1_LVT U705 ( .A(n431), .Y(n506) );
  INVX1_LVT U706 ( .A(n435), .Y(n511) );
  INVX1_LVT U707 ( .A(n386), .Y(n512) );
  INVX1_LVT U708 ( .A(n430), .Y(n505) );
  INVX1_LVT U709 ( .A(n448), .Y(n513) );
  NAND2X0_LVT U710 ( .A1(n1496), .A2(n745), .Y(n431) );
  INVX1_LVT U711 ( .A(n450), .Y(n515) );
  NAND2X0_LVT U712 ( .A1(n1479), .A2(n442), .Y(n386) );
  INVX1_LVT U713 ( .A(n449), .Y(n514) );
  INVX1_LVT U714 ( .A(n1483), .Y(wdata[2]) );
  MUX21X1_LVT U715 ( .A1(n668), .A2(n444), .S0(io_rw_wdata[2]), .Y(n1483) );
  AO22X1_LVT U716 ( .A1(io_rw_wdata[1]), .A2(n516), .A3(io_rw_rdata[1]), .A4(
        n1476), .Y(wdata[1]) );
  INVX1_LVT U717 ( .A(n1456), .Y(n1158) );
  INVX1_LVT U718 ( .A(n1457), .Y(n1151) );
  INVX1_LVT U719 ( .A(n444), .Y(n516) );
  NBUFFX2_LVT U720 ( .A(io_rw_cmd[1]), .Y(n589) );
  INVX1_LVT U721 ( .A(n387), .Y(n504) );
  NAND2X0_LVT U722 ( .A1(io_rw_cmd[2]), .A2(n597), .Y(n387) );
  INVX1_LVT U723 ( .A(n501), .Y(n500) );
  INVX1_LVT U724 ( .A(n1355), .Y(n501) );
  AND2X1_LVT U725 ( .A1(n1134), .A2(n942), .Y(n1356) );
  INVX1_LVT U726 ( .A(n451), .Y(n502) );
  OR2X1_LVT U727 ( .A1(n882), .A2(n1903), .Y(n451) );
  INVX1_LVT U728 ( .A(n1220), .Y(n899) );
  OR2X1_LVT U729 ( .A1(n1918), .A2(io_status_wfi), .Y(io_csr_stall) );
  NAND2X0_LVT U730 ( .A1(n1134), .A2(n600), .Y(n1697) );
  AND2X1_LVT U731 ( .A1(io_rw_cmd[2]), .A2(n598), .Y(n1134) );
  INVX1_LVT U732 ( .A(n1690), .Y(n481) );
  OR2X1_LVT U733 ( .A1(n749), .A2(n1650), .Y(n1690) );
  AND2X1_LVT U734 ( .A1(n640), .A2(n716), .Y(n1481) );
  AND2X1_LVT U735 ( .A1(n630), .A2(n1532), .Y(n1495) );
  AND2X1_LVT U736 ( .A1(n610), .A2(n1532), .Y(n1493) );
  AND2X1_LVT U737 ( .A1(n620), .A2(n1512), .Y(n1485) );
  AND2X1_LVT U738 ( .A1(n616), .A2(n662), .Y(n1494) );
  AND2X1_LVT U739 ( .A1(n616), .A2(n857), .Y(n1492) );
  AND2X1_LVT U740 ( .A1(n616), .A2(n676), .Y(n1473) );
  AND2X1_LVT U741 ( .A1(n616), .A2(n1512), .Y(n1480) );
  AND2X1_LVT U742 ( .A1(n630), .A2(n1531), .Y(n1162) );
  AND2X1_LVT U743 ( .A1(n1509), .A2(n676), .Y(n1160) );
  AND2X1_LVT U744 ( .A1(n858), .A2(n621), .Y(n1497) );
  AND2X1_LVT U745 ( .A1(n1509), .A2(n1512), .Y(n1508) );
  AND2X1_LVT U746 ( .A1(n620), .A2(n716), .Y(n1489) );
  AND2X1_LVT U747 ( .A1(n1509), .A2(n716), .Y(n1506) );
  AND2X1_LVT U748 ( .A1(n640), .A2(n857), .Y(n1490) );
  AND2X1_LVT U749 ( .A1(n616), .A2(n621), .Y(n1472) );
  NOR2X0_LVT U750 ( .A1(n605), .A2(n601), .Y(n1488) );
  AND2X1_LVT U751 ( .A1(n671), .A2(n1532), .Y(n1510) );
  AND2X1_LVT U752 ( .A1(n616), .A2(n716), .Y(n1496) );
  AND2X1_LVT U753 ( .A1(n616), .A2(n1505), .Y(n1491) );
  AND2X1_LVT U754 ( .A1(n1523), .A2(n1514), .Y(n616) );
  INVX1_LVT U755 ( .A(io_rw_addr[10]), .Y(n1514) );
  INVX1_LVT U756 ( .A(io_rw_addr[11]), .Y(n1513) );
  AND2X1_LVT U757 ( .A1(n1507), .A2(n504), .Y(n1463) );
  AND2X1_LVT U758 ( .A1(n744), .A2(n440), .Y(n745) );
  NBUFFX2_LVT U759 ( .A(n1150), .Y(n498) );
  NBUFFX2_LVT U760 ( .A(n1150), .Y(n497) );
  NBUFFX2_LVT U761 ( .A(n1150), .Y(n496) );
  AND2X1_LVT U762 ( .A1(n1147), .A2(io_time[5]), .Y(n1445) );
  NBUFFX2_LVT U763 ( .A(io_ungated_clock), .Y(n591) );
  NAND2X0_LVT U764 ( .A1(n504), .A2(n1493), .Y(n450) );
  NBUFFX2_LVT U765 ( .A(n1129), .Y(n495) );
  NBUFFX2_LVT U766 ( .A(n1129), .Y(n494) );
  NBUFFX2_LVT U767 ( .A(n1129), .Y(n493) );
  AND2X1_LVT U768 ( .A1(n961), .A2(n_T_45[5]), .Y(n673) );
  NAND2X0_LVT U769 ( .A1(n1489), .A2(n504), .Y(n449) );
  NAND2X0_LVT U770 ( .A1(n1506), .A2(n504), .Y(n448) );
  NAND2X0_LVT U771 ( .A1(n504), .A2(n1160), .Y(n1456) );
  NAND2X0_LVT U772 ( .A1(n504), .A2(n1153), .Y(n1457) );
  NAND2X0_LVT U773 ( .A1(n1903), .A2(n1697), .Y(io_eret) );
  AND3X1_LVT U774 ( .A1(io_rw_addr[10]), .A2(n1523), .A3(n1518), .Y(n1532) );
  NAND3X0_LVT U775 ( .A1(n1557), .A2(n1529), .A3(n596), .Y(n1674) );
  INVX1_LVT U776 ( .A(io_rw_addr[0]), .Y(n1520) );
  AND4X1_LVT U777 ( .A1(n1514), .A2(n1528), .A3(n1513), .A4(n1522), .Y(n1527)
         );
  AND2X1_LVT U778 ( .A1(n610), .A2(n1518), .Y(n716) );
  INVX1_LVT U779 ( .A(io_rw_addr[8]), .Y(n600) );
  NOR4X1_LVT U780 ( .A1(wdata[62]), .A2(wdata[61]), .A3(wdata[60]), .A4(n1673), 
        .Y(N1426) );
  XOR2X1_LVT U781 ( .A1(n1147), .A2(io_time[5]), .Y(n1148) );
  NBUFFX2_LVT U782 ( .A(net35324), .Y(n521) );
  NBUFFX2_LVT U783 ( .A(net35324), .Y(n518) );
  NBUFFX2_LVT U784 ( .A(net35324), .Y(n519) );
  NBUFFX2_LVT U785 ( .A(net35324), .Y(n517) );
  NBUFFX2_LVT U786 ( .A(net35324), .Y(n520) );
  AND2X1_LVT U787 ( .A1(n1460), .A2(n1499), .Y(n1498) );
  NBUFFX2_LVT U788 ( .A(net34722), .Y(n587) );
  NBUFFX2_LVT U789 ( .A(net34935), .Y(n557) );
  NBUFFX2_LVT U790 ( .A(net34885), .Y(n580) );
  NBUFFX2_LVT U791 ( .A(net34935), .Y(n558) );
  NBUFFX2_LVT U792 ( .A(net34920), .Y(n571) );
  NAND2X0_LVT U793 ( .A1(n1134), .A2(n655), .Y(n1903) );
  NOR4X1_LVT U794 ( .A1(n1567), .A2(n1566), .A3(n1565), .A4(n1564), .Y(n1570)
         );
  NOR4X1_LVT U795 ( .A1(n1611), .A2(n1610), .A3(n1609), .A4(n1608), .Y(n1613)
         );
  NOR4X1_LVT U796 ( .A1(n1537), .A2(n1536), .A3(n1535), .A4(n1534), .Y(n1544)
         );
  NOR4X1_LVT U797 ( .A1(n1551), .A2(n1550), .A3(n1549), .A4(n1548), .Y(n1555)
         );
  NOR4X1_LVT U798 ( .A1(n1574), .A2(n1573), .A3(n1572), .A4(n1571), .Y(n1581)
         );
  NOR4X1_LVT U799 ( .A1(n1578), .A2(n1577), .A3(n1576), .A4(n1575), .Y(n1580)
         );
  NOR4X1_LVT U800 ( .A1(n1670), .A2(n1669), .A3(n1668), .A4(n1667), .Y(n1671)
         );
  AND2X1_LVT U801 ( .A1(n1504), .A2(io_rw_addr[9]), .Y(n1502) );
  NOR4X1_LVT U802 ( .A1(n1601), .A2(n1600), .A3(n1599), .A4(n1598), .Y(n1605)
         );
  AOI22X1_LVT U803 ( .A1(n1478), .A2(reg_stvec[5]), .A3(n1162), .A4(io_time[5]), .Y(n379) );
  AND3X1_LVT U804 ( .A1(n468), .A2(n385), .A3(n487), .Y(n380) );
  AOI22X1_LVT U805 ( .A1(n1162), .A2(io_time[2]), .A3(n1689), .A4(n_T_45[2]), 
        .Y(n382) );
  AOI22X1_LVT U806 ( .A1(n1689), .A2(n_T_45[5]), .A3(n1477), .A4(io_fcsr_rm[0]), .Y(n384) );
  AOI22X1_LVT U807 ( .A1(n1452), .A2(n1923), .A3(reg_mepc[5]), .A4(n1489), .Y(
        n385) );
  AOI22X1_LVT U808 ( .A1(n1153), .A2(n_T_383[5]), .A3(reg_mtvec[5]), .A4(n1470), .Y(n388) );
  NBUFFX2_LVT U809 ( .A(n1128), .Y(n492) );
  NBUFFX2_LVT U810 ( .A(n1348), .Y(n499) );
  AND2X1_LVT U811 ( .A1(io_rw_cmd[0]), .A2(n589), .Y(n444) );
  AND2X1_LVT U812 ( .A1(n1512), .A2(n1514), .Y(n445) );
  AOI22X1_LVT U813 ( .A1(n1508), .A2(reg_sscratch[27]), .A3(n1506), .A4(
        reg_sepc[27]), .Y(n466) );
  AOI22X1_LVT U814 ( .A1(n1689), .A2(n_T_45[61]), .A3(n1510), .A4(
        reg_dscratch[61]), .Y(n467) );
  AOI22X1_LVT U815 ( .A1(n1160), .A2(n_T_444[5]), .A3(n1496), .A4(
        io_pmp_1_addr[5]), .Y(n468) );
  AOI22X1_LVT U816 ( .A1(n1502), .A2(reg_mie[5]), .A3(n1508), .A4(
        reg_sscratch[5]), .Y(n469) );
  AOI22X1_LVT U817 ( .A1(n1496), .A2(io_pmp_1_addr[2]), .A3(n1466), .A4(
        io_fcsr_rm[2]), .Y(n471) );
  AOI21X1_LVT U818 ( .A1(n1507), .A2(io_pmp_6_cfg_l), .A3(n755), .Y(n473) );
  AOI21X1_LVT U819 ( .A1(n1507), .A2(io_pmp_7_cfg_x), .A3(n969), .Y(n474) );
  AOI21X1_LVT U820 ( .A1(n1507), .A2(io_pmp_7_cfg_w), .A3(n971), .Y(n475) );
  AOI22X1_LVT U821 ( .A1(n1510), .A2(reg_dscratch[5]), .A3(n1485), .A4(
        reg_mscratch[5]), .Y(n476) );
  AOI21X1_LVT U822 ( .A1(n1493), .A2(reg_dpc[19]), .A3(n1591), .Y(n478) );
  NAND2X0_LVT U823 ( .A1(n1689), .A2(n_T_45[46]), .Y(n479) );
  NAND2X0_LVT U824 ( .A1(n1487), .A2(reg_stvec[30]), .Y(n480) );
  NAND3X0_LVT U825 ( .A1(n1241), .A2(n1240), .A3(n1242), .Y(io_evec[7]) );
  NAND3X0_LVT U826 ( .A1(n1234), .A2(n1233), .A3(n1235), .Y(io_evec[6]) );
  AND3X1_LVT U827 ( .A1(n1012), .A2(n1011), .A3(n1013), .Y(n1014) );
  AND3X1_LVT U828 ( .A1(n1004), .A2(n1003), .A3(n1005), .Y(n1006) );
  NAND3X0_LVT U829 ( .A1(n1000), .A2(n999), .A3(n1001), .Y(n1002) );
  AND3X1_LVT U830 ( .A1(n994), .A2(n993), .A3(n995), .Y(n996) );
  AND3X1_LVT U831 ( .A1(n990), .A2(n989), .A3(n991), .Y(n992) );
  AND3X1_LVT U832 ( .A1(n986), .A2(n985), .A3(n987), .Y(n988) );
  NAND3X0_LVT U833 ( .A1(n982), .A2(n981), .A3(n983), .Y(n984) );
  NAND3X0_LVT U834 ( .A1(n978), .A2(n977), .A3(n979), .Y(n980) );
  AND3X1_LVT U835 ( .A1(n974), .A2(n973), .A3(n975), .Y(n976) );
  NAND3X0_LVT U836 ( .A1(n963), .A2(n962), .A3(n964), .Y(n965) );
  NAND3X0_LVT U837 ( .A1(n824), .A2(n823), .A3(n825), .Y(n826) );
  AND3X1_LVT U838 ( .A1(n819), .A2(n818), .A3(n820), .Y(n821) );
  AND3X1_LVT U839 ( .A1(n815), .A2(n814), .A3(n816), .Y(n817) );
  AND3X1_LVT U840 ( .A1(n811), .A2(n810), .A3(n812), .Y(n813) );
  AND3X1_LVT U841 ( .A1(n807), .A2(n806), .A3(n808), .Y(n809) );
  NAND3X0_LVT U842 ( .A1(n776), .A2(n775), .A3(n777), .Y(n778) );
  NAND3X0_LVT U843 ( .A1(n768), .A2(n767), .A3(n769), .Y(n772) );
  NAND3X0_LVT U844 ( .A1(n752), .A2(n751), .A3(n753), .Y(n754) );
  AND3X1_LVT U845 ( .A1(n1220), .A2(n954), .A3(n1209), .Y(n707) );
  AND2X1_LVT U846 ( .A1(wdata[4]), .A2(n923), .Y(N1274) );
  AND2X1_LVT U847 ( .A1(n1508), .A2(reg_sscratch[7]), .Y(n832) );
  AND2X1_LVT U848 ( .A1(n1474), .A2(n1136), .Y(n736) );
  AND2X1_LVT U849 ( .A1(n1508), .A2(reg_sscratch[11]), .Y(n623) );
  NAND2X0_LVT U850 ( .A1(n1162), .A2(io_time[16]), .Y(n1124) );
  AND2X1_LVT U851 ( .A1(n1160), .A2(n_T_444[17]), .Y(n1577) );
  AND2X1_LVT U852 ( .A1(n1160), .A2(n_T_444[18]), .Y(n1105) );
  AND2X1_LVT U853 ( .A1(n1162), .A2(io_time[19]), .Y(n1092) );
  NAND2X0_LVT U854 ( .A1(n1508), .A2(reg_sscratch[20]), .Y(n1073) );
  AND2X1_LVT U855 ( .A1(n1489), .A2(reg_mepc[23]), .Y(n788) );
  NAND2X0_LVT U856 ( .A1(n1160), .A2(n_T_444[24]), .Y(n1060) );
  AND2X1_LVT U857 ( .A1(n1162), .A2(io_time[27]), .Y(n797) );
  AND2X1_LVT U858 ( .A1(n1160), .A2(n_T_444[29]), .Y(n1045) );
  AND2X1_LVT U859 ( .A1(n1510), .A2(reg_dscratch[32]), .Y(n1629) );
  AND2X1_LVT U860 ( .A1(n1493), .A2(reg_dpc[34]), .Y(n1636) );
  NAND2X0_LVT U861 ( .A1(n1506), .A2(reg_sepc[36]), .Y(n804) );
  AND2X1_LVT U862 ( .A1(n1485), .A2(reg_mscratch[37]), .Y(n1645) );
  NAND2X0_LVT U863 ( .A1(n1485), .A2(reg_mscratch[39]), .Y(n752) );
  NAND2X0_LVT U864 ( .A1(n1485), .A2(reg_mscratch[40]), .Y(n1013) );
  AND2X1_LVT U865 ( .A1(n1485), .A2(reg_mscratch[41]), .Y(n1008) );
  NAND2X0_LVT U866 ( .A1(n1508), .A2(reg_sscratch[42]), .Y(n1005) );
  NAND2X0_LVT U867 ( .A1(n1508), .A2(reg_sscratch[43]), .Y(n820) );
  NAND2X0_LVT U868 ( .A1(n1485), .A2(reg_mscratch[44]), .Y(n824) );
  NAND2X0_LVT U869 ( .A1(n1485), .A2(reg_mscratch[45]), .Y(n1000) );
  NAND2X0_LVT U870 ( .A1(n1485), .A2(reg_mscratch[47]), .Y(n808) );
  NAND2X0_LVT U871 ( .A1(n1508), .A2(reg_sscratch[48]), .Y(n995) );
  NAND2X0_LVT U872 ( .A1(n1485), .A2(reg_mscratch[49]), .Y(n991) );
  NAND2X0_LVT U873 ( .A1(n1508), .A2(reg_sscratch[50]), .Y(n987) );
  NAND2X0_LVT U874 ( .A1(n1508), .A2(reg_sscratch[51]), .Y(n812) );
  NAND2X0_LVT U875 ( .A1(n1485), .A2(reg_mscratch[52]), .Y(n816) );
  NAND2X0_LVT U876 ( .A1(n1485), .A2(reg_mscratch[53]), .Y(n982) );
  NAND2X0_LVT U877 ( .A1(n1485), .A2(reg_mscratch[54]), .Y(n978) );
  NAND2X0_LVT U878 ( .A1(n1485), .A2(reg_mscratch[55]), .Y(n756) );
  NAND2X0_LVT U879 ( .A1(n1485), .A2(reg_mscratch[56]), .Y(n975) );
  NAND2X0_LVT U880 ( .A1(n1162), .A2(n1942), .Y(n972) );
  NAND2X0_LVT U881 ( .A1(n1162), .A2(n1941), .Y(n970) );
  AND2X1_LVT U882 ( .A1(n1485), .A2(reg_mscratch[59]), .Y(n771) );
  NAND2X0_LVT U883 ( .A1(n1485), .A2(reg_mscratch[60]), .Y(n776) );
  NAND2X0_LVT U884 ( .A1(n1485), .A2(reg_mscratch[61]), .Y(n966) );
  NAND2X0_LVT U885 ( .A1(n1485), .A2(reg_mscratch[62]), .Y(n963) );
  AND2X1_LVT U886 ( .A1(n1477), .A2(io_fcsr_rm[2]), .Y(n827) );
  NAND2X0_LVT U887 ( .A1(n1153), .A2(n_T_383[9]), .Y(n733) );
  AND2X1_LVT U888 ( .A1(n1153), .A2(n_T_383[11]), .Y(n619) );
  NAND2X0_LVT U889 ( .A1(n1160), .A2(n_T_444[16]), .Y(n1123) );
  AND2X1_LVT U890 ( .A1(n1493), .A2(reg_dpc[17]), .Y(n1578) );
  AND2X1_LVT U891 ( .A1(n1497), .A2(reg_mtvec[18]), .Y(n1106) );
  AND2X1_LVT U892 ( .A1(n1485), .A2(reg_mscratch[19]), .Y(n1081) );
  NAND2X0_LVT U893 ( .A1(n1153), .A2(n_T_383[20]), .Y(n1072) );
  AND2X1_LVT U894 ( .A1(n1452), .A2(n1919), .Y(n784) );
  NAND2X0_LVT U895 ( .A1(n1497), .A2(reg_mtvec[24]), .Y(n1061) );
  AND2X1_LVT U896 ( .A1(n1160), .A2(n_T_444[27]), .Y(n794) );
  AND2X1_LVT U897 ( .A1(n1489), .A2(reg_mepc[29]), .Y(n1049) );
  NAND2X0_LVT U898 ( .A1(n1485), .A2(reg_mscratch[30]), .Y(n1040) );
  AND2X1_LVT U899 ( .A1(n1489), .A2(reg_mepc[32]), .Y(n1631) );
  AND2X1_LVT U900 ( .A1(n1489), .A2(reg_mepc[34]), .Y(n1634) );
  NAND2X0_LVT U901 ( .A1(n1507), .A2(io_pmp_4_cfg_a[1]), .Y(n802) );
  AND2X1_LVT U902 ( .A1(n1490), .A2(io_bp_0_address[37]), .Y(n1644) );
  AND2X1_LVT U903 ( .A1(n1689), .A2(n_T_45[41]), .Y(n1009) );
  AND2X1_LVT U904 ( .A1(n1510), .A2(reg_dscratch[46]), .Y(n998) );
  AND3X1_LVT U905 ( .A1(n384), .A2(n379), .A3(n476), .Y(n674) );
  NAND2X0_LVT U906 ( .A1(n1508), .A2(reg_sscratch[46]), .Y(n482) );
  NAND3X0_LVT U907 ( .A1(n479), .A2(n481), .A3(n482), .Y(n1679) );
  NAND2X0_LVT U908 ( .A1(reg_stvec[2]), .A2(n1478), .Y(n483) );
  NAND3X0_LVT U909 ( .A1(n382), .A2(n471), .A3(n483), .Y(n1669) );
  NAND2X0_LVT U910 ( .A1(n1489), .A2(reg_mepc[30]), .Y(n485) );
  NAND3X0_LVT U911 ( .A1(n480), .A2(n484), .A3(n485), .Y(n1627) );
  NAND2X0_LVT U912 ( .A1(n1490), .A2(io_bp_0_address[5]), .Y(n486) );
  NAND3X0_LVT U913 ( .A1(n388), .A2(n469), .A3(n486), .Y(n1540) );
  NAND2X0_LVT U914 ( .A1(read_mideleg_5), .A2(n1539), .Y(n487) );
  INVX1_LVT U915 ( .A(io_rw_addr[5]), .Y(n1517) );
  INVX1_LVT U916 ( .A(io_rw_addr[6]), .Y(n1516) );
  NOR2X0_LVT U917 ( .A1(io_rw_addr[8]), .A2(n605), .Y(n595) );
  AND3X1_LVT U918 ( .A1(n1557), .A2(n1529), .A3(n595), .Y(n1511) );
  AND2X1_LVT U919 ( .A1(n1516), .A2(io_rw_addr[9]), .Y(n615) );
  AND4X1_LVT U920 ( .A1(n615), .A2(io_rw_addr[11]), .A3(io_rw_addr[8]), .A4(
        n1514), .Y(n596) );
  AND2X1_LVT U921 ( .A1(n1520), .A2(io_rw_addr[1]), .Y(n671) );
  AND2X1_LVT U922 ( .A1(n1519), .A2(io_rw_addr[0]), .Y(n610) );
  OR2X1_LVT U923 ( .A1(io_rw_cmd[1]), .A2(io_rw_cmd[0]), .Y(n597) );
  AND3X1_LVT U924 ( .A1(n1134), .A2(io_rw_addr[9]), .A3(n1519), .Y(n599) );
  OA21X1_LVT U925 ( .A1(n1918), .A2(n599), .A3(n590), .Y(N1693) );
  NAND2X0_LVT U926 ( .A1(n1162), .A2(io_time[11]), .Y(n609) );
  NAND2X0_LVT U927 ( .A1(io_pmp_1_cfg_a[0]), .A2(n1507), .Y(n604) );
  AOI22X1_LVT U928 ( .A1(n1689), .A2(n_T_45[11]), .A3(n1510), .A4(
        reg_dscratch[11]), .Y(n603) );
  NAND4X0_LVT U929 ( .A1(n1513), .A2(io_rw_addr[7]), .A3(n1522), .A4(n445), 
        .Y(n601) );
  AOI22X1_LVT U930 ( .A1(n1493), .A2(reg_dpc[11]), .A3(n488), .A4(
        io_ptbr_ppn[11]), .Y(n602) );
  AND3X1_LVT U931 ( .A1(n604), .A2(n603), .A3(n602), .Y(n608) );
  NAND2X0_LVT U932 ( .A1(reg_stvec[11]), .A2(n1487), .Y(n607) );
  AND2X1_LVT U933 ( .A1(n1526), .A2(io_rw_addr[10]), .Y(n640) );
  AND2X1_LVT U934 ( .A1(n671), .A2(n1518), .Y(n857) );
  NAND2X0_LVT U935 ( .A1(io_bp_0_address[11]), .A2(n1490), .Y(n606) );
  NAND4X0_LVT U936 ( .A1(n609), .A2(n608), .A3(n607), .A4(n606), .Y(n614) );
  AND2X1_LVT U937 ( .A1(n630), .A2(io_rw_addr[2]), .Y(n1505) );
  AO22X1_LVT U938 ( .A1(n1479), .A2(io_pmp_7_addr[11]), .A3(n1491), .A4(
        io_pmp_4_addr[11]), .Y(n613) );
  AND2X1_LVT U939 ( .A1(n610), .A2(io_rw_addr[2]), .Y(n621) );
  AO22X1_LVT U940 ( .A1(n1480), .A2(io_pmp_0_addr[11]), .A3(n1472), .A4(
        io_pmp_5_addr[11]), .Y(n612) );
  AND3X1_LVT U941 ( .A1(n1518), .A2(io_rw_addr[1]), .A3(io_rw_addr[0]), .Y(
        n676) );
  AO22X1_LVT U942 ( .A1(n1492), .A2(io_pmp_2_addr[11]), .A3(n1473), .A4(
        io_pmp_3_addr[11]), .Y(n611) );
  NOR4X1_LVT U943 ( .A1(n614), .A2(n613), .A3(n612), .A4(n611), .Y(n628) );
  AND2X1_LVT U944 ( .A1(n620), .A2(n857), .Y(n1161) );
  AND2X1_LVT U945 ( .A1(n1527), .A2(n615), .Y(n858) );
  NAND2X0_LVT U946 ( .A1(n858), .A2(n1512), .Y(n1041) );
  AO22X1_LVT U947 ( .A1(n1474), .A2(io_interrupts_meip), .A3(n1157), .A4(
        n[1930]), .Y(n618) );
  AND2X1_LVT U948 ( .A1(n671), .A2(io_rw_addr[2]), .Y(n662) );
  AO22X1_LVT U949 ( .A1(n1494), .A2(io_pmp_6_addr[11]), .A3(n1496), .A4(
        io_pmp_1_addr[11]), .Y(n617) );
  NOR3X0_LVT U950 ( .A1(n619), .A2(n618), .A3(n617), .Y(n627) );
  AO22X1_LVT U951 ( .A1(n1485), .A2(reg_mscratch[11]), .A3(n1489), .A4(
        reg_mepc[11]), .Y(n625) );
  AO22X1_LVT U952 ( .A1(n1160), .A2(n_T_444[11]), .A3(n1497), .A4(
        reg_mtvec[11]), .Y(n624) );
  AND2X1_LVT U953 ( .A1(n1509), .A2(n857), .Y(n1168) );
  AO22X1_LVT U954 ( .A1(n1506), .A2(reg_sepc[11]), .A3(n1502), .A4(reg_mie[11]), .Y(n622) );
  NOR4X1_LVT U955 ( .A1(n625), .A2(n624), .A3(n623), .A4(n622), .Y(n626) );
  NAND3X0_LVT U956 ( .A1(n628), .A2(n627), .A3(n626), .Y(io_rw_rdata[11]) );
  INVX1_LVT U957 ( .A(n1674), .Y(n672) );
  NAND3X0_LVT U958 ( .A1(n503), .A2(n672), .A3(n630), .Y(n629) );
  AND2X1_LVT U959 ( .A1(n1142), .A2(io_time[2]), .Y(n1144) );
  AO22X1_LVT U960 ( .A1(n498), .A2(n_T_52[5]), .A3(wdata[11]), .A4(n1149), .Y(
        N1896) );
  NAND2X0_LVT U961 ( .A1(n504), .A2(n1168), .Y(n1455) );
  AND2X1_LVT U962 ( .A1(n1455), .A2(n1139), .Y(n1501) );
  AND2X1_LVT U963 ( .A1(n1501), .A2(n1697), .Y(n1500) );
  NAND2X0_LVT U964 ( .A1(n504), .A2(n1161), .Y(n1460) );
  AND2X1_LVT U965 ( .A1(n1139), .A2(n590), .Y(n1499) );
  AO22X1_LVT U966 ( .A1(n1151), .A2(wdata[11]), .A3(io_tval[11]), .A4(n1152), 
        .Y(N1004) );
  AO22X1_LVT U967 ( .A1(n1158), .A2(wdata[11]), .A3(io_tval[11]), .A4(n1159), 
        .Y(N1393) );
  NAND2X0_LVT U968 ( .A1(io_pmp_1_cfg_l), .A2(n1507), .Y(n632) );
  NAND2X0_LVT U969 ( .A1(n1493), .A2(reg_dpc[15]), .Y(n631) );
  AO22X1_LVT U970 ( .A1(n1150), .A2(n_T_52[9]), .A3(wdata[15]), .A4(n1149), 
        .Y(N1900) );
  AO22X1_LVT U971 ( .A1(n1152), .A2(io_tval[15]), .A3(wdata[15]), .A4(n1151), 
        .Y(N1008) );
  AO22X1_LVT U972 ( .A1(n1159), .A2(io_tval[15]), .A3(wdata[15]), .A4(n1158), 
        .Y(N1397) );
  MUX21X1_LVT U973 ( .A1(io_pc[15]), .A2(wdata[15]), .S0(n515), .Y(net35259)
         );
  MUX21X1_LVT U974 ( .A1(io_pc[15]), .A2(wdata[15]), .S0(n514), .Y(net35037)
         );
  NOR3X0_LVT U975 ( .A1(n1651), .A2(n1654), .A3(n1652), .Y(n652) );
  AO22X1_LVT U976 ( .A1(n1160), .A2(n_T_444[0]), .A3(n1497), .A4(n416), .Y(
        n649) );
  AO22X1_LVT U977 ( .A1(n1168), .A2(reg_scause[0]), .A3(n1162), .A4(io_time[0]), .Y(n648) );
  AND2X1_LVT U978 ( .A1(n858), .A2(n716), .Y(n1452) );
  AO22X1_LVT U979 ( .A1(n1153), .A2(n_T_383[0]), .A3(n1452), .A4(
        io_status_isa_0_), .Y(n646) );
  AND3X1_LVT U980 ( .A1(n1527), .A2(n633), .A3(n662), .Y(n1465) );
  NAND2X0_LVT U981 ( .A1(n1520), .A2(n1656), .Y(n637) );
  AOI22X1_LVT U982 ( .A1(n1689), .A2(n_T_45[0]), .A3(n1510), .A4(
        reg_dscratch[0]), .Y(n636) );
  AOI22X1_LVT U983 ( .A1(n1495), .A2(n_T_389_0), .A3(n488), .A4(io_ptbr_ppn[0]), .Y(n635) );
  NAND2X0_LVT U984 ( .A1(n1507), .A2(io_pmp_0_cfg_r), .Y(n634) );
  NAND4X0_LVT U985 ( .A1(n637), .A2(n636), .A3(n635), .A4(n634), .Y(n638) );
  AO21X1_LVT U986 ( .A1(read_scounteren[0]), .A2(n1465), .A3(n638), .Y(n639)
         );
  AO21X1_LVT U987 ( .A1(n1161), .A2(reg_mcause[0]), .A3(n639), .Y(n645) );
  NAND2X0_LVT U988 ( .A1(io_pmp_0_addr[0]), .A2(n1480), .Y(n643) );
  AOI22X1_LVT U989 ( .A1(n1481), .A2(io_bp_0_control_r), .A3(n1490), .A4(
        io_bp_0_address[0]), .Y(n642) );
  AND3X1_LVT U990 ( .A1(n1511), .A2(n1514), .A3(n1513), .Y(n1486) );
  AND2X1_LVT U991 ( .A1(n1486), .A2(io_rw_addr[0]), .Y(n1167) );
  AND2X1_LVT U992 ( .A1(n1486), .A2(n671), .Y(n1466) );
  AOI22X1_LVT U993 ( .A1(n1167), .A2(read_fcsr[0]), .A3(n1466), .A4(
        io_fcsr_rm[0]), .Y(n641) );
  NAND3X0_LVT U994 ( .A1(n643), .A2(n642), .A3(n641), .Y(n644) );
  OR3X1_LVT U995 ( .A1(n646), .A2(n645), .A3(n644), .Y(n647) );
  NOR4X1_LVT U996 ( .A1(n649), .A2(n648), .A3(n1655), .A4(n647), .Y(n651) );
  NAND3X0_LVT U997 ( .A1(n652), .A2(n651), .A3(n650), .Y(io_rw_rdata[0]) );
  NAND2X0_LVT U998 ( .A1(n1167), .A2(n504), .Y(n1163) );
  AND2X1_LVT U999 ( .A1(io_fcsr_flags_valid), .A2(n1163), .Y(n1164) );
  MUX21X1_LVT U1000 ( .A1(wdata[0]), .A2(read_fcsr[0]), .S0(n1163), .Y(n653)
         );
  AO21X1_LVT U1001 ( .A1(n1164), .A2(io_fcsr_flags_bits[0]), .A3(n653), .Y(
        n_GEN_345[0]) );
  NAND3X0_LVT U1002 ( .A1(n1517), .A2(n1518), .A3(io_rw_addr[8]), .Y(n654) );
  NAND2X0_LVT U1003 ( .A1(n654), .A2(n1514), .Y(n655) );
  AOI22X1_LVT U1004 ( .A1(n1160), .A2(n_T_444[2]), .A3(n1168), .A4(
        reg_scause[2]), .Y(n661) );
  AOI22X1_LVT U1005 ( .A1(n1510), .A2(reg_dscratch[2]), .A3(n1493), .A4(
        reg_dpc[2]), .Y(n660) );
  NAND2X0_LVT U1006 ( .A1(io_status_isa_2_), .A2(n1452), .Y(n657) );
  NAND2X0_LVT U1007 ( .A1(io_pmp_2_addr[2]), .A2(n1492), .Y(n656) );
  NAND4X0_LVT U1008 ( .A1(n661), .A2(n660), .A3(n657), .A4(n656), .Y(n666) );
  AO22X1_LVT U1009 ( .A1(n1153), .A2(n_T_383[2]), .A3(n1161), .A4(
        reg_mcause[2]), .Y(n664) );
  AND2X1_LVT U1010 ( .A1(n858), .A2(n662), .Y(n1484) );
  AO22X1_LVT U1011 ( .A1(n1485), .A2(reg_mscratch[2]), .A3(read_mcounteren[2]), 
        .A4(n1484), .Y(n663) );
  OR3X1_LVT U1012 ( .A1(n664), .A2(n663), .A3(n1659), .Y(n665) );
  NOR4X1_LVT U1013 ( .A1(n1660), .A2(n1658), .A3(n666), .A4(n665), .Y(n667) );
  NAND2X0_LVT U1014 ( .A1(n1671), .A2(n667), .Y(io_rw_rdata[2]) );
  NAND2X0_LVT U1015 ( .A1(io_rw_rdata[2]), .A2(n589), .Y(n668) );
  AND2X1_LVT U1016 ( .A1(io_cause[2]), .A2(n1697), .Y(n1220) );
  NAND2X0_LVT U1017 ( .A1(n1161), .A2(n503), .Y(n701) );
  AO22X1_LVT U1018 ( .A1(io_tval[2]), .A2(n1152), .A3(wdata[2]), .A4(n1151), 
        .Y(N995) );
  AO22X1_LVT U1019 ( .A1(io_tval[2]), .A2(n1159), .A3(wdata[2]), .A4(n1158), 
        .Y(N1384) );
  MUX21X1_LVT U1020 ( .A1(io_pc[2]), .A2(wdata[2]), .S0(n515), .Y(net35298) );
  AND2X1_LVT U1021 ( .A1(io_status_debug_BAR), .A2(n_T_389_2), .Y(
        io_singleStep) );
  INVX1_LVT U1022 ( .A(n1670), .Y(n1083) );
  AO22X1_LVT U1023 ( .A1(n1150), .A2(n_T_52[6]), .A3(wdata[12]), .A4(n1149), 
        .Y(N1897) );
  AO22X1_LVT U1024 ( .A1(io_tval[12]), .A2(n1152), .A3(wdata[12]), .A4(n1151), 
        .Y(N1005) );
  AO22X1_LVT U1025 ( .A1(io_tval[12]), .A2(n1159), .A3(wdata[12]), .A4(n1158), 
        .Y(N1394) );
  AND2X1_LVT U1026 ( .A1(n_T_45[1]), .A2(n_T_45[0]), .Y(n670) );
  AND2X1_LVT U1027 ( .A1(io_retire), .A2(n670), .Y(n956) );
  AND2X1_LVT U1028 ( .A1(n956), .A2(n_T_45[2]), .Y(n959) );
  AND2X1_LVT U1029 ( .A1(n959), .A2(n_T_45[3]), .Y(n960) );
  AND2X1_LVT U1030 ( .A1(n960), .A2(n_T_45[4]), .Y(n1459) );
  AND2X1_LVT U1031 ( .A1(n957), .A2(n590), .Y(n961) );
  AO22X1_LVT U1032 ( .A1(n495), .A2(n_T_44[6]), .A3(wdata[12]), .A4(n491), .Y(
        N1503) );
  AND2X1_LVT U1033 ( .A1(n1167), .A2(io_rw_addr[1]), .Y(n1477) );
  INVX1_LVT U1034 ( .A(n1477), .Y(n1696) );
  AND2X1_LVT U1035 ( .A1(n1487), .A2(n658), .Y(n1478) );
  NAND3X0_LVT U1036 ( .A1(n1544), .A2(n674), .A3(n380), .Y(n675) );
  OR2X1_LVT U1037 ( .A1(n675), .A2(n1543), .Y(io_rw_rdata[5]) );
  NAND2X0_LVT U1038 ( .A1(n676), .A2(n858), .Y(n1553) );
  NAND2X0_LVT U1039 ( .A1(n1935), .A2(n1154), .Y(n681) );
  AO21X1_LVT U1040 ( .A1(n_T_45[1]), .A2(n1689), .A3(n1554), .Y(n677) );
  AOI21X1_LVT U1041 ( .A1(n1495), .A2(n_T_389_1), .A3(n677), .Y(n680) );
  NAND2X0_LVT U1042 ( .A1(n1481), .A2(io_bp_0_control_w), .Y(n679) );
  NAND2X0_LVT U1043 ( .A1(n1507), .A2(io_pmp_0_cfg_w), .Y(n678) );
  NAND4X0_LVT U1044 ( .A1(n681), .A2(n680), .A3(n679), .A4(n678), .Y(n687) );
  AO22X1_LVT U1045 ( .A1(n1490), .A2(io_bp_0_address[1]), .A3(n1167), .A4(
        read_fcsr[1]), .Y(n682) );
  AO21X1_LVT U1046 ( .A1(n1153), .A2(n_T_383[1]), .A3(n682), .Y(n686) );
  AO22X1_LVT U1047 ( .A1(n1161), .A2(reg_mcause[1]), .A3(n1484), .A4(
        read_mcounteren[1]), .Y(n685) );
  NAND3X0_LVT U1048 ( .A1(n1553), .A2(n1552), .A3(n1692), .Y(n683) );
  AND2X1_LVT U1049 ( .A1(n683), .A2(read_mideleg_1), .Y(n684) );
  NOR4X1_LVT U1050 ( .A1(n687), .A2(n686), .A3(n685), .A4(n684), .Y(n696) );
  NAND2X0_LVT U1051 ( .A1(n1162), .A2(io_time[1]), .Y(n691) );
  NAND2X0_LVT U1052 ( .A1(n1160), .A2(n_T_444[1]), .Y(n690) );
  NAND2X0_LVT U1053 ( .A1(n1168), .A2(reg_scause[1]), .Y(n689) );
  NAND2X0_LVT U1054 ( .A1(n1508), .A2(reg_sscratch[1]), .Y(n688) );
  NAND4X0_LVT U1055 ( .A1(n691), .A2(n690), .A3(n689), .A4(n688), .Y(n692) );
  NOR4X1_LVT U1056 ( .A1(n692), .A2(n1546), .A3(n1547), .A4(n1545), .Y(n695)
         );
  AO222X1_LVT U1057 ( .A1(n1493), .A2(reg_dpc[1]), .A3(n1506), .A4(reg_sepc[1]), .A5(reg_mepc[1]), .A6(n1489), .Y(n693) );
  NAND2X0_LVT U1058 ( .A1(n693), .A2(io_status_isa_2_), .Y(n694) );
  NAND4X0_LVT U1059 ( .A1(n1555), .A2(n696), .A3(n695), .A4(n694), .Y(
        io_rw_rdata[1]) );
  AND2X1_LVT U1060 ( .A1(n697), .A2(n589), .Y(n1476) );
  MUX21X1_LVT U1061 ( .A1(wdata[1]), .A2(read_fcsr[1]), .S0(n1163), .Y(n698)
         );
  AO21X1_LVT U1062 ( .A1(n1164), .A2(io_fcsr_flags_bits[1]), .A3(n698), .Y(
        n_GEN_345[1]) );
  OR2X1_LVT U1063 ( .A1(io_status_prv[1]), .A2(io_rw_addr[0]), .Y(n700) );
  AO222X1_LVT U1064 ( .A1(n700), .A2(n699), .A3(wdata[1]), .A4(n923), .A5(
        n1500), .A6(io_cause[1]), .Y(N1271) );
  INVX1_LVT U1065 ( .A(n701), .Y(n955) );
  AO22X1_LVT U1066 ( .A1(n1498), .A2(n1209), .A3(wdata[1]), .A4(n955), .Y(N882) );
  NAND2X0_LVT U1067 ( .A1(n503), .A2(n1154), .Y(n702) );
  NAND2X0_LVT U1068 ( .A1(n590), .A2(n702), .Y(N290) );
  NAND2X0_LVT U1069 ( .A1(n500), .A2(n590), .Y(n917) );
  INVX1_LVT U1070 ( .A(N290), .Y(n1443) );
  INVX1_LVT U1071 ( .A(n917), .Y(n883) );
  AO22X1_LVT U1072 ( .A1(n1933), .A2(n883), .A3(wdata[1]), .A4(n949), .Y(n1062) );
  AO22X1_LVT U1073 ( .A1(wdata[1]), .A2(n1151), .A3(io_tval[1]), .A4(n1152), 
        .Y(N994) );
  AO22X1_LVT U1074 ( .A1(wdata[1]), .A2(n1158), .A3(io_tval[1]), .A4(n1159), 
        .Y(N1383) );
  AND2X1_LVT U1075 ( .A1(n381), .A2(n_T_1155[0]), .Y(n704) );
  MUX21X1_LVT U1076 ( .A1(n_T_1155[1]), .A2(n_T_1155_3), .S0(io_status_prv[1]), 
        .Y(n703) );
  MUX21X1_LVT U1077 ( .A1(n704), .A2(n703), .S0(io_status_prv[0]), .Y(n705) );
  NAND2X0_LVT U1078 ( .A1(n1210), .A2(n705), .Y(n706) );
  NAND3X0_LVT U1079 ( .A1(n706), .A2(n860), .A3(io_status_debug_BAR), .Y(n708)
         );
  AND2X1_LVT U1080 ( .A1(n707), .A2(n1226), .Y(n1467) );
  NAND3X0_LVT U1081 ( .A1(n1257), .A2(io_status_debug_BAR), .A3(n1139), .Y(
        n1448) );
  NAND2X0_LVT U1082 ( .A1(n1448), .A2(n590), .Y(N467) );
  NAND2X0_LVT U1083 ( .A1(n504), .A2(n1495), .Y(n1449) );
  INVX1_LVT U1084 ( .A(n1449), .Y(n932) );
  OR2X1_LVT U1085 ( .A1(n932), .A2(N467), .Y(n935) );
  NAND2X0_LVT U1086 ( .A1(n935), .A2(n590), .Y(n934) );
  AND2X1_LVT U1087 ( .A1(wdata[0]), .A2(wdata[1]), .Y(n709) );
  MUX21X1_LVT U1088 ( .A1(n709), .A2(io_status_prv[1]), .S0(n1449), .Y(n710)
         );
  OA22X1_LVT U1089 ( .A1(n_T_389_1), .A2(n935), .A3(n934), .A4(n710), .Y(n2155) );
  AO21X1_LVT U1090 ( .A1(n_T_45[0]), .A2(io_retire), .A3(n_T_45[1]), .Y(n711)
         );
  AO22X1_LVT U1091 ( .A1(n712), .A2(n711), .A3(wdata[1]), .A4(n491), .Y(N1429)
         );
  AND2X1_LVT U1092 ( .A1(n1509), .A2(n1505), .Y(n1475) );
  INVX1_LVT U1093 ( .A(n1475), .Y(n1898) );
  INVX1_LVT U1094 ( .A(n1474), .Y(n1899) );
  AND2X1_LVT U1095 ( .A1(io_rw_wdata[9]), .A2(n516), .Y(n714) );
  NAND2X0_LVT U1096 ( .A1(n1474), .A2(n1908), .Y(n713) );
  AO22X1_LVT U1097 ( .A1(n1474), .A2(n714), .A3(n_T_3694_9_), .A4(n713), .Y(
        n200) );
  AO22X1_LVT U1098 ( .A1(n1502), .A2(reg_mie[9]), .A3(n1162), .A4(io_time[9]), 
        .Y(n728) );
  AO22X1_LVT U1099 ( .A1(n1491), .A2(io_pmp_4_addr[9]), .A3(n1480), .A4(
        io_pmp_0_addr[9]), .Y(n727) );
  NAND2X0_LVT U1100 ( .A1(io_pmp_7_addr[9]), .A2(n1479), .Y(n724) );
  NAND2X0_LVT U1101 ( .A1(n1507), .A2(io_pmp_1_cfg_w), .Y(n720) );
  AOI22X1_LVT U1102 ( .A1(n1493), .A2(reg_dpc[9]), .A3(n1488), .A4(
        io_ptbr_ppn[9]), .Y(n719) );
  AND2X1_LVT U1103 ( .A1(io_rw_addr[10]), .A2(io_rw_addr[9]), .Y(n942) );
  AND4X1_LVT U1104 ( .A1(n1513), .A2(io_rw_addr[7]), .A3(io_rw_addr[6]), .A4(
        n1522), .Y(n715) );
  NAND3X0_LVT U1105 ( .A1(n716), .A2(n942), .A3(n715), .Y(n866) );
  AOI22X1_LVT U1106 ( .A1(n1689), .A2(n_T_45[9]), .A3(n1510), .A4(
        reg_dscratch[9]), .Y(n717) );
  OA21X1_LVT U1107 ( .A1(n1912), .A2(n866), .A3(n717), .Y(n718) );
  AND3X1_LVT U1108 ( .A1(n720), .A2(n719), .A3(n718), .Y(n723) );
  NAND2X0_LVT U1109 ( .A1(reg_stvec[9]), .A2(n1487), .Y(n722) );
  NAND2X0_LVT U1110 ( .A1(n1490), .A2(io_bp_0_address[9]), .Y(n721) );
  NAND4X0_LVT U1111 ( .A1(n724), .A2(n723), .A3(n722), .A4(n721), .Y(n726) );
  AO22X1_LVT U1112 ( .A1(n1472), .A2(io_pmp_5_addr[9]), .A3(n1473), .A4(
        io_pmp_3_addr[9]), .Y(n725) );
  NOR4X1_LVT U1113 ( .A1(n728), .A2(n727), .A3(n726), .A4(n725), .Y(n741) );
  AOI22X1_LVT U1114 ( .A1(n1492), .A2(io_pmp_2_addr[9]), .A3(n1494), .A4(
        io_pmp_6_addr[9]), .Y(n734) );
  AND2X1_LVT U1115 ( .A1(n1504), .A2(n1515), .Y(n1503) );
  NAND2X0_LVT U1116 ( .A1(reg_mie[9]), .A2(n1503), .Y(n742) );
  NAND2X0_LVT U1117 ( .A1(n1136), .A2(n1475), .Y(n729) );
  NAND3X0_LVT U1118 ( .A1(n742), .A2(n1553), .A3(n729), .Y(n730) );
  NAND2X0_LVT U1119 ( .A1(read_mideleg_9_), .A2(n730), .Y(n732) );
  NAND2X0_LVT U1120 ( .A1(io_pmp_1_addr[9]), .A2(n1496), .Y(n731) );
  AND4X1_LVT U1121 ( .A1(n734), .A2(n733), .A3(n732), .A4(n731), .Y(n740) );
  AO22X1_LVT U1122 ( .A1(n1485), .A2(reg_mscratch[9]), .A3(n1489), .A4(
        reg_mepc[9]), .Y(n738) );
  AO22X1_LVT U1123 ( .A1(n1160), .A2(n_T_444[9]), .A3(n1497), .A4(reg_mtvec[9]), .Y(n737) );
  AO22X1_LVT U1124 ( .A1(n1508), .A2(reg_sscratch[9]), .A3(n1506), .A4(
        reg_sepc[9]), .Y(n735) );
  NOR4X1_LVT U1125 ( .A1(n738), .A2(n737), .A3(n736), .A4(n735), .Y(n739) );
  NAND3X0_LVT U1126 ( .A1(n741), .A2(n740), .A3(n739), .Y(io_rw_rdata[9]) );
  NAND2X0_LVT U1127 ( .A1(n503), .A2(n743), .Y(n879) );
  AO22X1_LVT U1128 ( .A1(n498), .A2(n_T_52[3]), .A3(wdata[9]), .A4(n1149), .Y(
        N1894) );
  AO22X1_LVT U1129 ( .A1(n1151), .A2(wdata[9]), .A3(io_tval[9]), .A4(n1152), 
        .Y(N1002) );
  AO22X1_LVT U1130 ( .A1(n1158), .A2(wdata[9]), .A3(io_tval[9]), .A4(n1159), 
        .Y(N1391) );
  NAND3X0_LVT U1131 ( .A1(n463), .A2(io_pmp_2_cfg_l), .A3(io_pmp_2_cfg_a[0]), 
        .Y(n744) );
  MUX21X1_LVT U1132 ( .A1(io_pmp_1_addr[9]), .A2(wdata[9]), .S0(n506), .Y(
        n_GEN_265[9]) );
  MUX21X1_LVT U1133 ( .A1(io_pc[9]), .A2(wdata[9]), .S0(n513), .Y(net34853) );
  NAND2X0_LVT U1134 ( .A1(n_T_444[39]), .A2(n1160), .Y(n748) );
  AOI21X1_LVT U1135 ( .A1(n1493), .A2(reg_dpc[39]), .A3(n1649), .Y(n747) );
  NAND2X0_LVT U1136 ( .A1(n_T_383[39]), .A2(n1153), .Y(n746) );
  NAND3X0_LVT U1137 ( .A1(n748), .A2(n747), .A3(n746), .Y(n749) );
  AOI22X1_LVT U1138 ( .A1(n1508), .A2(reg_sscratch[39]), .A3(n1162), .A4(n1960), .Y(n753) );
  AO22X1_LVT U1139 ( .A1(n1689), .A2(n_T_45[39]), .A3(n1510), .A4(
        reg_dscratch[39]), .Y(n750) );
  AOI21X1_LVT U1140 ( .A1(n1507), .A2(io_pmp_4_cfg_l), .A3(n750), .Y(n751) );
  OR2X1_LVT U1141 ( .A1(n754), .A2(n1690), .Y(io_rw_rdata[39]) );
  AO22X1_LVT U1142 ( .A1(n1149), .A2(wdata[39]), .A3(n_T_52[33]), .A4(n496), 
        .Y(N1924) );
  AO22X1_LVT U1143 ( .A1(n492), .A2(wdata[39]), .A3(n_T_44[33]), .A4(n495), 
        .Y(N1530) );
  AO22X1_LVT U1144 ( .A1(wdata[39]), .A2(n1151), .A3(io_tval[39]), .A4(n1152), 
        .Y(N1032) );
  MUX21X1_LVT U1145 ( .A1(io_pc[39]), .A2(wdata[39]), .S0(n515), .Y(net35187)
         );
  AO22X1_LVT U1146 ( .A1(wdata[39]), .A2(n1158), .A3(io_tval[39]), .A4(n1159), 
        .Y(N1421) );
  AOI22X1_LVT U1147 ( .A1(n1508), .A2(reg_sscratch[55]), .A3(n1162), .A4(n1944), .Y(n757) );
  AO22X1_LVT U1148 ( .A1(n1689), .A2(n_T_45[55]), .A3(n1510), .A4(
        reg_dscratch[55]), .Y(n755) );
  NAND4X0_LVT U1149 ( .A1(n968), .A2(n757), .A3(n473), .A4(n756), .Y(
        io_rw_rdata[55]) );
  AO22X1_LVT U1150 ( .A1(n1149), .A2(wdata[55]), .A3(n_T_52[49]), .A4(n496), 
        .Y(N1940) );
  AO22X1_LVT U1151 ( .A1(n492), .A2(wdata[55]), .A3(n_T_44[49]), .A4(n494), 
        .Y(N1546) );
  NAND2X0_LVT U1152 ( .A1(n1510), .A2(reg_dscratch[13]), .Y(n758) );
  NAND2X0_LVT U1153 ( .A1(n1928), .A2(n1154), .Y(n1155) );
  AO22X1_LVT U1154 ( .A1(n1150), .A2(n_T_52[7]), .A3(wdata[13]), .A4(n1149), 
        .Y(N1898) );
  AO22X1_LVT U1155 ( .A1(n1152), .A2(io_tval[13]), .A3(wdata[13]), .A4(n1151), 
        .Y(N1006) );
  AO22X1_LVT U1156 ( .A1(n1159), .A2(io_tval[13]), .A3(wdata[13]), .A4(n1158), 
        .Y(N1395) );
  AO22X1_LVT U1157 ( .A1(n493), .A2(n_T_44[7]), .A3(wdata[13]), .A4(n491), .Y(
        N1504) );
  AO22X1_LVT U1158 ( .A1(n1150), .A2(n_T_52[8]), .A3(wdata[14]), .A4(n1149), 
        .Y(N1899) );
  AO22X1_LVT U1159 ( .A1(n1152), .A2(io_tval[14]), .A3(wdata[14]), .A4(n1151), 
        .Y(N1007) );
  AO22X1_LVT U1160 ( .A1(n1159), .A2(io_tval[14]), .A3(wdata[14]), .A4(n1158), 
        .Y(N1396) );
  MUX21X1_LVT U1161 ( .A1(io_pc[14]), .A2(wdata[14]), .S0(n514), .Y(net35040)
         );
  INVX1_LVT U1162 ( .A(wdata[14]), .Y(n51) );
  AO22X1_LVT U1163 ( .A1(n1129), .A2(n_T_44[8]), .A3(wdata[14]), .A4(n491), 
        .Y(N1505) );
  AOI22X1_LVT U1164 ( .A1(n1161), .A2(reg_mcause[63]), .A3(n1168), .A4(
        reg_scause[63]), .Y(n765) );
  AOI22X1_LVT U1165 ( .A1(n1689), .A2(n_T_45[63]), .A3(n1510), .A4(
        reg_dscratch[63]), .Y(n761) );
  NAND2X0_LVT U1166 ( .A1(n1507), .A2(io_pmp_7_cfg_l), .Y(n760) );
  NAND2X0_LVT U1167 ( .A1(n488), .A2(io_ptbr_mode[3]), .Y(n759) );
  AND4X1_LVT U1168 ( .A1(n1155), .A2(n761), .A3(n760), .A4(n759), .Y(n764) );
  NAND2X0_LVT U1169 ( .A1(n1452), .A2(n_T_3678_63_), .Y(n763) );
  NAND2X0_LVT U1170 ( .A1(n1162), .A2(n1936), .Y(n762) );
  NAND4X0_LVT U1171 ( .A1(n765), .A2(n764), .A3(n763), .A4(n762), .Y(n766) );
  OR3X1_LVT U1172 ( .A1(n766), .A2(n1672), .A3(n1690), .Y(io_rw_rdata[63]) );
  AND2X1_LVT U1173 ( .A1(io_cause[63]), .A2(n1697), .Y(n1201) );
  AO22X1_LVT U1174 ( .A1(n1501), .A2(n1201), .A3(wdata[63]), .A4(n923), .Y(
        N1333) );
  AO22X1_LVT U1175 ( .A1(n1498), .A2(n1201), .A3(wdata[63]), .A4(n955), .Y(
        N944) );
  AO21X1_LVT U1176 ( .A1(n_T_3678_63_), .A2(n504), .A3(n376), .Y(N1622) );
  AOI22X1_LVT U1177 ( .A1(n1689), .A2(n_T_45[59]), .A3(n1510), .A4(
        reg_dscratch[59]), .Y(n769) );
  NAND2X0_LVT U1178 ( .A1(n1481), .A2(n_T_366_59_), .Y(n768) );
  NAND2X0_LVT U1179 ( .A1(n1507), .A2(io_pmp_7_cfg_a[0]), .Y(n767) );
  AO22X1_LVT U1180 ( .A1(n1508), .A2(reg_sscratch[59]), .A3(n1162), .A4(n1940), 
        .Y(n770) );
  OR3X1_LVT U1181 ( .A1(n772), .A2(n771), .A3(n770), .Y(n773) );
  OR2X1_LVT U1182 ( .A1(n773), .A2(n1690), .Y(io_rw_rdata[59]) );
  AO22X1_LVT U1183 ( .A1(n1149), .A2(wdata[59]), .A3(n_T_52[53]), .A4(n496), 
        .Y(N1944) );
  AO22X1_LVT U1184 ( .A1(n1128), .A2(wdata[59]), .A3(n_T_44[53]), .A4(n495), 
        .Y(N1550) );
  AOI22X1_LVT U1185 ( .A1(n1508), .A2(reg_sscratch[60]), .A3(n1162), .A4(n1939), .Y(n777) );
  AO22X1_LVT U1186 ( .A1(n1689), .A2(n_T_45[60]), .A3(n1510), .A4(
        reg_dscratch[60]), .Y(n774) );
  AOI21X1_LVT U1187 ( .A1(n1507), .A2(io_pmp_7_cfg_a[1]), .A3(n774), .Y(n775)
         );
  OR2X1_LVT U1188 ( .A1(n778), .A2(n1690), .Y(io_rw_rdata[60]) );
  AO22X1_LVT U1189 ( .A1(n1149), .A2(wdata[60]), .A3(n_T_52[54]), .A4(n496), 
        .Y(N1945) );
  AO22X1_LVT U1190 ( .A1(n1128), .A2(wdata[60]), .A3(n_T_44[54]), .A4(n494), 
        .Y(N1551) );
  MUX21X1_LVT U1191 ( .A1(io_pmp_6_addr[9]), .A2(wdata[9]), .S0(n511), .Y(
        n_GEN_300[9]) );
  MUX21X1_LVT U1192 ( .A1(io_pc[9]), .A2(wdata[9]), .S0(n515), .Y(net35277) );
  AO22X1_LVT U1193 ( .A1(n1508), .A2(reg_sscratch[23]), .A3(n1162), .A4(
        io_time[23]), .Y(n787) );
  NAND2X0_LVT U1194 ( .A1(n1153), .A2(n_T_383[23]), .Y(n782) );
  AOI21X1_LVT U1195 ( .A1(n_T_45[23]), .A2(n1689), .A3(n1604), .Y(n781) );
  NAND2X0_LVT U1196 ( .A1(n1507), .A2(io_pmp_2_cfg_l), .Y(n780) );
  NAND2X0_LVT U1197 ( .A1(n1510), .A2(reg_dscratch[23]), .Y(n779) );
  NAND4X0_LVT U1198 ( .A1(n782), .A2(n781), .A3(n780), .A4(n779), .Y(n785) );
  AO22X1_LVT U1199 ( .A1(n1480), .A2(io_pmp_0_addr[23]), .A3(n1492), .A4(
        io_pmp_2_addr[23]), .Y(n783) );
  OR3X1_LVT U1200 ( .A1(n785), .A2(n784), .A3(n783), .Y(n786) );
  NOR4X1_LVT U1201 ( .A1(n788), .A2(n787), .A3(n786), .A4(n1602), .Y(n789) );
  NAND2X0_LVT U1202 ( .A1(n1605), .A2(n789), .Y(io_rw_rdata[23]) );
  AO22X1_LVT U1203 ( .A1(n1150), .A2(n_T_52[17]), .A3(wdata[23]), .A4(n1149), 
        .Y(N1908) );
  AO22X1_LVT U1204 ( .A1(n1152), .A2(io_tval[23]), .A3(wdata[23]), .A4(n1151), 
        .Y(N1016) );
  AO21X1_LVT U1205 ( .A1(n1919), .A2(n504), .A3(n376), .Y(N1582) );
  MUX21X1_LVT U1206 ( .A1(io_pc[23]), .A2(wdata[23]), .S0(n514), .Y(net35013)
         );
  AO22X1_LVT U1207 ( .A1(n493), .A2(n_T_44[17]), .A3(wdata[23]), .A4(n492), 
        .Y(N1514) );
  AO22X1_LVT U1208 ( .A1(n1149), .A2(wdata[31]), .A3(n_T_52[25]), .A4(n496), 
        .Y(N1916) );
  AO22X1_LVT U1209 ( .A1(n1151), .A2(wdata[31]), .A3(io_tval[31]), .A4(n1152), 
        .Y(N1024) );
  AO22X1_LVT U1210 ( .A1(n1158), .A2(wdata[31]), .A3(io_tval[31]), .A4(n1159), 
        .Y(N1413) );
  AO22X1_LVT U1211 ( .A1(n1128), .A2(wdata[31]), .A3(n_T_44[25]), .A4(n494), 
        .Y(N1522) );
  NAND2X0_LVT U1212 ( .A1(n1153), .A2(n_T_383[27]), .Y(n793) );
  AOI21X1_LVT U1213 ( .A1(n_T_45[27]), .A2(n1689), .A3(n1617), .Y(n792) );
  NAND2X0_LVT U1214 ( .A1(n1507), .A2(io_pmp_3_cfg_a[0]), .Y(n791) );
  NAND2X0_LVT U1215 ( .A1(n1493), .A2(reg_dpc[27]), .Y(n790) );
  NAND4X0_LVT U1216 ( .A1(n793), .A2(n792), .A3(n791), .A4(n790), .Y(n795) );
  NOR4X1_LVT U1217 ( .A1(n1619), .A2(n795), .A3(n794), .A4(n1618), .Y(n800) );
  AO22X1_LVT U1218 ( .A1(n1491), .A2(io_pmp_4_addr[27]), .A3(n1496), .A4(
        io_pmp_1_addr[27]), .Y(n796) );
  NOR3X0_LVT U1219 ( .A1(n797), .A2(n796), .A3(n1614), .Y(n799) );
  NOR2X0_LVT U1220 ( .A1(n1615), .A2(n1616), .Y(n798) );
  NAND4X0_LVT U1221 ( .A1(n800), .A2(n799), .A3(n798), .A4(n466), .Y(
        io_rw_rdata[27]) );
  AO22X1_LVT U1222 ( .A1(n1150), .A2(n_T_52[21]), .A3(wdata[27]), .A4(n1149), 
        .Y(N1912) );
  AO22X1_LVT U1223 ( .A1(n1152), .A2(io_tval[27]), .A3(wdata[27]), .A4(n1151), 
        .Y(N1020) );
  AO22X1_LVT U1224 ( .A1(n1159), .A2(io_tval[27]), .A3(wdata[27]), .A4(n1158), 
        .Y(N1409) );
  MUX21X1_LVT U1225 ( .A1(io_pc[27]), .A2(wdata[27]), .S0(n515), .Y(net35223)
         );
  AO22X1_LVT U1226 ( .A1(n495), .A2(n_T_44[21]), .A3(wdata[27]), .A4(n492), 
        .Y(N1518) );
  AO22X1_LVT U1227 ( .A1(n497), .A2(n_T_52[22]), .A3(wdata[28]), .A4(n1149), 
        .Y(N1913) );
  AO22X1_LVT U1228 ( .A1(n1152), .A2(io_tval[28]), .A3(wdata[28]), .A4(n1151), 
        .Y(N1021) );
  AO22X1_LVT U1229 ( .A1(n1159), .A2(io_tval[28]), .A3(wdata[28]), .A4(n1158), 
        .Y(N1410) );
  MUX21X1_LVT U1230 ( .A1(io_pc[28]), .A2(wdata[28]), .S0(n515), .Y(net35220)
         );
  AO22X1_LVT U1231 ( .A1(n493), .A2(n_T_44[22]), .A3(wdata[28]), .A4(n492), 
        .Y(N1519) );
  AO22X1_LVT U1232 ( .A1(n1149), .A2(wdata[35]), .A3(n_T_52[29]), .A4(n496), 
        .Y(N1920) );
  AO22X1_LVT U1233 ( .A1(wdata[35]), .A2(n1151), .A3(n1152), .A4(io_tval[35]), 
        .Y(N1028) );
  AO22X1_LVT U1234 ( .A1(wdata[35]), .A2(n1158), .A3(n1159), .A4(io_tval[35]), 
        .Y(N1417) );
  MUX21X1_LVT U1235 ( .A1(io_pc[35]), .A2(wdata[35]), .S0(n515), .Y(net35199)
         );
  MUX21X1_LVT U1236 ( .A1(io_pc[35]), .A2(wdata[35]), .S0(n514), .Y(net34977)
         );
  AO22X1_LVT U1237 ( .A1(n1128), .A2(wdata[35]), .A3(n_T_44[29]), .A4(n1129), 
        .Y(N1526) );
  AOI22X1_LVT U1238 ( .A1(n1153), .A2(n_T_383[36]), .A3(n1160), .A4(
        n_T_444[36]), .Y(n803) );
  NAND2X0_LVT U1239 ( .A1(n1162), .A2(n1963), .Y(n801) );
  NAND4X0_LVT U1240 ( .A1(n804), .A2(n803), .A3(n802), .A4(n801), .Y(n805) );
  OR2X1_LVT U1241 ( .A1(n805), .A2(n1643), .Y(io_rw_rdata[36]) );
  AO22X1_LVT U1242 ( .A1(n_T_52[30]), .A2(n1150), .A3(n1149), .A4(wdata[36]), 
        .Y(N1921) );
  AO22X1_LVT U1243 ( .A1(n1152), .A2(io_tval[36]), .A3(wdata[36]), .A4(n1151), 
        .Y(N1029) );
  AO22X1_LVT U1244 ( .A1(n1159), .A2(io_tval[36]), .A3(wdata[36]), .A4(n1158), 
        .Y(N1418) );
  MUX21X1_LVT U1245 ( .A1(io_pc[36]), .A2(wdata[36]), .S0(n513), .Y(net34772)
         );
  MUX21X1_LVT U1246 ( .A1(io_pmp_3_addr[9]), .A2(wdata[9]), .S0(n508), .Y(
        n_GEN_279[9]) );
  AOI22X1_LVT U1247 ( .A1(n1689), .A2(n_T_45[47]), .A3(n1507), .A4(
        io_pmp_5_cfg_l), .Y(n807) );
  NAND2X0_LVT U1248 ( .A1(n1162), .A2(n1952), .Y(n806) );
  NAND3X0_LVT U1249 ( .A1(n481), .A2(n1680), .A3(n809), .Y(io_rw_rdata[47]) );
  AO22X1_LVT U1250 ( .A1(n1149), .A2(wdata[47]), .A3(n_T_52[41]), .A4(n497), 
        .Y(N1932) );
  AO22X1_LVT U1251 ( .A1(n1128), .A2(wdata[47]), .A3(n_T_44[41]), .A4(n1129), 
        .Y(N1538) );
  AOI22X1_LVT U1252 ( .A1(n1689), .A2(n_T_45[51]), .A3(n1507), .A4(
        io_pmp_6_cfg_a[0]), .Y(n811) );
  NAND2X0_LVT U1253 ( .A1(n1162), .A2(n1948), .Y(n810) );
  NAND3X0_LVT U1254 ( .A1(n481), .A2(n1684), .A3(n813), .Y(io_rw_rdata[51]) );
  AO22X1_LVT U1255 ( .A1(n1149), .A2(wdata[51]), .A3(n_T_52[45]), .A4(n497), 
        .Y(N1936) );
  AO22X1_LVT U1256 ( .A1(n1128), .A2(wdata[51]), .A3(n_T_44[45]), .A4(n1129), 
        .Y(N1542) );
  AOI22X1_LVT U1257 ( .A1(n1689), .A2(n_T_45[52]), .A3(n1507), .A4(
        io_pmp_6_cfg_a[1]), .Y(n815) );
  NAND2X0_LVT U1258 ( .A1(n1162), .A2(n1947), .Y(n814) );
  NAND3X0_LVT U1259 ( .A1(n481), .A2(n1685), .A3(n817), .Y(io_rw_rdata[52]) );
  AO22X1_LVT U1260 ( .A1(n1149), .A2(wdata[52]), .A3(n_T_52[46]), .A4(n1150), 
        .Y(N1937) );
  AO22X1_LVT U1261 ( .A1(n1128), .A2(wdata[52]), .A3(n_T_44[46]), .A4(n1129), 
        .Y(N1543) );
  MUX21X1_LVT U1262 ( .A1(io_pmp_5_addr[9]), .A2(wdata[9]), .S0(n510), .Y(
        n_GEN_293[9]) );
  AOI22X1_LVT U1263 ( .A1(n1689), .A2(n_T_45[43]), .A3(n1507), .A4(
        io_pmp_5_cfg_a[0]), .Y(n819) );
  NAND2X0_LVT U1264 ( .A1(n1162), .A2(n1956), .Y(n818) );
  NAND3X0_LVT U1265 ( .A1(n481), .A2(n1678), .A3(n821), .Y(io_rw_rdata[43]) );
  AO22X1_LVT U1266 ( .A1(n1149), .A2(wdata[43]), .A3(n_T_52[37]), .A4(n497), 
        .Y(N1928) );
  AO22X1_LVT U1267 ( .A1(n1128), .A2(wdata[43]), .A3(n_T_44[37]), .A4(n495), 
        .Y(N1534) );
  AOI22X1_LVT U1268 ( .A1(n1508), .A2(reg_sscratch[44]), .A3(n1162), .A4(n1955), .Y(n825) );
  AO22X1_LVT U1269 ( .A1(n1689), .A2(n_T_45[44]), .A3(n1510), .A4(
        reg_dscratch[44]), .Y(n822) );
  AOI21X1_LVT U1270 ( .A1(n1507), .A2(io_pmp_5_cfg_a[1]), .A3(n822), .Y(n823)
         );
  OR2X1_LVT U1271 ( .A1(n826), .A2(n1690), .Y(io_rw_rdata[44]) );
  AO22X1_LVT U1272 ( .A1(n1149), .A2(wdata[44]), .A3(n_T_52[38]), .A4(n1150), 
        .Y(N1929) );
  AO22X1_LVT U1273 ( .A1(n1128), .A2(wdata[44]), .A3(n_T_44[38]), .A4(n494), 
        .Y(N1535) );
  MUX21X1_LVT U1274 ( .A1(io_pmp_4_addr[9]), .A2(wdata[9]), .S0(n509), .Y(
        n_GEN_286[9]) );
  AO22X1_LVT U1275 ( .A1(n1479), .A2(io_pmp_7_addr[7]), .A3(n1472), .A4(
        io_pmp_5_addr[7]), .Y(n831) );
  AO22X1_LVT U1276 ( .A1(n1491), .A2(io_pmp_4_addr[7]), .A3(n1492), .A4(
        io_pmp_2_addr[7]), .Y(n830) );
  AO22X1_LVT U1277 ( .A1(n1473), .A2(io_pmp_3_addr[7]), .A3(n1494), .A4(
        io_pmp_6_addr[7]), .Y(n829) );
  AO21X1_LVT U1278 ( .A1(n1496), .A2(io_pmp_1_addr[7]), .A3(n827), .Y(n828) );
  NOR4X1_LVT U1279 ( .A1(n831), .A2(n830), .A3(n829), .A4(n828), .Y(n850) );
  AO22X1_LVT U1280 ( .A1(n1153), .A2(n_T_383[7]), .A3(n1474), .A4(
        io_interrupts_mtip), .Y(n835) );
  AO22X1_LVT U1281 ( .A1(n1485), .A2(reg_mscratch[7]), .A3(n1157), .A4(n1932), 
        .Y(n834) );
  AO22X1_LVT U1282 ( .A1(n1160), .A2(n_T_444[7]), .A3(reg_mepc[7]), .A4(n1489), 
        .Y(n833) );
  NOR4X1_LVT U1283 ( .A1(n835), .A2(n834), .A3(n833), .A4(n832), .Y(n849) );
  AO22X1_LVT U1284 ( .A1(n1502), .A2(reg_mie[7]), .A3(n1162), .A4(io_time[7]), 
        .Y(n847) );
  AO22X1_LVT U1285 ( .A1(n1506), .A2(reg_sepc[7]), .A3(reg_stvec[7]), .A4(
        n1478), .Y(n846) );
  NAND2X0_LVT U1286 ( .A1(io_pmp_0_addr[7]), .A2(n1480), .Y(n843) );
  NAND2X0_LVT U1287 ( .A1(io_pmp_0_cfg_l), .A2(n1507), .Y(n839) );
  AOI22X1_LVT U1288 ( .A1(n1493), .A2(reg_dpc[7]), .A3(n1495), .A4(n_T_389[7]), 
        .Y(n838) );
  AOI22X1_LVT U1289 ( .A1(n1689), .A2(n_T_45[7]), .A3(n1510), .A4(
        reg_dscratch[7]), .Y(n837) );
  NAND2X0_LVT U1290 ( .A1(io_ptbr_ppn[7]), .A2(n488), .Y(n836) );
  AND4X1_LVT U1291 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .Y(n842) );
  NAND2X0_LVT U1292 ( .A1(io_bp_0_control_tmatch[0]), .A2(n1481), .Y(n841) );
  NAND2X0_LVT U1293 ( .A1(io_bp_0_address[7]), .A2(n1490), .Y(n840) );
  NAND4X0_LVT U1294 ( .A1(n843), .A2(n842), .A3(n841), .A4(n840), .Y(n845) );
  AND2X1_LVT U1295 ( .A1(n1497), .A2(n659), .Y(n1470) );
  AND2X1_LVT U1296 ( .A1(n1470), .A2(reg_mtvec[7]), .Y(n844) );
  NOR4X1_LVT U1297 ( .A1(n847), .A2(n846), .A3(n845), .A4(n844), .Y(n848) );
  NAND3X0_LVT U1298 ( .A1(n850), .A2(n849), .A3(n848), .Y(io_rw_rdata[7]) );
  AO22X1_LVT U1299 ( .A1(n498), .A2(n_T_52[1]), .A3(wdata[7]), .A4(n1149), .Y(
        N1892) );
  AO22X1_LVT U1300 ( .A1(n1151), .A2(wdata[7]), .A3(io_tval[7]), .A4(n1152), 
        .Y(N1000) );
  AO22X1_LVT U1301 ( .A1(n1158), .A2(wdata[7]), .A3(io_tval[7]), .A4(n1159), 
        .Y(N1389) );
  AO22X1_LVT U1302 ( .A1(reg_mie[7]), .A2(n1503), .A3(wdata[7]), .A4(n1502), 
        .Y(N613) );
  AND2X1_LVT U1303 ( .A1(n1499), .A2(n860), .Y(n1471) );
  AND2X1_LVT U1304 ( .A1(n1467), .A2(n1471), .Y(N469) );
  MUX21X1_LVT U1305 ( .A1(io_pmp_1_addr[7]), .A2(wdata[7]), .S0(n506), .Y(
        n_GEN_265[7]) );
  MUX21X1_LVT U1306 ( .A1(io_pmp_6_addr[7]), .A2(wdata[7]), .S0(n511), .Y(
        n_GEN_300[7]) );
  MUX21X1_LVT U1307 ( .A1(io_pmp_2_addr[7]), .A2(wdata[7]), .S0(n507), .Y(
        n_GEN_272[7]) );
  MUX21X1_LVT U1308 ( .A1(io_pmp_3_addr[7]), .A2(wdata[7]), .S0(n508), .Y(
        n_GEN_279[7]) );
  MUX21X1_LVT U1309 ( .A1(io_pmp_5_addr[7]), .A2(wdata[7]), .S0(n510), .Y(
        n_GEN_293[7]) );
  MUX21X1_LVT U1310 ( .A1(io_pmp_4_addr[7]), .A2(wdata[7]), .S0(n509), .Y(
        n_GEN_286[7]) );
  MUX21X1_LVT U1311 ( .A1(io_pmp_0_addr[7]), .A2(wdata[7]), .S0(n505), .Y(
        n_GEN_258[7]) );
  MUX21X1_LVT U1312 ( .A1(io_pmp_7_addr[7]), .A2(wdata[7]), .S0(n512), .Y(
        n_GEN_307[7]) );
  MUX21X1_LVT U1313 ( .A1(wdata[7]), .A2(wdata[2]), .S0(n1696), .Y(
        n_GEN_155[2]) );
  AO22X1_LVT U1314 ( .A1(n1480), .A2(io_pmp_0_addr[3]), .A3(n1473), .A4(
        io_pmp_3_addr[3]), .Y(n856) );
  AO22X1_LVT U1315 ( .A1(n1472), .A2(io_pmp_5_addr[3]), .A3(n1492), .A4(
        io_pmp_2_addr[3]), .Y(n855) );
  AO22X1_LVT U1316 ( .A1(n1494), .A2(io_pmp_6_addr[3]), .A3(n1496), .A4(
        io_pmp_1_addr[3]), .Y(n854) );
  AO22X1_LVT U1317 ( .A1(n1153), .A2(n_T_383[3]), .A3(n1452), .A4(
        io_status_isa_3_), .Y(n852) );
  AO22X1_LVT U1318 ( .A1(n1161), .A2(reg_mcause[3]), .A3(n1157), .A4(n1934), 
        .Y(n851) );
  OR2X1_LVT U1319 ( .A1(n852), .A2(n851), .Y(n853) );
  NOR4X1_LVT U1320 ( .A1(n856), .A2(n855), .A3(n854), .A4(n853), .Y(n878) );
  AO22X1_LVT U1321 ( .A1(n1474), .A2(io_interrupts_msip), .A3(read_medeleg[3]), 
        .A4(n1469), .Y(n863) );
  AO22X1_LVT U1322 ( .A1(n1485), .A2(reg_mscratch[3]), .A3(reg_mepc[3]), .A4(
        n1489), .Y(n862) );
  AO22X1_LVT U1323 ( .A1(n1160), .A2(n_T_444[3]), .A3(n1168), .A4(
        reg_scause[3]), .Y(n861) );
  AO22X1_LVT U1324 ( .A1(n1508), .A2(reg_sscratch[3]), .A3(reg_sepc[3]), .A4(
        n1506), .Y(n859) );
  NOR4X1_LVT U1325 ( .A1(n863), .A2(n862), .A3(n861), .A4(n859), .Y(n877) );
  AO22X1_LVT U1326 ( .A1(n1502), .A2(reg_mie[3]), .A3(reg_stvec[3]), .A4(n1478), .Y(n864) );
  AOI21X1_LVT U1327 ( .A1(reg_mtvec[3]), .A2(n1470), .A3(n864), .Y(n876) );
  AND2X1_LVT U1328 ( .A1(n1162), .A2(io_time[3]), .Y(n874) );
  NAND2X0_LVT U1329 ( .A1(n1490), .A2(io_bp_0_address[3]), .Y(n870) );
  AOI22X1_LVT U1330 ( .A1(n1493), .A2(reg_dpc[3]), .A3(n488), .A4(
        io_ptbr_ppn[3]), .Y(n869) );
  AOI22X1_LVT U1331 ( .A1(n1689), .A2(n_T_45[3]), .A3(n1510), .A4(
        reg_dscratch[3]), .Y(n865) );
  OA21X1_LVT U1332 ( .A1(n1910), .A2(n866), .A3(n865), .Y(n868) );
  NAND2X0_LVT U1333 ( .A1(n1507), .A2(io_pmp_0_cfg_a[0]), .Y(n867) );
  NAND4X0_LVT U1334 ( .A1(n870), .A2(n869), .A3(n868), .A4(n867), .Y(n873) );
  AO22X1_LVT U1335 ( .A1(n1481), .A2(io_bp_0_control_u), .A3(n1167), .A4(
        read_fcsr[3]), .Y(n872) );
  AO22X1_LVT U1336 ( .A1(n1479), .A2(io_pmp_7_addr[3]), .A3(n1491), .A4(
        io_pmp_4_addr[3]), .Y(n871) );
  NOR4X1_LVT U1337 ( .A1(n874), .A2(n873), .A3(n872), .A4(n871), .Y(n875) );
  NAND4X0_LVT U1338 ( .A1(n878), .A2(n877), .A3(n876), .A4(n875), .Y(
        io_rw_rdata[3]) );
  AND2X1_LVT U1339 ( .A1(n590), .A2(n1910), .Y(n880) );
  MUX21X1_LVT U1340 ( .A1(wdata[3]), .A2(read_fcsr[3]), .S0(n1163), .Y(n881)
         );
  AO21X1_LVT U1341 ( .A1(n1164), .A2(io_fcsr_flags_bits[3]), .A3(n881), .Y(
        n_GEN_345[3]) );
  AO22X1_LVT U1342 ( .A1(n1501), .A2(n1226), .A3(wdata[3]), .A4(n923), .Y(
        N1273) );
  AND2X1_LVT U1343 ( .A1(wdata[3]), .A2(n503), .Y(n1468) );
  AO22X1_LVT U1344 ( .A1(n1498), .A2(n1226), .A3(n1468), .A4(n1161), .Y(N884)
         );
  AO22X1_LVT U1345 ( .A1(wdata[3]), .A2(n1151), .A3(n1152), .A4(io_tval[3]), 
        .Y(N996) );
  AO22X1_LVT U1346 ( .A1(wdata[3]), .A2(n1158), .A3(n1159), .A4(io_tval[3]), 
        .Y(N1385) );
  AO22X1_LVT U1347 ( .A1(reg_mie[3]), .A2(n1503), .A3(wdata[3]), .A4(n1502), 
        .Y(N609) );
  MUX21X1_LVT U1348 ( .A1(io_pc[3]), .A2(wdata[3]), .S0(n513), .Y(net34871) );
  MUX21X1_LVT U1349 ( .A1(io_pmp_6_addr[3]), .A2(wdata[3]), .S0(n511), .Y(
        n_GEN_300[3]) );
  MUX21X1_LVT U1350 ( .A1(io_pmp_2_addr[3]), .A2(wdata[3]), .S0(n507), .Y(
        n_GEN_272[3]) );
  MUX21X1_LVT U1351 ( .A1(io_pmp_3_addr[3]), .A2(wdata[3]), .S0(n508), .Y(
        n_GEN_279[3]) );
  MUX21X1_LVT U1352 ( .A1(io_pmp_5_addr[3]), .A2(wdata[3]), .S0(n510), .Y(
        n_GEN_293[3]) );
  MUX21X1_LVT U1353 ( .A1(io_pmp_4_addr[3]), .A2(wdata[3]), .S0(n509), .Y(
        n_GEN_286[3]) );
  MUX21X1_LVT U1354 ( .A1(io_pmp_0_addr[3]), .A2(wdata[3]), .S0(n505), .Y(
        n_GEN_258[3]) );
  MUX21X1_LVT U1355 ( .A1(io_pmp_7_addr[3]), .A2(wdata[3]), .S0(n512), .Y(
        n_GEN_307[3]) );
  MUX21X1_LVT U1356 ( .A1(io_pc[3]), .A2(wdata[3]), .S0(n514), .Y(net35073) );
  NAND2X0_LVT U1357 ( .A1(n1514), .A2(io_rw_addr[9]), .Y(n882) );
  NAND2X0_LVT U1358 ( .A1(n590), .A2(n1932), .Y(n907) );
  AO21X1_LVT U1359 ( .A1(n503), .A2(n1041), .A3(n883), .Y(n1451) );
  NAND2X0_LVT U1360 ( .A1(n1451), .A2(n1934), .Y(n916) );
  MUX21X1_LVT U1361 ( .A1(read_medeleg[4]), .A2(read_medeleg_6), .S0(n1209), 
        .Y(n884) );
  NAND2X0_LVT U1362 ( .A1(n884), .A2(n954), .Y(n887) );
  MUX21X1_LVT U1363 ( .A1(read_medeleg_13), .A2(read_medeleg_15), .S0(n1209), 
        .Y(n885) );
  NAND2X0_LVT U1364 ( .A1(n885), .A2(io_cause[0]), .Y(n886) );
  MUX21X1_LVT U1365 ( .A1(n887), .A2(n886), .S0(n1226), .Y(n890) );
  AND3X1_LVT U1366 ( .A1(n1226), .A2(n891), .A3(n888), .Y(n896) );
  NAND2X0_LVT U1367 ( .A1(n896), .A2(read_medeleg_12), .Y(n889) );
  NAND2X0_LVT U1368 ( .A1(n890), .A2(n889), .Y(n898) );
  MUX21X1_LVT U1369 ( .A1(read_medeleg_0), .A2(read_medeleg[2]), .S0(n1209), 
        .Y(n893) );
  AND2X1_LVT U1370 ( .A1(read_medeleg[3]), .A2(n1209), .Y(n892) );
  MUX21X1_LVT U1371 ( .A1(n893), .A2(n892), .S0(n1202), .Y(n894) );
  AO22X1_LVT U1372 ( .A1(n896), .A2(read_medeleg_8), .A3(n895), .A4(n894), .Y(
        n897) );
  MUX21X1_LVT U1373 ( .A1(n898), .A2(n897), .S0(n899), .Y(n905) );
  MUX21X1_LVT U1374 ( .A1(read_mideleg_1), .A2(read_mideleg_9_), .S0(n1226), 
        .Y(n900) );
  MUX21X1_LVT U1375 ( .A1(n901), .A2(n900), .S0(n899), .Y(n903) );
  AND3X1_LVT U1376 ( .A1(n903), .A2(n1202), .A3(n902), .Y(n904) );
  OA22X1_LVT U1377 ( .A1(n451), .A2(n907), .A3(n916), .A4(n1255), .Y(n914) );
  INVX1_LVT U1378 ( .A(n1257), .Y(n1198) );
  AND2X1_LVT U1379 ( .A1(n1198), .A2(n1139), .Y(n908) );
  AO21X1_LVT U1380 ( .A1(n1026), .A2(n1903), .A3(n1515), .Y(n910) );
  AND3X1_LVT U1381 ( .A1(n451), .A2(n387), .A3(n501), .Y(n909) );
  AND2X1_LVT U1382 ( .A1(n908), .A2(n1255), .Y(n925) );
  AND2X1_LVT U1383 ( .A1(n909), .A2(n1461), .Y(n930) );
  AO21X1_LVT U1384 ( .A1(n911), .A2(n910), .A3(n930), .Y(n912) );
  NAND3X0_LVT U1385 ( .A1(n912), .A2(n1934), .A3(n590), .Y(n913) );
  AND2X1_LVT U1386 ( .A1(n914), .A2(n913), .Y(n194) );
  MUX21X1_LVT U1387 ( .A1(n1932), .A2(n1934), .S0(n925), .Y(n915) );
  NOR2X0_LVT U1388 ( .A1(n389), .A2(n1041), .Y(n1450) );
  NAND2X0_LVT U1389 ( .A1(n1450), .A2(wdata[7]), .Y(n920) );
  NAND2X0_LVT U1390 ( .A1(n502), .A2(n590), .Y(n919) );
  AO21X1_LVT U1391 ( .A1(n1442), .A2(n917), .A3(n916), .Y(n918) );
  NAND4X0_LVT U1392 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .Y(N360) );
  AO22X1_LVT U1393 ( .A1(n494), .A2(n_T_44[1]), .A3(wdata[7]), .A4(n492), .Y(
        N1498) );
  AO22X1_LVT U1394 ( .A1(n1129), .A2(n_T_44[3]), .A3(wdata[9]), .A4(n492), .Y(
        N1500) );
  MUX21X1_LVT U1395 ( .A1(wdata[4]), .A2(read_fcsr[4]), .S0(n1163), .Y(n922)
         );
  AO21X1_LVT U1396 ( .A1(n1164), .A2(io_fcsr_flags_bits[4]), .A3(n922), .Y(
        n_GEN_345[4]) );
  AO22X1_LVT U1397 ( .A1(n1152), .A2(io_tval[4]), .A3(wdata[4]), .A4(n1151), 
        .Y(N997) );
  AO22X1_LVT U1398 ( .A1(n1159), .A2(io_tval[4]), .A3(wdata[4]), .A4(n1158), 
        .Y(N1386) );
  NAND2X0_LVT U1399 ( .A1(n_T_383[6]), .A2(n1153), .Y(n924) );
  AO22X1_LVT U1400 ( .A1(n498), .A2(n456), .A3(wdata[6]), .A4(n1149), .Y(N1891) );
  AO22X1_LVT U1401 ( .A1(n1152), .A2(io_tval[6]), .A3(wdata[6]), .A4(n1151), 
        .Y(N999) );
  AO22X1_LVT U1402 ( .A1(n1159), .A2(io_tval[6]), .A3(wdata[6]), .A4(n1158), 
        .Y(N1388) );
  MUX21X1_LVT U1403 ( .A1(io_pc[6]), .A2(wdata[6]), .S0(n513), .Y(net34862) );
  AO22X1_LVT U1404 ( .A1(n493), .A2(n455), .A3(wdata[6]), .A4(n492), .Y(N1497)
         );
  NAND2X0_LVT U1405 ( .A1(n1041), .A2(io_exception), .Y(n927) );
  NAND2X0_LVT U1406 ( .A1(n925), .A2(n451), .Y(n926) );
  NAND2X0_LVT U1407 ( .A1(n928), .A2(n501), .Y(n929) );
  NAND2X0_LVT U1408 ( .A1(wdata[11]), .A2(n1450), .Y(n931) );
  MUX21X1_LVT U1409 ( .A1(io_status_prv[0]), .A2(wdata[0]), .S0(n932), .Y(n933) );
  OA22X1_LVT U1410 ( .A1(n_T_389_0), .A2(n935), .A3(n934), .A4(n933), .Y(n2156) );
  OR2X1_LVT U1411 ( .A1(n1257), .A2(n1255), .Y(n1441) );
  AND3X1_LVT U1412 ( .A1(n1139), .A2(n1903), .A3(io_status_debug_BAR), .Y(n952) );
  NAND2X0_LVT U1413 ( .A1(n1441), .A2(n952), .Y(n940) );
  MUX21X1_LVT U1414 ( .A1(n[1930]), .A2(n_T_389_0), .S0(io_rw_addr[10]), .Y(
        n936) );
  AO21X1_LVT U1415 ( .A1(n1199), .A2(n936), .A3(n500), .Y(n951) );
  MUX21X1_LVT U1416 ( .A1(n[1929]), .A2(n_T_389_1), .S0(io_rw_addr[10]), .Y(
        n937) );
  NAND3X0_LVT U1417 ( .A1(n951), .A2(io_rw_addr[9]), .A3(n937), .Y(n939) );
  AND2X1_LVT U1418 ( .A1(io_status_prv[0]), .A2(n1903), .Y(n950) );
  NAND2X0_LVT U1419 ( .A1(n950), .A2(io_status_prv[1]), .Y(n938) );
  AND2X1_LVT U1420 ( .A1(n1499), .A2(n941), .Y(n946) );
  AO21X1_LVT U1421 ( .A1(n1257), .A2(n1139), .A3(n1356), .Y(n945) );
  INVX1_LVT U1422 ( .A(n942), .Y(n943) );
  MUX21X1_LVT U1423 ( .A1(io_status_debug), .A2(n943), .S0(n945), .Y(n944) );
  AO22X1_LVT U1424 ( .A1(n946), .A2(n945), .A3(n944), .A4(n590), .Y(n2161) );
  NAND2X0_LVT U1425 ( .A1(n1490), .A2(io_bp_0_address[8]), .Y(n948) );
  NAND2X0_LVT U1426 ( .A1(n1495), .A2(n_T_389[8]), .Y(n947) );
  AO22X1_LVT U1427 ( .A1(n1498), .A2(n1202), .A3(wdata[0]), .A4(n955), .Y(N881) );
  AO22X1_LVT U1428 ( .A1(io_tval[0]), .A2(n1152), .A3(wdata[0]), .A4(n1151), 
        .Y(N993) );
  AO22X1_LVT U1429 ( .A1(io_tval[0]), .A2(n1159), .A3(wdata[0]), .A4(n1158), 
        .Y(N1382) );
  OAI22X1_LVT U1430 ( .A1(n959), .A2(n958), .A3(n957), .A4(n1483), .Y(N1430)
         );
  AO22X1_LVT U1431 ( .A1(n1128), .A2(wdata[63]), .A3(n_T_44[57]), .A4(n1129), 
        .Y(N1554) );
  AOI22X1_LVT U1432 ( .A1(n1508), .A2(reg_sscratch[62]), .A3(n1162), .A4(n1937), .Y(n964) );
  AOI22X1_LVT U1433 ( .A1(n1689), .A2(n_T_45[62]), .A3(n1510), .A4(
        reg_dscratch[62]), .Y(n962) );
  OR2X1_LVT U1434 ( .A1(n965), .A2(n1690), .Y(io_rw_rdata[62]) );
  AO22X1_LVT U1435 ( .A1(n1149), .A2(wdata[62]), .A3(n_T_52[56]), .A4(n1150), 
        .Y(N1947) );
  AO22X1_LVT U1436 ( .A1(n1128), .A2(wdata[62]), .A3(n_T_44[56]), .A4(n494), 
        .Y(N1553) );
  AOI22X1_LVT U1437 ( .A1(n1508), .A2(reg_sscratch[61]), .A3(n1162), .A4(n1938), .Y(n967) );
  NAND4X0_LVT U1438 ( .A1(n968), .A2(n967), .A3(n467), .A4(n966), .Y(
        io_rw_rdata[61]) );
  AO22X1_LVT U1439 ( .A1(n1149), .A2(wdata[61]), .A3(n_T_52[55]), .A4(n1150), 
        .Y(N1946) );
  AO22X1_LVT U1440 ( .A1(n1128), .A2(wdata[61]), .A3(n_T_44[55]), .A4(n1129), 
        .Y(N1552) );
  AO22X1_LVT U1441 ( .A1(n1689), .A2(n_T_45[58]), .A3(n1510), .A4(
        reg_dscratch[58]), .Y(n969) );
  NAND4X0_LVT U1442 ( .A1(n481), .A2(n1688), .A3(n474), .A4(n970), .Y(
        io_rw_rdata[58]) );
  AO22X1_LVT U1443 ( .A1(n1689), .A2(n_T_45[57]), .A3(n1510), .A4(
        reg_dscratch[57]), .Y(n971) );
  NAND4X0_LVT U1444 ( .A1(n481), .A2(n1687), .A3(n475), .A4(n972), .Y(
        io_rw_rdata[57]) );
  AO22X1_LVT U1445 ( .A1(n1149), .A2(wdata[57]), .A3(n_T_52[51]), .A4(n497), 
        .Y(N1942) );
  AOI22X1_LVT U1446 ( .A1(n1689), .A2(n_T_45[56]), .A3(n1510), .A4(
        reg_dscratch[56]), .Y(n974) );
  NAND2X0_LVT U1447 ( .A1(n1162), .A2(n1943), .Y(n973) );
  NAND3X0_LVT U1448 ( .A1(n481), .A2(n1686), .A3(n976), .Y(io_rw_rdata[56]) );
  AO22X1_LVT U1449 ( .A1(n1149), .A2(wdata[56]), .A3(n_T_52[50]), .A4(n497), 
        .Y(N1941) );
  AO22X1_LVT U1450 ( .A1(n1128), .A2(wdata[56]), .A3(n_T_44[50]), .A4(n494), 
        .Y(N1547) );
  AO22X1_LVT U1451 ( .A1(n1128), .A2(wdata[57]), .A3(n_T_44[51]), .A4(n495), 
        .Y(N1548) );
  AOI22X1_LVT U1452 ( .A1(n1508), .A2(reg_sscratch[54]), .A3(n1162), .A4(n1945), .Y(n979) );
  AOI22X1_LVT U1453 ( .A1(n1689), .A2(n_T_45[54]), .A3(n1510), .A4(
        reg_dscratch[54]), .Y(n977) );
  OR2X1_LVT U1454 ( .A1(n980), .A2(n1690), .Y(io_rw_rdata[54]) );
  AO22X1_LVT U1455 ( .A1(n1128), .A2(wdata[54]), .A3(n_T_44[48]), .A4(n494), 
        .Y(N1545) );
  AOI22X1_LVT U1456 ( .A1(n1508), .A2(reg_sscratch[53]), .A3(n1162), .A4(n1946), .Y(n983) );
  AOI22X1_LVT U1457 ( .A1(n1689), .A2(n_T_45[53]), .A3(n1510), .A4(
        reg_dscratch[53]), .Y(n981) );
  OR2X1_LVT U1458 ( .A1(n984), .A2(n1690), .Y(io_rw_rdata[53]) );
  AO22X1_LVT U1459 ( .A1(n1149), .A2(wdata[53]), .A3(n_T_52[47]), .A4(n497), 
        .Y(N1938) );
  AO22X1_LVT U1460 ( .A1(n1128), .A2(wdata[53]), .A3(n_T_44[47]), .A4(n1129), 
        .Y(N1544) );
  AOI22X1_LVT U1461 ( .A1(n1689), .A2(n_T_45[50]), .A3(n1510), .A4(
        reg_dscratch[50]), .Y(n986) );
  NAND2X0_LVT U1462 ( .A1(n1162), .A2(n1949), .Y(n985) );
  NAND3X0_LVT U1463 ( .A1(n481), .A2(n1683), .A3(n988), .Y(io_rw_rdata[50]) );
  AOI22X1_LVT U1464 ( .A1(n1689), .A2(n_T_45[49]), .A3(n1507), .A4(
        io_pmp_6_cfg_w), .Y(n990) );
  NAND2X0_LVT U1465 ( .A1(n1162), .A2(n1950), .Y(n989) );
  NAND3X0_LVT U1466 ( .A1(n481), .A2(n1682), .A3(n992), .Y(io_rw_rdata[49]) );
  AO22X1_LVT U1467 ( .A1(n1149), .A2(wdata[49]), .A3(n_T_52[43]), .A4(n496), 
        .Y(N1934) );
  AOI22X1_LVT U1468 ( .A1(n1689), .A2(n_T_45[48]), .A3(n1507), .A4(
        io_pmp_6_cfg_r), .Y(n994) );
  NAND2X0_LVT U1469 ( .A1(n1162), .A2(n1951), .Y(n993) );
  NAND3X0_LVT U1470 ( .A1(n481), .A2(n1681), .A3(n996), .Y(io_rw_rdata[48]) );
  AO22X1_LVT U1471 ( .A1(n1149), .A2(wdata[48]), .A3(n_T_52[42]), .A4(n497), 
        .Y(N1933) );
  AO22X1_LVT U1472 ( .A1(n1128), .A2(wdata[48]), .A3(n_T_44[42]), .A4(n1129), 
        .Y(N1539) );
  AO22X1_LVT U1473 ( .A1(n1128), .A2(wdata[49]), .A3(n_T_44[43]), .A4(n495), 
        .Y(N1540) );
  AO22X1_LVT U1474 ( .A1(n1485), .A2(reg_mscratch[46]), .A3(n1162), .A4(n1953), 
        .Y(n997) );
  OR3X1_LVT U1475 ( .A1(n998), .A2(n997), .A3(n1679), .Y(io_rw_rdata[46]) );
  AO22X1_LVT U1476 ( .A1(n_T_52[40]), .A2(n1150), .A3(n1149), .A4(wdata[46]), 
        .Y(N1931) );
  AO22X1_LVT U1477 ( .A1(n_T_44[40]), .A2(n1129), .A3(n492), .A4(wdata[46]), 
        .Y(N1537) );
  AOI22X1_LVT U1478 ( .A1(n1508), .A2(reg_sscratch[45]), .A3(n1162), .A4(n1954), .Y(n1001) );
  AOI22X1_LVT U1479 ( .A1(n1689), .A2(n_T_45[45]), .A3(n1510), .A4(
        reg_dscratch[45]), .Y(n999) );
  OR2X1_LVT U1480 ( .A1(n1002), .A2(n1690), .Y(io_rw_rdata[45]) );
  AO22X1_LVT U1481 ( .A1(n1149), .A2(wdata[45]), .A3(n_T_52[39]), .A4(n496), 
        .Y(N1930) );
  AO22X1_LVT U1482 ( .A1(n1128), .A2(wdata[45]), .A3(n_T_44[39]), .A4(n495), 
        .Y(N1536) );
  AOI22X1_LVT U1483 ( .A1(n1689), .A2(n_T_45[42]), .A3(n1507), .A4(
        io_pmp_5_cfg_x), .Y(n1004) );
  NAND2X0_LVT U1484 ( .A1(n1162), .A2(n1957), .Y(n1003) );
  NAND3X0_LVT U1485 ( .A1(n481), .A2(n1677), .A3(n1006), .Y(io_rw_rdata[42])
         );
  AO22X1_LVT U1486 ( .A1(n1149), .A2(wdata[42]), .A3(n_T_52[36]), .A4(n497), 
        .Y(N1927) );
  AO22X1_LVT U1487 ( .A1(n1128), .A2(wdata[42]), .A3(n_T_44[36]), .A4(n495), 
        .Y(N1533) );
  AO22X1_LVT U1488 ( .A1(n1508), .A2(reg_sscratch[41]), .A3(n1162), .A4(n1958), 
        .Y(n1007) );
  NOR3X0_LVT U1489 ( .A1(n1009), .A2(n1008), .A3(n1007), .Y(n1010) );
  NAND3X0_LVT U1490 ( .A1(n481), .A2(n1676), .A3(n1010), .Y(io_rw_rdata[41])
         );
  AO22X1_LVT U1491 ( .A1(n1149), .A2(wdata[41]), .A3(n_T_52[35]), .A4(n496), 
        .Y(N1926) );
  AO22X1_LVT U1492 ( .A1(n1128), .A2(wdata[41]), .A3(n_T_44[35]), .A4(n494), 
        .Y(N1532) );
  AOI22X1_LVT U1493 ( .A1(n1689), .A2(n_T_45[40]), .A3(n1510), .A4(
        reg_dscratch[40]), .Y(n1012) );
  NAND2X0_LVT U1494 ( .A1(n1162), .A2(n1959), .Y(n1011) );
  NAND3X0_LVT U1495 ( .A1(n481), .A2(n1675), .A3(n1014), .Y(io_rw_rdata[40])
         );
  AO22X1_LVT U1496 ( .A1(n1149), .A2(wdata[40]), .A3(n_T_52[34]), .A4(n496), 
        .Y(N1925) );
  AO22X1_LVT U1497 ( .A1(n1128), .A2(wdata[40]), .A3(n_T_44[34]), .A4(n495), 
        .Y(N1531) );
  AO22X1_LVT U1498 ( .A1(wdata[38]), .A2(n1151), .A3(n1152), .A4(io_tval[38]), 
        .Y(N1031) );
  AO22X1_LVT U1499 ( .A1(wdata[38]), .A2(n1158), .A3(n1159), .A4(io_tval[38]), 
        .Y(N1420) );
  MUX21X1_LVT U1500 ( .A1(io_pc[38]), .A2(wdata[38]), .S0(n513), .Y(net34766)
         );
  MUX21X1_LVT U1501 ( .A1(io_pc[38]), .A2(wdata[38]), .S0(n515), .Y(net35190)
         );
  MUX21X1_LVT U1502 ( .A1(io_pc[38]), .A2(wdata[38]), .S0(n514), .Y(net34968)
         );
  AOI22X1_LVT U1503 ( .A1(n1160), .A2(n_T_444[37]), .A3(n1508), .A4(
        reg_sscratch[37]), .Y(n1018) );
  AOI22X1_LVT U1504 ( .A1(n1689), .A2(n_T_45[37]), .A3(n1487), .A4(
        reg_stvec[37]), .Y(n1017) );
  NAND2X0_LVT U1505 ( .A1(n1153), .A2(n_T_383[37]), .Y(n1016) );
  NAND2X0_LVT U1506 ( .A1(n1162), .A2(n1962), .Y(n1015) );
  NAND4X0_LVT U1507 ( .A1(n1018), .A2(n1017), .A3(n1016), .A4(n1015), .Y(n1019) );
  OR2X1_LVT U1508 ( .A1(n1019), .A2(n1648), .Y(io_rw_rdata[37]) );
  AO22X1_LVT U1509 ( .A1(n498), .A2(n_T_52[31]), .A3(wdata[37]), .A4(n1149), 
        .Y(N1922) );
  AO22X1_LVT U1510 ( .A1(n1152), .A2(io_tval[37]), .A3(wdata[37]), .A4(n1151), 
        .Y(N1030) );
  AO22X1_LVT U1511 ( .A1(n1159), .A2(io_tval[37]), .A3(wdata[37]), .A4(n1158), 
        .Y(N1419) );
  AO22X1_LVT U1512 ( .A1(n495), .A2(n_T_44[31]), .A3(wdata[37]), .A4(n491), 
        .Y(N1528) );
  AO22X1_LVT U1513 ( .A1(n_T_44[30]), .A2(n495), .A3(wdata[36]), .A4(n491), 
        .Y(N1527) );
  AO22X1_LVT U1514 ( .A1(n1160), .A2(n_T_444[34]), .A3(n1508), .A4(
        reg_sscratch[34]), .Y(n1025) );
  NAND2X0_LVT U1515 ( .A1(n1506), .A2(reg_sepc[34]), .Y(n1023) );
  NAND2X0_LVT U1516 ( .A1(n1153), .A2(n_T_383[34]), .Y(n1022) );
  AOI22X1_LVT U1517 ( .A1(n1689), .A2(n_T_45[34]), .A3(n1510), .A4(
        reg_dscratch[34]), .Y(n1021) );
  NAND2X0_LVT U1518 ( .A1(n1490), .A2(io_bp_0_address[34]), .Y(n1020) );
  NAND4X0_LVT U1519 ( .A1(n1023), .A2(n1022), .A3(n1021), .A4(n1020), .Y(n1024) );
  OR3X1_LVT U1520 ( .A1(n1025), .A2(n1024), .A3(n1638), .Y(io_rw_rdata[34]) );
  AO22X1_LVT U1521 ( .A1(n1152), .A2(io_tval[34]), .A3(wdata[34]), .A4(n1151), 
        .Y(N1027) );
  AO22X1_LVT U1522 ( .A1(n1159), .A2(io_tval[34]), .A3(wdata[34]), .A4(n1158), 
        .Y(N1416) );
  MUX21X1_LVT U1523 ( .A1(io_pc[34]), .A2(wdata[34]), .S0(n513), .Y(net34778)
         );
  AO22X1_LVT U1524 ( .A1(n1129), .A2(n_T_44[28]), .A3(wdata[34]), .A4(n491), 
        .Y(N1525) );
  AO22X1_LVT U1525 ( .A1(n1149), .A2(wdata[33]), .A3(n_T_52[27]), .A4(n496), 
        .Y(N1918) );
  AO22X1_LVT U1526 ( .A1(n1151), .A2(wdata[33]), .A3(io_tval[33]), .A4(n1152), 
        .Y(N1026) );
  AO22X1_LVT U1527 ( .A1(n1158), .A2(wdata[33]), .A3(io_tval[33]), .A4(n1159), 
        .Y(N1415) );
  MUX21X1_LVT U1528 ( .A1(io_pc[33]), .A2(wdata[33]), .S0(n513), .Y(net34781)
         );
  MUX21X1_LVT U1529 ( .A1(io_pc[33]), .A2(wdata[33]), .S0(n515), .Y(net35205)
         );
  MUX21X1_LVT U1530 ( .A1(io_pc[33]), .A2(wdata[33]), .S0(n514), .Y(net34983)
         );
  AO22X1_LVT U1531 ( .A1(n1128), .A2(wdata[33]), .A3(n_T_44[27]), .A4(n495), 
        .Y(N1524) );
  AO22X1_LVT U1532 ( .A1(n1160), .A2(n_T_444[32]), .A3(n1485), .A4(
        reg_mscratch[32]), .Y(n1032) );
  NAND2X0_LVT U1533 ( .A1(n1506), .A2(reg_sepc[32]), .Y(n1030) );
  NAND2X0_LVT U1534 ( .A1(n1153), .A2(n_T_383[32]), .Y(n1029) );
  AOI22X1_LVT U1535 ( .A1(n1689), .A2(n_T_45[32]), .A3(n1493), .A4(reg_dpc[32]), .Y(n1028) );
  NAND2X0_LVT U1536 ( .A1(n1490), .A2(io_bp_0_address[32]), .Y(n1027) );
  NAND4X0_LVT U1537 ( .A1(n1030), .A2(n1029), .A3(n1028), .A4(n1027), .Y(n1031) );
  OR3X1_LVT U1538 ( .A1(n1032), .A2(n1031), .A3(n1633), .Y(io_rw_rdata[32]) );
  AO22X1_LVT U1539 ( .A1(n1152), .A2(io_tval[32]), .A3(wdata[32]), .A4(n1151), 
        .Y(N1025) );
  AO22X1_LVT U1540 ( .A1(n1159), .A2(io_tval[32]), .A3(wdata[32]), .A4(n1158), 
        .Y(N1414) );
  MUX21X1_LVT U1541 ( .A1(io_pc[32]), .A2(wdata[32]), .S0(n513), .Y(net34784)
         );
  MUX21X1_LVT U1542 ( .A1(io_pc[32]), .A2(wdata[32]), .S0(n515), .Y(net35208)
         );
  AO22X1_LVT U1543 ( .A1(n495), .A2(n_T_44[26]), .A3(wdata[32]), .A4(n491), 
        .Y(N1523) );
  AOI22X1_LVT U1544 ( .A1(n1160), .A2(n_T_444[30]), .A3(n1506), .A4(
        reg_sepc[30]), .Y(n1042) );
  NAND2X0_LVT U1545 ( .A1(n1490), .A2(io_bp_0_address[30]), .Y(n1036) );
  AOI21X1_LVT U1546 ( .A1(n_T_45[30]), .A2(n1689), .A3(n1627), .Y(n1035) );
  NAND2X0_LVT U1547 ( .A1(n1493), .A2(reg_dpc[30]), .Y(n1034) );
  NAND2X0_LVT U1548 ( .A1(n1510), .A2(reg_dscratch[30]), .Y(n1033) );
  NAND4X0_LVT U1549 ( .A1(n1036), .A2(n1035), .A3(n1034), .A4(n1033), .Y(n1037) );
  AOI21X1_LVT U1550 ( .A1(n1153), .A2(n_T_383[30]), .A3(n1037), .Y(n1039) );
  NAND2X0_LVT U1551 ( .A1(n1162), .A2(io_time[30]), .Y(n1038) );
  NAND4X0_LVT U1552 ( .A1(n1042), .A2(n1040), .A3(n1039), .A4(n1038), .Y(n1043) );
  OR2X1_LVT U1553 ( .A1(n1043), .A2(n1628), .Y(io_rw_rdata[30]) );
  AO22X1_LVT U1554 ( .A1(n498), .A2(n_T_52[24]), .A3(wdata[30]), .A4(n1149), 
        .Y(N1915) );
  AO22X1_LVT U1555 ( .A1(wdata[30]), .A2(n1151), .A3(n1152), .A4(io_tval[30]), 
        .Y(N1023) );
  AO22X1_LVT U1556 ( .A1(wdata[30]), .A2(n1158), .A3(n1159), .A4(io_tval[30]), 
        .Y(N1412) );
  MUX21X1_LVT U1557 ( .A1(io_pc[30]), .A2(wdata[30]), .S0(n513), .Y(net34790)
         );
  MUX21X1_LVT U1558 ( .A1(io_pc[30]), .A2(wdata[30]), .S0(n515), .Y(net35214)
         );
  AO22X1_LVT U1559 ( .A1(n494), .A2(n_T_44[24]), .A3(wdata[30]), .A4(n491), 
        .Y(N1521) );
  AO22X1_LVT U1560 ( .A1(n1162), .A2(io_time[29]), .A3(n1480), .A4(
        io_pmp_0_addr[29]), .Y(n1044) );
  OR3X1_LVT U1561 ( .A1(n1045), .A2(n1044), .A3(n1625), .Y(n1046) );
  NOR3X0_LVT U1562 ( .A1(n1622), .A2(n1620), .A3(n1046), .Y(n1053) );
  AO22X1_LVT U1563 ( .A1(n1689), .A2(n_T_45[29]), .A3(n1493), .A4(reg_dpc[29]), 
        .Y(n1047) );
  AO21X1_LVT U1564 ( .A1(n1487), .A2(reg_stvec[29]), .A3(n1047), .Y(n1048) );
  AO21X1_LVT U1565 ( .A1(n1153), .A2(n_T_383[29]), .A3(n1048), .Y(n1050) );
  NOR4X1_LVT U1566 ( .A1(n1626), .A2(n1050), .A3(n1049), .A4(n1623), .Y(n1051)
         );
  NAND3X0_LVT U1567 ( .A1(n1053), .A2(n1052), .A3(n1051), .Y(io_rw_rdata[29])
         );
  AO22X1_LVT U1568 ( .A1(n496), .A2(n_T_52[23]), .A3(wdata[29]), .A4(n1149), 
        .Y(N1914) );
  AO22X1_LVT U1569 ( .A1(n1152), .A2(io_tval[29]), .A3(wdata[29]), .A4(n1151), 
        .Y(N1022) );
  AO22X1_LVT U1570 ( .A1(n1159), .A2(io_tval[29]), .A3(wdata[29]), .A4(n1158), 
        .Y(N1411) );
  MUX21X1_LVT U1571 ( .A1(io_pc[29]), .A2(wdata[29]), .S0(n515), .Y(net35217)
         );
  MUX21X1_LVT U1572 ( .A1(io_pc[29]), .A2(wdata[29]), .S0(n514), .Y(net34995)
         );
  AO22X1_LVT U1573 ( .A1(n494), .A2(n_T_44[23]), .A3(wdata[29]), .A4(n491), 
        .Y(N1520) );
  AO22X1_LVT U1574 ( .A1(n498), .A2(n_T_52[20]), .A3(wdata[26]), .A4(n1149), 
        .Y(N1911) );
  AO22X1_LVT U1575 ( .A1(n1152), .A2(io_tval[26]), .A3(wdata[26]), .A4(n1151), 
        .Y(N1019) );
  AO22X1_LVT U1576 ( .A1(n1159), .A2(io_tval[26]), .A3(wdata[26]), .A4(n1158), 
        .Y(N1408) );
  MUX21X1_LVT U1577 ( .A1(io_pc[26]), .A2(wdata[26]), .S0(n514), .Y(net35004)
         );
  AO22X1_LVT U1578 ( .A1(n1129), .A2(n_T_44[20]), .A3(wdata[26]), .A4(n491), 
        .Y(N1517) );
  AO22X1_LVT U1579 ( .A1(n497), .A2(n_T_52[19]), .A3(wdata[25]), .A4(n1149), 
        .Y(N1910) );
  AO22X1_LVT U1580 ( .A1(n1152), .A2(io_tval[25]), .A3(wdata[25]), .A4(n1151), 
        .Y(N1018) );
  AO22X1_LVT U1581 ( .A1(n1159), .A2(io_tval[25]), .A3(wdata[25]), .A4(n1158), 
        .Y(N1407) );
  MUX21X1_LVT U1582 ( .A1(io_pc[25]), .A2(wdata[25]), .S0(n513), .Y(net34805)
         );
  AO22X1_LVT U1583 ( .A1(n494), .A2(n_T_44[19]), .A3(wdata[25]), .A4(n491), 
        .Y(N1516) );
  NAND2X0_LVT U1584 ( .A1(n1153), .A2(n_T_383[24]), .Y(n1057) );
  AOI22X1_LVT U1585 ( .A1(n1689), .A2(n_T_45[24]), .A3(n1493), .A4(reg_dpc[24]), .Y(n1056) );
  NAND2X0_LVT U1586 ( .A1(n1487), .A2(reg_stvec[24]), .Y(n1055) );
  NAND2X0_LVT U1587 ( .A1(n1507), .A2(io_pmp_3_cfg_r), .Y(n1054) );
  AND4X1_LVT U1588 ( .A1(n1057), .A2(n1056), .A3(n1055), .A4(n1054), .Y(n1059)
         );
  NAND2X0_LVT U1589 ( .A1(n1162), .A2(io_time[24]), .Y(n1058) );
  NAND4X0_LVT U1590 ( .A1(n1061), .A2(n1060), .A3(n1059), .A4(n1058), .Y(n1063) );
  NOR4X1_LVT U1591 ( .A1(n1612), .A2(n1063), .A3(n1606), .A4(n1607), .Y(n1064)
         );
  NAND2X0_LVT U1592 ( .A1(n1613), .A2(n1064), .Y(io_rw_rdata[24]) );
  AO22X1_LVT U1593 ( .A1(n496), .A2(n_T_52[18]), .A3(wdata[24]), .A4(n1149), 
        .Y(N1909) );
  AO22X1_LVT U1594 ( .A1(n1152), .A2(io_tval[24]), .A3(wdata[24]), .A4(n1151), 
        .Y(N1017) );
  AO22X1_LVT U1595 ( .A1(n1159), .A2(io_tval[24]), .A3(wdata[24]), .A4(n1158), 
        .Y(N1406) );
  MUX21X1_LVT U1596 ( .A1(io_pc[24]), .A2(wdata[24]), .S0(n515), .Y(net35232)
         );
  AO22X1_LVT U1597 ( .A1(n493), .A2(n_T_44[18]), .A3(wdata[24]), .A4(n491), 
        .Y(N1515) );
  AO22X1_LVT U1598 ( .A1(n498), .A2(n_T_52[16]), .A3(wdata[22]), .A4(n1149), 
        .Y(N1907) );
  AO22X1_LVT U1599 ( .A1(n1152), .A2(io_tval[22]), .A3(wdata[22]), .A4(n1151), 
        .Y(N1015) );
  AO22X1_LVT U1600 ( .A1(n1159), .A2(io_tval[22]), .A3(wdata[22]), .A4(n1158), 
        .Y(N1404) );
  MUX21X1_LVT U1601 ( .A1(io_pc[22]), .A2(wdata[22]), .S0(n515), .Y(net35238)
         );
  AO22X1_LVT U1602 ( .A1(n493), .A2(n_T_44[16]), .A3(wdata[22]), .A4(n491), 
        .Y(N1513) );
  AO22X1_LVT U1603 ( .A1(n497), .A2(n_T_52[15]), .A3(wdata[21]), .A4(n1149), 
        .Y(N1906) );
  AO22X1_LVT U1604 ( .A1(n1152), .A2(io_tval[21]), .A3(wdata[21]), .A4(n1151), 
        .Y(N1014) );
  AO22X1_LVT U1605 ( .A1(n1159), .A2(io_tval[21]), .A3(wdata[21]), .A4(n1158), 
        .Y(N1403) );
  MUX21X1_LVT U1606 ( .A1(io_pc[21]), .A2(wdata[21]), .S0(n514), .Y(net35019)
         );
  AO22X1_LVT U1607 ( .A1(n493), .A2(n_T_44[15]), .A3(wdata[21]), .A4(n1128), 
        .Y(N1512) );
  AOI22X1_LVT U1608 ( .A1(n1162), .A2(io_time[20]), .A3(n1506), .A4(
        reg_sepc[20]), .Y(n1071) );
  NAND2X0_LVT U1609 ( .A1(io_pmp_2_cfg_a[1]), .A2(n1507), .Y(n1067) );
  NAND2X0_LVT U1610 ( .A1(n1493), .A2(reg_dpc[20]), .Y(n1066) );
  NAND2X0_LVT U1611 ( .A1(n1510), .A2(reg_dscratch[20]), .Y(n1065) );
  AND4X1_LVT U1612 ( .A1(n1067), .A2(n1083), .A3(n1066), .A4(n1065), .Y(n1070)
         );
  NAND2X0_LVT U1613 ( .A1(n1920), .A2(n1452), .Y(n1069) );
  NAND2X0_LVT U1614 ( .A1(io_pmp_2_addr[20]), .A2(n1492), .Y(n1068) );
  NAND4X0_LVT U1615 ( .A1(n1071), .A2(n1070), .A3(n1069), .A4(n1068), .Y(n1077) );
  AOI22X1_LVT U1616 ( .A1(n1485), .A2(reg_mscratch[20]), .A3(n1157), .A4(n1926), .Y(n1075) );
  AOI22X1_LVT U1617 ( .A1(n1160), .A2(n_T_444[20]), .A3(n1489), .A4(
        reg_mepc[20]), .Y(n1074) );
  NAND4X0_LVT U1618 ( .A1(n1075), .A2(n1074), .A3(n1073), .A4(n1072), .Y(n1076) );
  NOR4X1_LVT U1619 ( .A1(n1077), .A2(n1076), .A3(n1592), .A4(n1595), .Y(n1079)
         );
  NOR3X0_LVT U1620 ( .A1(n1594), .A2(n1597), .A3(n1593), .Y(n1078) );
  NAND2X0_LVT U1621 ( .A1(n1079), .A2(n1078), .Y(io_rw_rdata[20]) );
  AO22X1_LVT U1622 ( .A1(n496), .A2(n_T_52[14]), .A3(wdata[20]), .A4(n1149), 
        .Y(N1905) );
  AO22X1_LVT U1623 ( .A1(n1152), .A2(io_tval[20]), .A3(wdata[20]), .A4(n1151), 
        .Y(N1013) );
  AO22X1_LVT U1624 ( .A1(n1159), .A2(io_tval[20]), .A3(wdata[20]), .A4(n1158), 
        .Y(N1402) );
  AO21X1_LVT U1625 ( .A1(n1920), .A2(n504), .A3(n376), .Y(N1579) );
  MUX21X1_LVT U1626 ( .A1(io_pc[20]), .A2(wdata[20]), .S0(n513), .Y(net34820)
         );
  MUX21X1_LVT U1627 ( .A1(io_pc[20]), .A2(wdata[20]), .S0(n515), .Y(net35244)
         );
  MUX21X1_LVT U1628 ( .A1(io_pc[20]), .A2(wdata[20]), .S0(n514), .Y(net35022)
         );
  AO22X1_LVT U1629 ( .A1(n493), .A2(n_T_44[14]), .A3(wdata[20]), .A4(n491), 
        .Y(N1511) );
  AO22X1_LVT U1630 ( .A1(n1160), .A2(n_T_444[19]), .A3(n1497), .A4(
        reg_mtvec[19]), .Y(n1080) );
  NOR4X1_LVT U1631 ( .A1(n1587), .A2(n1081), .A3(n1080), .A4(n1588), .Y(n1095)
         );
  AO22X1_LVT U1632 ( .A1(n1479), .A2(io_pmp_7_addr[19]), .A3(n1480), .A4(
        io_pmp_0_addr[19]), .Y(n1091) );
  AO22X1_LVT U1633 ( .A1(n1472), .A2(io_pmp_5_addr[19]), .A3(n1492), .A4(
        io_pmp_2_addr[19]), .Y(n1090) );
  NAND2X0_LVT U1634 ( .A1(io_pmp_6_addr[19]), .A2(n1494), .Y(n1088) );
  NAND2X0_LVT U1635 ( .A1(io_pmp_2_cfg_a[0]), .A2(n1507), .Y(n1084) );
  NAND2X0_LVT U1636 ( .A1(n488), .A2(io_ptbr_ppn[19]), .Y(n1082) );
  AND4X1_LVT U1637 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n478), .Y(n1087)
         );
  NAND2X0_LVT U1638 ( .A1(n_T_383[19]), .A2(n1153), .Y(n1086) );
  NAND2X0_LVT U1639 ( .A1(io_status_mxr), .A2(n1154), .Y(n1085) );
  NAND4X0_LVT U1640 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .Y(n1089) );
  NOR4X1_LVT U1641 ( .A1(n1092), .A2(n1091), .A3(n1090), .A4(n1089), .Y(n1093)
         );
  NAND3X0_LVT U1642 ( .A1(n1095), .A2(n1094), .A3(n1093), .Y(io_rw_rdata[19])
         );
  AO22X1_LVT U1643 ( .A1(n498), .A2(n_T_52[13]), .A3(wdata[19]), .A4(n1149), 
        .Y(N1904) );
  AO22X1_LVT U1644 ( .A1(n1152), .A2(io_tval[19]), .A3(wdata[19]), .A4(n1151), 
        .Y(N1012) );
  AO22X1_LVT U1645 ( .A1(n1159), .A2(io_tval[19]), .A3(wdata[19]), .A4(n1158), 
        .Y(N1401) );
  AO22X1_LVT U1646 ( .A1(n493), .A2(n_T_44[13]), .A3(wdata[19]), .A4(n1128), 
        .Y(N1510) );
  AO22X1_LVT U1647 ( .A1(n1491), .A2(io_pmp_4_addr[18]), .A3(n1496), .A4(
        io_pmp_1_addr[18]), .Y(n1102) );
  NAND2X0_LVT U1648 ( .A1(reg_stvec[18]), .A2(n1487), .Y(n1099) );
  NAND2X0_LVT U1649 ( .A1(io_status_sum), .A2(n1154), .Y(n1098) );
  AOI22X1_LVT U1650 ( .A1(n1689), .A2(n_T_45[18]), .A3(n1510), .A4(
        reg_dscratch[18]), .Y(n1097) );
  NAND2X0_LVT U1651 ( .A1(io_pmp_2_cfg_x), .A2(n1507), .Y(n1096) );
  NAND4X0_LVT U1652 ( .A1(n1099), .A2(n1098), .A3(n1097), .A4(n1096), .Y(n1101) );
  AO22X1_LVT U1653 ( .A1(n1153), .A2(n_T_383[18]), .A3(n1452), .A4(n1921), .Y(
        n1100) );
  NOR4X1_LVT U1654 ( .A1(n1102), .A2(n1101), .A3(n1100), .A4(n1582), .Y(n1110)
         );
  AO22X1_LVT U1655 ( .A1(n1162), .A2(io_time[18]), .A3(n1480), .A4(
        io_pmp_0_addr[18]), .Y(n1104) );
  AO22X1_LVT U1656 ( .A1(n1479), .A2(io_pmp_7_addr[18]), .A3(n1473), .A4(
        io_pmp_3_addr[18]), .Y(n1103) );
  NOR4X1_LVT U1657 ( .A1(n1106), .A2(n1105), .A3(n1104), .A4(n1103), .Y(n1108)
         );
  NAND4X0_LVT U1658 ( .A1(n1110), .A2(n1109), .A3(n1108), .A4(n1107), .Y(
        io_rw_rdata[18]) );
  AO22X1_LVT U1659 ( .A1(n498), .A2(n_T_52[12]), .A3(wdata[18]), .A4(n1149), 
        .Y(N1903) );
  AO22X1_LVT U1660 ( .A1(n1152), .A2(io_tval[18]), .A3(wdata[18]), .A4(n1151), 
        .Y(N1011) );
  AO22X1_LVT U1661 ( .A1(n1159), .A2(io_tval[18]), .A3(wdata[18]), .A4(n1158), 
        .Y(N1400) );
  AO21X1_LVT U1662 ( .A1(n1921), .A2(n504), .A3(n376), .Y(N1577) );
  AO22X1_LVT U1663 ( .A1(n493), .A2(n_T_44[12]), .A3(wdata[18]), .A4(n492), 
        .Y(N1509) );
  NAND2X0_LVT U1664 ( .A1(io_pmp_2_cfg_w), .A2(n1507), .Y(n1113) );
  NAND2X0_LVT U1665 ( .A1(n1488), .A2(io_ptbr_ppn[17]), .Y(n1112) );
  NAND2X0_LVT U1666 ( .A1(n1689), .A2(n_T_45[17]), .Y(n1111) );
  NAND4X0_LVT U1667 ( .A1(n1113), .A2(n1579), .A3(n1112), .A4(n1111), .Y(n1114) );
  AO21X1_LVT U1668 ( .A1(n1153), .A2(n_T_383[17]), .A3(n1114), .Y(n1118) );
  AND2X1_LVT U1669 ( .A1(n1494), .A2(io_pmp_6_addr[17]), .Y(n1117) );
  AO22X1_LVT U1670 ( .A1(n1489), .A2(reg_mepc[17]), .A3(n1162), .A4(
        io_time[17]), .Y(n1116) );
  AO22X1_LVT U1671 ( .A1(n1491), .A2(io_pmp_4_addr[17]), .A3(n1492), .A4(
        io_pmp_2_addr[17]), .Y(n1115) );
  NOR4X1_LVT U1672 ( .A1(n1118), .A2(n1117), .A3(n1116), .A4(n1115), .Y(n1119)
         );
  NAND3X0_LVT U1673 ( .A1(n1580), .A2(n1581), .A3(n1119), .Y(io_rw_rdata[17])
         );
  AO22X1_LVT U1674 ( .A1(n498), .A2(n_T_52[11]), .A3(wdata[17]), .A4(n1149), 
        .Y(N1902) );
  AO22X1_LVT U1675 ( .A1(n1152), .A2(io_tval[17]), .A3(wdata[17]), .A4(n1151), 
        .Y(N1010) );
  MUX21X1_LVT U1676 ( .A1(io_pc[17]), .A2(wdata[17]), .S0(n514), .Y(net35031)
         );
  AO22X1_LVT U1677 ( .A1(n493), .A2(n_T_44[11]), .A3(wdata[17]), .A4(n1128), 
        .Y(N1508) );
  AO22X1_LVT U1678 ( .A1(n1689), .A2(n_T_45[16]), .A3(n1510), .A4(
        reg_dscratch[16]), .Y(n1120) );
  AOI21X1_LVT U1679 ( .A1(n1493), .A2(reg_dpc[16]), .A3(n1120), .Y(n1122) );
  NAND2X0_LVT U1680 ( .A1(n1153), .A2(n_T_383[16]), .Y(n1121) );
  NAND4X0_LVT U1681 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .Y(n1125) );
  OR2X1_LVT U1682 ( .A1(n1125), .A2(n1563), .Y(n1126) );
  NOR4X1_LVT U1683 ( .A1(n1562), .A2(n1561), .A3(n1126), .A4(n1569), .Y(n1127)
         );
  NAND2X0_LVT U1684 ( .A1(n1127), .A2(n1570), .Y(io_rw_rdata[16]) );
  AO22X1_LVT U1685 ( .A1(n498), .A2(n_T_52[10]), .A3(wdata[16]), .A4(n1149), 
        .Y(N1901) );
  AO22X1_LVT U1686 ( .A1(n1152), .A2(io_tval[16]), .A3(wdata[16]), .A4(n1151), 
        .Y(N1009) );
  AO22X1_LVT U1687 ( .A1(n1159), .A2(io_tval[16]), .A3(wdata[16]), .A4(n1158), 
        .Y(N1398) );
  MUX21X1_LVT U1688 ( .A1(io_pc[16]), .A2(wdata[16]), .S0(n515), .Y(net35256)
         );
  AO22X1_LVT U1689 ( .A1(n493), .A2(n_T_44[10]), .A3(wdata[16]), .A4(n492), 
        .Y(N1507) );
  AO22X1_LVT U1690 ( .A1(n494), .A2(n_T_44[5]), .A3(wdata[11]), .A4(n491), .Y(
        N1502) );
  AO22X1_LVT U1691 ( .A1(n498), .A2(n_T_52[4]), .A3(wdata[10]), .A4(n1149), 
        .Y(N1895) );
  AO22X1_LVT U1692 ( .A1(n1152), .A2(io_tval[10]), .A3(wdata[10]), .A4(n1151), 
        .Y(N1003) );
  AO22X1_LVT U1693 ( .A1(n1159), .A2(io_tval[10]), .A3(wdata[10]), .A4(n1158), 
        .Y(N1392) );
  MUX21X1_LVT U1694 ( .A1(io_pc[10]), .A2(wdata[10]), .S0(n514), .Y(net35052)
         );
  AO22X1_LVT U1695 ( .A1(n493), .A2(n_T_44[4]), .A3(wdata[10]), .A4(n491), .Y(
        N1501) );
  AO22X1_LVT U1696 ( .A1(n493), .A2(n_T_44[2]), .A3(wdata[8]), .A4(n1128), .Y(
        N1499) );
  AO22X1_LVT U1697 ( .A1(n493), .A2(n_T_44[9]), .A3(wdata[15]), .A4(n1128), 
        .Y(N1506) );
  MUX21X1_LVT U1698 ( .A1(io_pmp_1_addr[11]), .A2(wdata[11]), .S0(n506), .Y(
        n_GEN_265[11]) );
  MUX21X1_LVT U1699 ( .A1(io_pmp_6_addr[11]), .A2(wdata[11]), .S0(n511), .Y(
        n_GEN_300[11]) );
  MUX21X1_LVT U1700 ( .A1(io_pmp_2_addr[11]), .A2(wdata[11]), .S0(n507), .Y(
        n_GEN_272[11]) );
  MUX21X1_LVT U1701 ( .A1(io_pmp_3_addr[11]), .A2(wdata[11]), .S0(n508), .Y(
        n_GEN_279[11]) );
  MUX21X1_LVT U1702 ( .A1(io_pmp_5_addr[11]), .A2(wdata[11]), .S0(n510), .Y(
        n_GEN_293[11]) );
  MUX21X1_LVT U1703 ( .A1(io_pmp_4_addr[11]), .A2(wdata[11]), .S0(n509), .Y(
        n_GEN_286[11]) );
  MUX21X1_LVT U1704 ( .A1(io_pmp_0_addr[11]), .A2(wdata[11]), .S0(n505), .Y(
        n_GEN_258[11]) );
  MUX21X1_LVT U1705 ( .A1(io_pmp_7_addr[11]), .A2(wdata[11]), .S0(n512), .Y(
        n_GEN_307[11]) );
  MUX21X1_LVT U1706 ( .A1(io_pc[11]), .A2(wdata[11]), .S0(n514), .Y(net35049)
         );
  AO22X1_LVT U1707 ( .A1(reg_mie[11]), .A2(n1503), .A3(wdata[11]), .A4(n1502), 
        .Y(N617) );
  INVX1_LVT U1708 ( .A(n1692), .Y(n1130) );
  AO22X1_LVT U1709 ( .A1(n1693), .A2(n1504), .A3(n407), .A4(n1130), .Y(N607)
         );
  AO222X1_LVT U1710 ( .A1(wdata[1]), .A2(n1901), .A3(n1902), .A4(n_T_61_1), 
        .A5(n1474), .A6(n1900), .Y(n2162) );
  AND2X1_LVT U1711 ( .A1(io_rw_wdata[5]), .A2(n516), .Y(n1131) );
  AO22X1_LVT U1712 ( .A1(n1474), .A2(n1131), .A3(n_T_61_5_), .A4(n1906), .Y(
        n199) );
  INVX1_LVT U1713 ( .A(n1694), .Y(n1132) );
  AO22X1_LVT U1714 ( .A1(n1695), .A2(n1504), .A3(n427), .A4(n1132), .Y(N611)
         );
  NOR3X0_LVT U1715 ( .A1(io_status_debug), .A2(n_T_389_2), .A3(io_rw_addr[9]), 
        .Y(n1133) );
  NAND4X0_LVT U1716 ( .A1(n1134), .A2(n1133), .A3(n1519), .A4(n1517), .Y(n1135) );
  NAND2X0_LVT U1717 ( .A1(n1135), .A2(n472), .Y(n1138) );
  NAND2X0_LVT U1718 ( .A1(reg_mie[11]), .A2(io_interrupts_meip), .Y(n1188) );
  NAND2X0_LVT U1719 ( .A1(reg_mie[3]), .A2(io_interrupts_msip), .Y(n1193) );
  AND2X1_LVT U1720 ( .A1(n1188), .A2(n1193), .Y(n1183) );
  NAND2X0_LVT U1721 ( .A1(n1136), .A2(reg_mie[9]), .Y(n1171) );
  NAND2X0_LVT U1722 ( .A1(n_T_61_1), .A2(reg_mie[1]), .Y(n1178) );
  AND2X1_LVT U1723 ( .A1(n1171), .A2(n1178), .Y(n1182) );
  NAND2X0_LVT U1724 ( .A1(n_T_61_5_), .A2(reg_mie[5]), .Y(n1179) );
  NAND2X0_LVT U1725 ( .A1(reg_mie[7]), .A2(io_interrupts_mtip), .Y(n1172) );
  AND4X1_LVT U1726 ( .A1(n1179), .A2(n1172), .A3(n590), .A4(n1186), .Y(n1137)
         );
  NAND4X0_LVT U1727 ( .A1(n1138), .A2(n1183), .A3(n1182), .A4(n1137), .Y(n1140) );
  OA21X1_LVT U1728 ( .A1(n1142), .A2(io_time[2]), .A3(n1141), .Y(n1143) );
  AO22X1_LVT U1729 ( .A1(n1446), .A2(n1143), .A3(wdata[2]), .A4(n1149), .Y(
        N1824) );
  NAND2X0_LVT U1730 ( .A1(n1144), .A2(io_time[3]), .Y(n1145) );
  AOI21X1_LVT U1731 ( .A1(n1145), .A2(n454), .A3(n1147), .Y(n1146) );
  AO22X1_LVT U1732 ( .A1(n1446), .A2(n1146), .A3(wdata[4]), .A4(n1149), .Y(
        N1826) );
  AO22X1_LVT U1733 ( .A1(n1446), .A2(n1148), .A3(wdata[5]), .A4(n1149), .Y(
        N1827) );
  AO22X1_LVT U1734 ( .A1(n1149), .A2(wdata[63]), .A3(n_T_52[57]), .A4(n496), 
        .Y(N1948) );
  AO22X1_LVT U1735 ( .A1(n498), .A2(n_T_52[28]), .A3(wdata[34]), .A4(n1149), 
        .Y(N1919) );
  AO22X1_LVT U1736 ( .A1(n498), .A2(n_T_52[26]), .A3(wdata[32]), .A4(n1149), 
        .Y(N1917) );
  AO22X1_LVT U1737 ( .A1(n1150), .A2(n_T_52[2]), .A3(wdata[8]), .A4(n1149), 
        .Y(N1893) );
  AO22X1_LVT U1738 ( .A1(n1152), .A2(io_tval[8]), .A3(wdata[8]), .A4(n1151), 
        .Y(N1001) );
  AO22X1_LVT U1739 ( .A1(n1159), .A2(io_tval[8]), .A3(wdata[8]), .A4(n1158), 
        .Y(N1390) );
  AO21X1_LVT U1740 ( .A1(n1922), .A2(n504), .A3(n376), .Y(N1567) );
  MUX21X1_LVT U1741 ( .A1(io_pc[8]), .A2(wdata[8]), .S0(n513), .Y(net34856) );
  MUX21X1_LVT U1742 ( .A1(io_pc[8]), .A2(wdata[8]), .S0(n514), .Y(net35058) );
  MUX21X1_LVT U1743 ( .A1(io_pc[8]), .A2(wdata[8]), .S0(n515), .Y(net35280) );
  MUX21X1_LVT U1744 ( .A1(io_pc[5]), .A2(wdata[5]), .S0(n513), .Y(net34865) );
  MUX21X1_LVT U1745 ( .A1(io_pc[5]), .A2(wdata[5]), .S0(n514), .Y(net35067) );
  AO22X1_LVT U1746 ( .A1(io_tval[5]), .A2(n1159), .A3(wdata[5]), .A4(n1158), 
        .Y(N1387) );
  MUX21X1_LVT U1747 ( .A1(io_pc[5]), .A2(wdata[5]), .S0(n515), .Y(net35289) );
  AO22X1_LVT U1748 ( .A1(n1152), .A2(io_tval[5]), .A3(wdata[5]), .A4(n1151), 
        .Y(N998) );
  AO22X1_LVT U1749 ( .A1(n1154), .A2(n1933), .A3(n1480), .A4(io_pmp_0_addr[5]), 
        .Y(n1541) );
  MUX21X1_LVT U1750 ( .A1(io_pc[10]), .A2(wdata[10]), .S0(n515), .Y(net35274)
         );
  MUX21X1_LVT U1751 ( .A1(io_pc[10]), .A2(wdata[10]), .S0(n513), .Y(net34850)
         );
  MUX21X1_LVT U1752 ( .A1(io_pc[12]), .A2(wdata[12]), .S0(n515), .Y(net35268)
         );
  MUX21X1_LVT U1753 ( .A1(io_pc[12]), .A2(wdata[12]), .S0(n514), .Y(net35046)
         );
  MUX21X1_LVT U1754 ( .A1(io_pc[12]), .A2(wdata[12]), .S0(n513), .Y(net34844)
         );
  MUX21X1_LVT U1755 ( .A1(io_pc[13]), .A2(wdata[13]), .S0(n515), .Y(net35265)
         );
  MUX21X1_LVT U1756 ( .A1(io_pc[13]), .A2(wdata[13]), .S0(n513), .Y(net34841)
         );
  MUX21X1_LVT U1757 ( .A1(io_pc[13]), .A2(wdata[13]), .S0(n514), .Y(net35043)
         );
  MUX21X1_LVT U1758 ( .A1(io_pc[14]), .A2(wdata[14]), .S0(n515), .Y(net35262)
         );
  MUX21X1_LVT U1759 ( .A1(io_pc[14]), .A2(wdata[14]), .S0(n513), .Y(net34838)
         );
  MUX21X1_LVT U1760 ( .A1(io_pc[15]), .A2(wdata[15]), .S0(n513), .Y(net34835)
         );
  MUX21X1_LVT U1761 ( .A1(io_pc[16]), .A2(wdata[16]), .S0(n514), .Y(net35034)
         );
  MUX21X1_LVT U1762 ( .A1(io_pc[16]), .A2(wdata[16]), .S0(n513), .Y(net34832)
         );
  AO22X1_LVT U1763 ( .A1(n1157), .A2(n1927), .A3(n1480), .A4(io_pmp_0_addr[17]), .Y(n1573) );
  MUX21X1_LVT U1764 ( .A1(io_pc[17]), .A2(wdata[17]), .S0(n513), .Y(net34829)
         );
  MUX21X1_LVT U1765 ( .A1(io_pc[17]), .A2(wdata[17]), .S0(n515), .Y(net35253)
         );
  AO22X1_LVT U1766 ( .A1(n1159), .A2(io_tval[17]), .A3(wdata[17]), .A4(n1158), 
        .Y(N1399) );
  MUX21X1_LVT U1767 ( .A1(io_pc[18]), .A2(wdata[18]), .S0(n513), .Y(net34826)
         );
  MUX21X1_LVT U1768 ( .A1(io_pc[18]), .A2(wdata[18]), .S0(n514), .Y(net35028)
         );
  MUX21X1_LVT U1769 ( .A1(io_pc[18]), .A2(wdata[18]), .S0(n515), .Y(net35250)
         );
  MUX21X1_LVT U1770 ( .A1(io_pc[19]), .A2(wdata[19]), .S0(n514), .Y(net35025)
         );
  MUX21X1_LVT U1771 ( .A1(io_pc[19]), .A2(wdata[19]), .S0(n513), .Y(net34823)
         );
  MUX21X1_LVT U1772 ( .A1(io_pc[19]), .A2(wdata[19]), .S0(n515), .Y(net35247)
         );
  AO22X1_LVT U1773 ( .A1(n1689), .A2(n_T_45[19]), .A3(n1487), .A4(
        reg_stvec[19]), .Y(n1591) );
  AO22X1_LVT U1774 ( .A1(n1689), .A2(n_T_45[20]), .A3(n1487), .A4(
        reg_stvec[20]), .Y(n1596) );
  MUX21X1_LVT U1775 ( .A1(io_pc[21]), .A2(wdata[21]), .S0(n515), .Y(net35241)
         );
  MUX21X1_LVT U1776 ( .A1(io_pc[21]), .A2(wdata[21]), .S0(n513), .Y(net34817)
         );
  MUX21X1_LVT U1777 ( .A1(io_pc[22]), .A2(wdata[22]), .S0(n513), .Y(net34814)
         );
  MUX21X1_LVT U1778 ( .A1(io_pc[22]), .A2(wdata[22]), .S0(n514), .Y(net35016)
         );
  MUX21X1_LVT U1779 ( .A1(io_pc[23]), .A2(wdata[23]), .S0(n515), .Y(net35235)
         );
  AO22X1_LVT U1780 ( .A1(n1159), .A2(io_tval[23]), .A3(wdata[23]), .A4(n1158), 
        .Y(N1405) );
  MUX21X1_LVT U1781 ( .A1(io_pc[23]), .A2(wdata[23]), .S0(n513), .Y(net34811)
         );
  AO22X1_LVT U1782 ( .A1(n1160), .A2(n_T_444[23]), .A3(n1506), .A4(
        reg_sepc[23]), .Y(n1603) );
  MUX21X1_LVT U1783 ( .A1(io_pc[24]), .A2(wdata[24]), .S0(n513), .Y(net34808)
         );
  MUX21X1_LVT U1784 ( .A1(io_pc[24]), .A2(wdata[24]), .S0(n514), .Y(net35010)
         );
  MUX21X1_LVT U1785 ( .A1(io_pc[25]), .A2(wdata[25]), .S0(n514), .Y(net35007)
         );
  MUX21X1_LVT U1786 ( .A1(io_pc[25]), .A2(wdata[25]), .S0(n515), .Y(net35229)
         );
  MUX21X1_LVT U1787 ( .A1(io_pc[26]), .A2(wdata[26]), .S0(n513), .Y(net34802)
         );
  MUX21X1_LVT U1788 ( .A1(io_pc[26]), .A2(wdata[26]), .S0(n515), .Y(net35226)
         );
  MUX21X1_LVT U1789 ( .A1(io_pc[27]), .A2(wdata[27]), .S0(n514), .Y(net35001)
         );
  MUX21X1_LVT U1790 ( .A1(io_pc[27]), .A2(wdata[27]), .S0(n513), .Y(net34799)
         );
  MUX21X1_LVT U1791 ( .A1(io_pc[28]), .A2(wdata[28]), .S0(n514), .Y(net34998)
         );
  MUX21X1_LVT U1792 ( .A1(io_pc[28]), .A2(wdata[28]), .S0(n513), .Y(net34796)
         );
  MUX21X1_LVT U1793 ( .A1(io_pc[29]), .A2(wdata[29]), .S0(n513), .Y(net34793)
         );
  MUX21X1_LVT U1794 ( .A1(io_pc[30]), .A2(wdata[30]), .S0(n514), .Y(net34992)
         );
  MUX21X1_LVT U1795 ( .A1(io_pc[31]), .A2(wdata[31]), .S0(n514), .Y(net34989)
         );
  MUX21X1_LVT U1796 ( .A1(io_pc[31]), .A2(wdata[31]), .S0(n513), .Y(net34787)
         );
  MUX21X1_LVT U1797 ( .A1(io_pc[31]), .A2(wdata[31]), .S0(n515), .Y(net35211)
         );
  MUX21X1_LVT U1798 ( .A1(io_pc[32]), .A2(wdata[32]), .S0(n514), .Y(net34986)
         );
  AO22X1_LVT U1799 ( .A1(n1162), .A2(n1967), .A3(n1487), .A4(reg_stvec[32]), 
        .Y(n1630) );
  MUX21X1_LVT U1800 ( .A1(io_pc[34]), .A2(wdata[34]), .S0(n515), .Y(net35202)
         );
  AO22X1_LVT U1801 ( .A1(n1162), .A2(n1965), .A3(n1487), .A4(reg_stvec[34]), 
        .Y(n1635) );
  MUX21X1_LVT U1802 ( .A1(io_pc[34]), .A2(wdata[34]), .S0(n514), .Y(net34980)
         );
  MUX21X1_LVT U1803 ( .A1(io_pc[35]), .A2(wdata[35]), .S0(n513), .Y(net34775)
         );
  MUX21X1_LVT U1804 ( .A1(io_pc[36]), .A2(wdata[36]), .S0(n514), .Y(net34974)
         );
  MUX21X1_LVT U1805 ( .A1(io_pc[36]), .A2(wdata[36]), .S0(n515), .Y(net35196)
         );
  AO22X1_LVT U1806 ( .A1(n1689), .A2(n_T_45[36]), .A3(n1487), .A4(
        reg_stvec[36]), .Y(n1640) );
  MUX21X1_LVT U1807 ( .A1(io_pc[37]), .A2(wdata[37]), .S0(n514), .Y(net34971)
         );
  MUX21X1_LVT U1808 ( .A1(io_pc[37]), .A2(wdata[37]), .S0(n515), .Y(net35193)
         );
  MUX21X1_LVT U1809 ( .A1(io_pc[37]), .A2(wdata[37]), .S0(n513), .Y(net34769)
         );
  MUX21X1_LVT U1810 ( .A1(io_pc[39]), .A2(wdata[39]), .S0(n514), .Y(net34965)
         );
  MUX21X1_LVT U1811 ( .A1(io_pc[39]), .A2(wdata[39]), .S0(n513), .Y(net34763)
         );
  MUX21X1_LVT U1812 ( .A1(io_pc[2]), .A2(wdata[2]), .S0(n513), .Y(net34874) );
  MUX21X1_LVT U1813 ( .A1(io_pc[2]), .A2(wdata[2]), .S0(n514), .Y(net35076) );
  MUX21X1_LVT U1814 ( .A1(n1483), .A2(n477), .S0(n1163), .Y(n1166) );
  NAND2X0_LVT U1815 ( .A1(n1164), .A2(io_fcsr_flags_bits[2]), .Y(n1165) );
  NAND2X0_LVT U1816 ( .A1(n1166), .A2(n1165), .Y(n_GEN_345[2]) );
  AO22X1_LVT U1817 ( .A1(read_fcsr[2]), .A2(n1167), .A3(n1465), .A4(
        read_scounteren[2]), .Y(n1663) );
  AO22X1_LVT U1818 ( .A1(n1481), .A2(io_bp_0_control_x), .A3(n1495), .A4(
        n_T_389_2), .Y(n1666) );
  MUX21X1_LVT U1819 ( .A1(io_pc[4]), .A2(wdata[4]), .S0(n514), .Y(net35070) );
  MUX21X1_LVT U1820 ( .A1(io_pc[4]), .A2(wdata[4]), .S0(n515), .Y(net35292) );
  MUX21X1_LVT U1821 ( .A1(io_pc[4]), .A2(wdata[4]), .S0(n513), .Y(net34868) );
  MUX21X1_LVT U1822 ( .A1(io_pc[6]), .A2(wdata[6]), .S0(n515), .Y(net35286) );
  MUX21X1_LVT U1823 ( .A1(io_pc[6]), .A2(wdata[6]), .S0(n514), .Y(net35064) );
  INVX1_LVT U1824 ( .A(n1553), .Y(n1691) );
  INVX1_LVT U1825 ( .A(n_T_241[9]), .Y(n1698) );
  INVX1_LVT U1826 ( .A(n_T_241[11]), .Y(n1699) );
  INVX1_LVT U1827 ( .A(n_T_241[13]), .Y(n1700) );
  INVX1_LVT U1828 ( .A(n_T_241[14]), .Y(n1701) );
  INVX1_LVT U1829 ( .A(n_T_241[15]), .Y(n1702) );
  INVX1_LVT U1830 ( .A(n_T_241[16]), .Y(n1703) );
  INVX1_LVT U1831 ( .A(n_T_241[17]), .Y(n1704) );
  INVX1_LVT U1832 ( .A(n_T_241[18]), .Y(n1705) );
  INVX1_LVT U1833 ( .A(n_T_241[19]), .Y(n1706) );
  INVX1_LVT U1834 ( .A(n_T_241[20]), .Y(n1707) );
  INVX1_LVT U1835 ( .A(n_T_241[21]), .Y(n1708) );
  INVX1_LVT U1836 ( .A(n_T_241[22]), .Y(n1709) );
  INVX1_LVT U1837 ( .A(n_T_241[23]), .Y(n1710) );
  INVX1_LVT U1838 ( .A(n_T_241[24]), .Y(n1711) );
  INVX1_LVT U1839 ( .A(n_T_241[25]), .Y(n1712) );
  INVX1_LVT U1840 ( .A(n_T_241[26]), .Y(n1713) );
  INVX1_LVT U1841 ( .A(n_T_241[27]), .Y(n1714) );
  INVX1_LVT U1842 ( .A(n_T_241[28]), .Y(n1715) );
  INVX1_LVT U1843 ( .A(n_T_241[29]), .Y(n1716) );
  INVX1_LVT U1844 ( .A(n_T_241[1]), .Y(n1717) );
  INVX1_LVT U1845 ( .A(n_T_241[2]), .Y(n1718) );
  INVX1_LVT U1846 ( .A(n_T_241[3]), .Y(n1719) );
  INVX1_LVT U1847 ( .A(n_T_241[5]), .Y(n1720) );
  INVX1_LVT U1848 ( .A(n_T_241[6]), .Y(n1721) );
  INVX1_LVT U1849 ( .A(n_T_241[7]), .Y(n1722) );
  INVX1_LVT U1850 ( .A(n_T_250[9]), .Y(n1723) );
  INVX1_LVT U1851 ( .A(n_T_250[11]), .Y(n1724) );
  INVX1_LVT U1852 ( .A(n_T_250[13]), .Y(n1725) );
  INVX1_LVT U1853 ( .A(n_T_250[14]), .Y(n1726) );
  INVX1_LVT U1854 ( .A(n_T_250[15]), .Y(n1727) );
  INVX1_LVT U1855 ( .A(n_T_250[16]), .Y(n1728) );
  INVX1_LVT U1856 ( .A(n_T_250[17]), .Y(n1729) );
  INVX1_LVT U1857 ( .A(n_T_250[18]), .Y(n1730) );
  INVX1_LVT U1858 ( .A(n_T_250[19]), .Y(n1731) );
  INVX1_LVT U1859 ( .A(n_T_250[20]), .Y(n1732) );
  INVX1_LVT U1860 ( .A(n_T_250[21]), .Y(n1733) );
  INVX1_LVT U1861 ( .A(n_T_250[22]), .Y(n1734) );
  INVX1_LVT U1862 ( .A(n_T_250[23]), .Y(n1735) );
  INVX1_LVT U1863 ( .A(n_T_250[24]), .Y(n1736) );
  INVX1_LVT U1864 ( .A(n_T_250[25]), .Y(n1737) );
  INVX1_LVT U1865 ( .A(n_T_250[26]), .Y(n1738) );
  INVX1_LVT U1866 ( .A(n_T_250[27]), .Y(n1739) );
  INVX1_LVT U1867 ( .A(n_T_250[28]), .Y(n1740) );
  INVX1_LVT U1868 ( .A(n_T_250[29]), .Y(n1741) );
  INVX1_LVT U1869 ( .A(n_T_250[1]), .Y(n1742) );
  INVX1_LVT U1870 ( .A(n_T_250[2]), .Y(n1743) );
  INVX1_LVT U1871 ( .A(n_T_250[3]), .Y(n1744) );
  INVX1_LVT U1872 ( .A(n_T_250[5]), .Y(n1745) );
  INVX1_LVT U1873 ( .A(n_T_250[6]), .Y(n1746) );
  INVX1_LVT U1874 ( .A(n_T_250[7]), .Y(n1747) );
  INVX1_LVT U1875 ( .A(n_T_259[9]), .Y(n1748) );
  INVX1_LVT U1876 ( .A(n_T_259[11]), .Y(n1749) );
  INVX1_LVT U1877 ( .A(n_T_259[13]), .Y(n1750) );
  INVX1_LVT U1878 ( .A(n_T_259[14]), .Y(n1751) );
  INVX1_LVT U1879 ( .A(n_T_259[15]), .Y(n1752) );
  INVX1_LVT U1880 ( .A(n_T_259[16]), .Y(n1753) );
  INVX1_LVT U1881 ( .A(n_T_259[17]), .Y(n1754) );
  INVX1_LVT U1882 ( .A(n_T_259[18]), .Y(n1755) );
  INVX1_LVT U1883 ( .A(n_T_259[19]), .Y(n1756) );
  INVX1_LVT U1884 ( .A(n_T_259[20]), .Y(n1757) );
  INVX1_LVT U1885 ( .A(n_T_259[21]), .Y(n1758) );
  INVX1_LVT U1886 ( .A(n_T_259[22]), .Y(n1759) );
  INVX1_LVT U1887 ( .A(n_T_259[23]), .Y(n1760) );
  INVX1_LVT U1888 ( .A(n_T_259[24]), .Y(n1761) );
  INVX1_LVT U1889 ( .A(n_T_259[25]), .Y(n1762) );
  INVX1_LVT U1890 ( .A(n_T_259[26]), .Y(n1763) );
  INVX1_LVT U1891 ( .A(n_T_259[27]), .Y(n1764) );
  INVX1_LVT U1892 ( .A(n_T_259[28]), .Y(n1765) );
  INVX1_LVT U1893 ( .A(n_T_259[29]), .Y(n1766) );
  INVX1_LVT U1894 ( .A(n_T_259[1]), .Y(n1767) );
  INVX1_LVT U1895 ( .A(n_T_259[2]), .Y(n1768) );
  INVX1_LVT U1896 ( .A(n_T_259[3]), .Y(n1769) );
  INVX1_LVT U1897 ( .A(n_T_259[5]), .Y(n1770) );
  INVX1_LVT U1898 ( .A(n_T_259[6]), .Y(n1771) );
  INVX1_LVT U1899 ( .A(n_T_259[7]), .Y(n1772) );
  INVX1_LVT U1900 ( .A(n_T_268[9]), .Y(n1773) );
  INVX1_LVT U1901 ( .A(n_T_268[11]), .Y(n1774) );
  INVX1_LVT U1902 ( .A(n_T_268[13]), .Y(n1775) );
  INVX1_LVT U1903 ( .A(n_T_268[14]), .Y(n1776) );
  INVX1_LVT U1904 ( .A(n_T_268[15]), .Y(n1777) );
  INVX1_LVT U1905 ( .A(n_T_268[16]), .Y(n1778) );
  INVX1_LVT U1906 ( .A(n_T_268[17]), .Y(n1779) );
  INVX1_LVT U1907 ( .A(n_T_268[18]), .Y(n1780) );
  INVX1_LVT U1908 ( .A(n_T_268[19]), .Y(n1781) );
  INVX1_LVT U1909 ( .A(n_T_268[20]), .Y(n1782) );
  INVX1_LVT U1910 ( .A(n_T_268[21]), .Y(n1783) );
  INVX1_LVT U1911 ( .A(n_T_268[22]), .Y(n1784) );
  INVX1_LVT U1912 ( .A(n_T_268[23]), .Y(n1785) );
  INVX1_LVT U1913 ( .A(n_T_268[24]), .Y(n1786) );
  INVX1_LVT U1914 ( .A(n_T_268[25]), .Y(n1787) );
  INVX1_LVT U1915 ( .A(n_T_268[26]), .Y(n1788) );
  INVX1_LVT U1916 ( .A(n_T_268[27]), .Y(n1789) );
  INVX1_LVT U1917 ( .A(n_T_268[28]), .Y(n1790) );
  INVX1_LVT U1918 ( .A(n_T_268[29]), .Y(n1791) );
  INVX1_LVT U1919 ( .A(n_T_268[1]), .Y(n1792) );
  INVX1_LVT U1920 ( .A(n_T_268[2]), .Y(n1793) );
  INVX1_LVT U1921 ( .A(n_T_268[3]), .Y(n1794) );
  INVX1_LVT U1922 ( .A(n_T_268[5]), .Y(n1795) );
  INVX1_LVT U1923 ( .A(n_T_268[6]), .Y(n1796) );
  INVX1_LVT U1924 ( .A(n_T_268[7]), .Y(n1797) );
  INVX1_LVT U1925 ( .A(n_T_277[9]), .Y(n1798) );
  INVX1_LVT U1926 ( .A(n_T_277[11]), .Y(n1799) );
  INVX1_LVT U1927 ( .A(n_T_277[13]), .Y(n1800) );
  INVX1_LVT U1928 ( .A(n_T_277[14]), .Y(n1801) );
  INVX1_LVT U1929 ( .A(n_T_277[15]), .Y(n1802) );
  INVX1_LVT U1930 ( .A(n_T_277[16]), .Y(n1803) );
  INVX1_LVT U1931 ( .A(n_T_277[17]), .Y(n1804) );
  INVX1_LVT U1932 ( .A(n_T_277[18]), .Y(n1805) );
  INVX1_LVT U1933 ( .A(n_T_277[19]), .Y(n1806) );
  INVX1_LVT U1934 ( .A(n_T_277[20]), .Y(n1807) );
  INVX1_LVT U1935 ( .A(n_T_277[21]), .Y(n1808) );
  INVX1_LVT U1936 ( .A(n_T_277[22]), .Y(n1809) );
  INVX1_LVT U1937 ( .A(n_T_277[23]), .Y(n1810) );
  INVX1_LVT U1938 ( .A(n_T_277[24]), .Y(n1811) );
  INVX1_LVT U1939 ( .A(n_T_277[25]), .Y(n1812) );
  INVX1_LVT U1940 ( .A(n_T_277[26]), .Y(n1813) );
  INVX1_LVT U1941 ( .A(n_T_277[27]), .Y(n1814) );
  INVX1_LVT U1942 ( .A(n_T_277[28]), .Y(n1815) );
  INVX1_LVT U1943 ( .A(n_T_277[29]), .Y(n1816) );
  INVX1_LVT U1944 ( .A(n_T_277[1]), .Y(n1817) );
  INVX1_LVT U1945 ( .A(n_T_277[2]), .Y(n1818) );
  INVX1_LVT U1946 ( .A(n_T_277[3]), .Y(n1819) );
  INVX1_LVT U1947 ( .A(n_T_277[5]), .Y(n1820) );
  INVX1_LVT U1948 ( .A(n_T_277[6]), .Y(n1821) );
  INVX1_LVT U1949 ( .A(n_T_277[7]), .Y(n1822) );
  INVX1_LVT U1950 ( .A(n_T_286[9]), .Y(n1823) );
  INVX1_LVT U1951 ( .A(n_T_286[11]), .Y(n1824) );
  INVX1_LVT U1952 ( .A(n_T_286[13]), .Y(n1825) );
  INVX1_LVT U1953 ( .A(n_T_286[14]), .Y(n1826) );
  INVX1_LVT U1954 ( .A(n_T_286[15]), .Y(n1827) );
  INVX1_LVT U1955 ( .A(n_T_286[16]), .Y(n1828) );
  INVX1_LVT U1956 ( .A(n_T_286[17]), .Y(n1829) );
  INVX1_LVT U1957 ( .A(n_T_286[18]), .Y(n1830) );
  INVX1_LVT U1958 ( .A(n_T_286[19]), .Y(n1831) );
  INVX1_LVT U1959 ( .A(n_T_286[20]), .Y(n1832) );
  INVX1_LVT U1960 ( .A(n_T_286[21]), .Y(n1833) );
  INVX1_LVT U1961 ( .A(n_T_286[22]), .Y(n1834) );
  INVX1_LVT U1962 ( .A(n_T_286[23]), .Y(n1835) );
  INVX1_LVT U1963 ( .A(n_T_286[24]), .Y(n1836) );
  INVX1_LVT U1964 ( .A(n_T_286[25]), .Y(n1837) );
  INVX1_LVT U1965 ( .A(n_T_286[26]), .Y(n1838) );
  INVX1_LVT U1966 ( .A(n_T_286[27]), .Y(n1839) );
  INVX1_LVT U1967 ( .A(n_T_286[28]), .Y(n1840) );
  INVX1_LVT U1968 ( .A(n_T_286[29]), .Y(n1841) );
  INVX1_LVT U1969 ( .A(n_T_286[1]), .Y(n1842) );
  INVX1_LVT U1970 ( .A(n_T_286[2]), .Y(n1843) );
  INVX1_LVT U1971 ( .A(n_T_286[3]), .Y(n1844) );
  INVX1_LVT U1972 ( .A(n_T_286[5]), .Y(n1845) );
  INVX1_LVT U1973 ( .A(n_T_286[6]), .Y(n1846) );
  INVX1_LVT U1974 ( .A(n_T_286[7]), .Y(n1847) );
  INVX1_LVT U1975 ( .A(n_T_295[9]), .Y(n1848) );
  INVX1_LVT U1976 ( .A(n_T_295[11]), .Y(n1849) );
  INVX1_LVT U1977 ( .A(n_T_295[13]), .Y(n1850) );
  INVX1_LVT U1978 ( .A(n_T_295[14]), .Y(n1851) );
  INVX1_LVT U1979 ( .A(n_T_295[15]), .Y(n1852) );
  INVX1_LVT U1980 ( .A(n_T_295[16]), .Y(n1853) );
  INVX1_LVT U1981 ( .A(n_T_295[17]), .Y(n1854) );
  INVX1_LVT U1982 ( .A(n_T_295[18]), .Y(n1855) );
  INVX1_LVT U1983 ( .A(n_T_295[19]), .Y(n1856) );
  INVX1_LVT U1984 ( .A(n_T_295[20]), .Y(n1857) );
  INVX1_LVT U1985 ( .A(n_T_295[21]), .Y(n1858) );
  INVX1_LVT U1986 ( .A(n_T_295[22]), .Y(n1859) );
  INVX1_LVT U1987 ( .A(n_T_295[23]), .Y(n1860) );
  INVX1_LVT U1988 ( .A(n_T_295[24]), .Y(n1861) );
  INVX1_LVT U1989 ( .A(n_T_295[25]), .Y(n1862) );
  INVX1_LVT U1990 ( .A(n_T_295[26]), .Y(n1863) );
  INVX1_LVT U1991 ( .A(n_T_295[27]), .Y(n1864) );
  INVX1_LVT U1992 ( .A(n_T_295[28]), .Y(n1865) );
  INVX1_LVT U1993 ( .A(n_T_295[29]), .Y(n1866) );
  INVX1_LVT U1994 ( .A(n_T_295[1]), .Y(n1867) );
  INVX1_LVT U1995 ( .A(n_T_295[2]), .Y(n1868) );
  INVX1_LVT U1996 ( .A(n_T_295[3]), .Y(n1869) );
  INVX1_LVT U1997 ( .A(n_T_295[5]), .Y(n1870) );
  INVX1_LVT U1998 ( .A(n_T_295[6]), .Y(n1871) );
  INVX1_LVT U1999 ( .A(n_T_295[7]), .Y(n1872) );
  INVX1_LVT U2000 ( .A(n_T_304[9]), .Y(n1873) );
  INVX1_LVT U2001 ( .A(n_T_304[11]), .Y(n1874) );
  INVX1_LVT U2002 ( .A(n_T_304[13]), .Y(n1875) );
  INVX1_LVT U2003 ( .A(n_T_304[14]), .Y(n1876) );
  INVX1_LVT U2004 ( .A(n_T_304[15]), .Y(n1877) );
  INVX1_LVT U2005 ( .A(n_T_304[16]), .Y(n1878) );
  INVX1_LVT U2006 ( .A(n_T_304[17]), .Y(n1879) );
  INVX1_LVT U2007 ( .A(n_T_304[18]), .Y(n1880) );
  INVX1_LVT U2008 ( .A(n_T_304[19]), .Y(n1881) );
  INVX1_LVT U2009 ( .A(n_T_304[20]), .Y(n1882) );
  INVX1_LVT U2010 ( .A(n_T_304[21]), .Y(n1883) );
  INVX1_LVT U2011 ( .A(n_T_304[22]), .Y(n1884) );
  INVX1_LVT U2012 ( .A(n_T_304[23]), .Y(n1885) );
  INVX1_LVT U2013 ( .A(n_T_304[24]), .Y(n1886) );
  INVX1_LVT U2014 ( .A(n_T_304[25]), .Y(n1887) );
  INVX1_LVT U2015 ( .A(n_T_304[26]), .Y(n1888) );
  INVX1_LVT U2016 ( .A(n_T_304[27]), .Y(n1889) );
  INVX1_LVT U2017 ( .A(n_T_304[28]), .Y(n1890) );
  INVX1_LVT U2018 ( .A(n_T_304[29]), .Y(n1891) );
  INVX1_LVT U2019 ( .A(n_T_304[1]), .Y(n1892) );
  INVX1_LVT U2020 ( .A(n_T_304[2]), .Y(n1893) );
  INVX1_LVT U2021 ( .A(n_T_304[3]), .Y(n1894) );
  INVX1_LVT U2022 ( .A(n_T_304[5]), .Y(n1895) );
  INVX1_LVT U2023 ( .A(n_T_304[6]), .Y(n1896) );
  INVX1_LVT U2024 ( .A(n_T_304[7]), .Y(n1897) );
  NOR2X0_LVT U2025 ( .A1(n_T_304[4]), .A2(n412), .Y(io_pmp_7_mask[6]) );
  NOR2X0_LVT U2026 ( .A1(n_T_304[8]), .A2(n394), .Y(io_pmp_7_mask[10]) );
  NOR2X0_LVT U2027 ( .A1(n_T_304[10]), .A2(n424), .Y(io_pmp_7_mask[12]) );
  NOR2X0_LVT U2028 ( .A1(n_T_304[12]), .A2(n403), .Y(io_pmp_7_mask[14]) );
  NOR2X0_LVT U2029 ( .A1(n_T_295[4]), .A2(n413), .Y(io_pmp_6_mask[6]) );
  NOR2X0_LVT U2030 ( .A1(n_T_295[8]), .A2(n391), .Y(io_pmp_6_mask[10]) );
  NOR2X0_LVT U2031 ( .A1(n_T_295[10]), .A2(n420), .Y(io_pmp_6_mask[12]) );
  NOR2X0_LVT U2032 ( .A1(n_T_295[12]), .A2(n404), .Y(io_pmp_6_mask[14]) );
  NOR2X0_LVT U2033 ( .A1(n_T_286[4]), .A2(n414), .Y(io_pmp_5_mask[6]) );
  NOR2X0_LVT U2034 ( .A1(n_T_286[8]), .A2(n392), .Y(io_pmp_5_mask[10]) );
  NOR2X0_LVT U2035 ( .A1(n_T_286[10]), .A2(n422), .Y(io_pmp_5_mask[12]) );
  NOR2X0_LVT U2036 ( .A1(n_T_286[12]), .A2(n399), .Y(io_pmp_5_mask[14]) );
  NOR2X0_LVT U2037 ( .A1(n_T_277[4]), .A2(n408), .Y(io_pmp_4_mask[6]) );
  NOR2X0_LVT U2038 ( .A1(n_T_277[8]), .A2(n395), .Y(io_pmp_4_mask[10]) );
  NOR2X0_LVT U2039 ( .A1(n_T_277[10]), .A2(n423), .Y(io_pmp_4_mask[12]) );
  NOR2X0_LVT U2040 ( .A1(n_T_277[12]), .A2(n400), .Y(io_pmp_4_mask[14]) );
  NOR2X0_LVT U2041 ( .A1(n_T_268[4]), .A2(n409), .Y(io_pmp_3_mask[6]) );
  NOR2X0_LVT U2042 ( .A1(n_T_268[8]), .A2(n396), .Y(io_pmp_3_mask[10]) );
  NOR2X0_LVT U2043 ( .A1(n_T_268[10]), .A2(n418), .Y(io_pmp_3_mask[12]) );
  NOR2X0_LVT U2044 ( .A1(n_T_268[12]), .A2(n401), .Y(io_pmp_3_mask[14]) );
  NOR2X0_LVT U2045 ( .A1(n_T_259[4]), .A2(n410), .Y(io_pmp_2_mask[6]) );
  NOR2X0_LVT U2046 ( .A1(n_T_259[8]), .A2(n393), .Y(io_pmp_2_mask[10]) );
  NOR2X0_LVT U2047 ( .A1(n_T_259[10]), .A2(n421), .Y(io_pmp_2_mask[12]) );
  NOR2X0_LVT U2048 ( .A1(n_T_259[12]), .A2(n405), .Y(io_pmp_2_mask[14]) );
  NOR2X0_LVT U2049 ( .A1(n_T_250[4]), .A2(n411), .Y(io_pmp_1_mask[6]) );
  NOR2X0_LVT U2050 ( .A1(n_T_250[8]), .A2(n397), .Y(io_pmp_1_mask[10]) );
  NOR2X0_LVT U2051 ( .A1(n_T_250[10]), .A2(n425), .Y(io_pmp_1_mask[12]) );
  NOR2X0_LVT U2052 ( .A1(n_T_250[12]), .A2(n402), .Y(io_pmp_1_mask[14]) );
  NOR2X0_LVT U2053 ( .A1(n_T_241[4]), .A2(n415), .Y(io_pmp_0_mask[6]) );
  NOR2X0_LVT U2054 ( .A1(n_T_241[8]), .A2(n398), .Y(io_pmp_0_mask[10]) );
  NOR2X0_LVT U2055 ( .A1(n_T_241[10]), .A2(n419), .Y(io_pmp_0_mask[12]) );
  NOR2X0_LVT U2056 ( .A1(n_T_241[12]), .A2(n406), .Y(io_pmp_0_mask[14]) );
  NAND2X0_LVT U2057 ( .A1(n383), .A2(io_status_prv[1]), .Y(n1176) );
  NAND3X0_LVT U2058 ( .A1(n1169), .A2(n427), .A3(n1176), .Y(n1174) );
  OA21X1_LVT U2059 ( .A1(n1935), .A2(n429), .A3(n381), .Y(n1175) );
  AND2X1_LVT U2060 ( .A1(n1174), .A2(n1175), .Y(n1181) );
  AND2X1_LVT U2061 ( .A1(n1181), .A2(n1170), .Y(n1191) );
  NOR3X0_LVT U2062 ( .A1(read_mideleg_9_), .A2(n1187), .A3(n1171), .Y(n1189)
         );
  NAND2X0_LVT U2063 ( .A1(n1176), .A2(n1173), .Y(n1192) );
  NAND3X0_LVT U2064 ( .A1(n1177), .A2(n407), .A3(n1176), .Y(n1190) );
  OR3X1_LVT U2065 ( .A1(io_interrupts_debug), .A2(n1184), .A3(n1180), .Y(
        io_interrupt_cause[1]) );
  OA21X1_LVT U2066 ( .A1(io_interrupts_debug), .A2(n1194), .A3(n452), .Y(n1196) );
  NOR2X0_LVT U2067 ( .A1(io_status_debug), .A2(n1918), .Y(n1195) );
  OA21X1_LVT U2068 ( .A1(n426), .A2(n1196), .A3(n1195), .Y(io_interrupt) );
  AO222X1_LVT U2069 ( .A1(n502), .A2(reg_mepc[1]), .A3(n1356), .A4(reg_dpc[1]), 
        .A5(n1355), .A6(reg_sepc[1]), .Y(n1197) );
  AND2X1_LVT U2070 ( .A1(io_status_isa_2_), .A2(n1197), .Y(io_evec[1]) );
  NAND3X0_LVT U2071 ( .A1(n1255), .A2(n1198), .A3(n1903), .Y(n1204) );
  OAI22X1_LVT U2072 ( .A1(n659), .A2(n1204), .A3(n658), .A4(n1352), .Y(n1200)
         );
  AND2X1_LVT U2073 ( .A1(n1201), .A2(n1200), .Y(n1236) );
  NAND2X0_LVT U2074 ( .A1(n1236), .A2(n1202), .Y(n1208) );
  AO22X1_LVT U2075 ( .A1(n1356), .A2(reg_dpc[2]), .A3(n1355), .A4(reg_sepc[2]), 
        .Y(n1203) );
  AOI21X1_LVT U2076 ( .A1(n502), .A2(reg_mepc[2]), .A3(n1203), .Y(n1207) );
  AND2X1_LVT U2077 ( .A1(n1348), .A2(n658), .Y(n1238) );
  NAND2X0_LVT U2078 ( .A1(n1238), .A2(reg_stvec[2]), .Y(n1206) );
  AND2X1_LVT U2079 ( .A1(n1333), .A2(n659), .Y(n1239) );
  NAND2X0_LVT U2080 ( .A1(n1239), .A2(reg_mtvec[2]), .Y(n1205) );
  NAND4X0_LVT U2081 ( .A1(n1208), .A2(n1207), .A3(n1206), .A4(n1205), .Y(
        io_evec[2]) );
  NAND2X0_LVT U2082 ( .A1(n1236), .A2(n1209), .Y(n1219) );
  NAND2X0_LVT U2083 ( .A1(reg_sepc[3]), .A2(n500), .Y(n1215) );
  NAND2X0_LVT U2084 ( .A1(reg_mepc[3]), .A2(n502), .Y(n1214) );
  NAND2X0_LVT U2085 ( .A1(n1356), .A2(reg_dpc[3]), .Y(n1213) );
  NAND3X0_LVT U2086 ( .A1(n1211), .A2(io_status_debug), .A3(n1903), .Y(n1212)
         );
  AND4X1_LVT U2087 ( .A1(n1215), .A2(n1214), .A3(n1213), .A4(n1212), .Y(n1218)
         );
  NAND2X0_LVT U2088 ( .A1(n1238), .A2(reg_stvec[3]), .Y(n1217) );
  NAND2X0_LVT U2089 ( .A1(n1239), .A2(reg_mtvec[3]), .Y(n1216) );
  NAND4X0_LVT U2090 ( .A1(n1219), .A2(n1218), .A3(n1217), .A4(n1216), .Y(
        io_evec[3]) );
  NAND2X0_LVT U2091 ( .A1(n1236), .A2(n1220), .Y(n1225) );
  AO22X1_LVT U2092 ( .A1(n1356), .A2(reg_dpc[4]), .A3(n500), .A4(reg_sepc[4]), 
        .Y(n1221) );
  AOI21X1_LVT U2093 ( .A1(n502), .A2(reg_mepc[4]), .A3(n1221), .Y(n1224) );
  NAND2X0_LVT U2094 ( .A1(n1238), .A2(reg_stvec[4]), .Y(n1223) );
  NAND2X0_LVT U2095 ( .A1(n1239), .A2(reg_mtvec[4]), .Y(n1222) );
  NAND4X0_LVT U2096 ( .A1(n1225), .A2(n1224), .A3(n1223), .A4(n1222), .Y(
        io_evec[4]) );
  NAND2X0_LVT U2097 ( .A1(n1236), .A2(n1226), .Y(n1231) );
  AO22X1_LVT U2098 ( .A1(n1356), .A2(reg_dpc[5]), .A3(n1355), .A4(reg_sepc[5]), 
        .Y(n1227) );
  AOI21X1_LVT U2099 ( .A1(n502), .A2(reg_mepc[5]), .A3(n1227), .Y(n1230) );
  NAND2X0_LVT U2100 ( .A1(n1238), .A2(reg_stvec[5]), .Y(n1229) );
  NAND2X0_LVT U2101 ( .A1(n1239), .A2(reg_mtvec[5]), .Y(n1228) );
  NAND4X0_LVT U2102 ( .A1(n1231), .A2(n1230), .A3(n1229), .A4(n1228), .Y(
        io_evec[5]) );
  AO22X1_LVT U2103 ( .A1(n1356), .A2(reg_dpc[6]), .A3(n500), .A4(reg_sepc[6]), 
        .Y(n1232) );
  AOI21X1_LVT U2104 ( .A1(n502), .A2(reg_mepc[6]), .A3(n1232), .Y(n1235) );
  NAND2X0_LVT U2105 ( .A1(n1238), .A2(reg_stvec[6]), .Y(n1234) );
  NAND2X0_LVT U2106 ( .A1(n1239), .A2(reg_mtvec[6]), .Y(n1233) );
  AO22X1_LVT U2107 ( .A1(n1356), .A2(reg_dpc[7]), .A3(n1355), .A4(reg_sepc[7]), 
        .Y(n1237) );
  AOI21X1_LVT U2108 ( .A1(n502), .A2(reg_mepc[7]), .A3(n1237), .Y(n1242) );
  NAND2X0_LVT U2109 ( .A1(n1238), .A2(reg_stvec[7]), .Y(n1241) );
  NAND2X0_LVT U2110 ( .A1(n1239), .A2(reg_mtvec[7]), .Y(n1240) );
  NAND2X0_LVT U2111 ( .A1(n1348), .A2(reg_stvec[8]), .Y(n1246) );
  AOI22X1_LVT U2112 ( .A1(n1356), .A2(reg_dpc[8]), .A3(n500), .A4(reg_sepc[8]), 
        .Y(n1245) );
  NAND2X0_LVT U2113 ( .A1(n1333), .A2(reg_mtvec[8]), .Y(n1244) );
  NAND2X0_LVT U2114 ( .A1(n502), .A2(reg_mepc[8]), .Y(n1243) );
  NAND4X0_LVT U2115 ( .A1(n1246), .A2(n1245), .A3(n1244), .A4(n1243), .Y(
        io_evec[8]) );
  NAND2X0_LVT U2116 ( .A1(n1348), .A2(reg_stvec[9]), .Y(n1250) );
  AOI22X1_LVT U2117 ( .A1(n1356), .A2(reg_dpc[9]), .A3(n1355), .A4(reg_sepc[9]), .Y(n1249) );
  NAND2X0_LVT U2118 ( .A1(n1333), .A2(reg_mtvec[9]), .Y(n1248) );
  NAND2X0_LVT U2119 ( .A1(n502), .A2(reg_mepc[9]), .Y(n1247) );
  NAND4X0_LVT U2120 ( .A1(n1250), .A2(n1249), .A3(n1248), .A4(n1247), .Y(
        io_evec[9]) );
  NAND2X0_LVT U2121 ( .A1(n1348), .A2(reg_stvec[10]), .Y(n1254) );
  AOI22X1_LVT U2122 ( .A1(n1356), .A2(reg_dpc[10]), .A3(n500), .A4(
        reg_sepc[10]), .Y(n1253) );
  NAND2X0_LVT U2123 ( .A1(n1333), .A2(reg_mtvec[10]), .Y(n1252) );
  NAND2X0_LVT U2124 ( .A1(n502), .A2(reg_mepc[10]), .Y(n1251) );
  NAND4X0_LVT U2125 ( .A1(n1254), .A2(n1253), .A3(n1252), .A4(n1251), .Y(
        io_evec[10]) );
  AND2X1_LVT U2126 ( .A1(n502), .A2(reg_mepc[11]), .Y(n1260) );
  AO22X1_LVT U2127 ( .A1(n1356), .A2(reg_dpc[11]), .A3(n500), .A4(reg_sepc[11]), .Y(n1259) );
  MUX21X1_LVT U2128 ( .A1(reg_stvec[11]), .A2(reg_mtvec[11]), .S0(n1255), .Y(
        n1256) );
  OA21X1_LVT U2129 ( .A1(n1257), .A2(n1256), .A3(n1903), .Y(n1258) );
  OR3X1_LVT U2130 ( .A1(n1260), .A2(n1259), .A3(n1258), .Y(io_evec[11]) );
  NAND2X0_LVT U2131 ( .A1(n1348), .A2(reg_stvec[12]), .Y(n1264) );
  AOI22X1_LVT U2132 ( .A1(n1356), .A2(reg_dpc[12]), .A3(n1355), .A4(
        reg_sepc[12]), .Y(n1263) );
  NAND2X0_LVT U2133 ( .A1(n1333), .A2(reg_mtvec[12]), .Y(n1262) );
  NAND2X0_LVT U2134 ( .A1(n502), .A2(reg_mepc[12]), .Y(n1261) );
  NAND4X0_LVT U2135 ( .A1(n1264), .A2(n1263), .A3(n1262), .A4(n1261), .Y(
        io_evec[12]) );
  NAND2X0_LVT U2136 ( .A1(n1348), .A2(reg_stvec[13]), .Y(n1268) );
  AOI22X1_LVT U2137 ( .A1(n1356), .A2(reg_dpc[13]), .A3(n500), .A4(
        reg_sepc[13]), .Y(n1267) );
  NAND2X0_LVT U2138 ( .A1(n1333), .A2(reg_mtvec[13]), .Y(n1266) );
  NAND2X0_LVT U2139 ( .A1(n502), .A2(reg_mepc[13]), .Y(n1265) );
  NAND4X0_LVT U2140 ( .A1(n1268), .A2(n1267), .A3(n1266), .A4(n1265), .Y(
        io_evec[13]) );
  NAND2X0_LVT U2141 ( .A1(n1348), .A2(reg_stvec[14]), .Y(n1272) );
  AOI22X1_LVT U2142 ( .A1(n1356), .A2(reg_dpc[14]), .A3(n1355), .A4(
        reg_sepc[14]), .Y(n1271) );
  NAND2X0_LVT U2143 ( .A1(n1333), .A2(reg_mtvec[14]), .Y(n1270) );
  NAND2X0_LVT U2144 ( .A1(n502), .A2(reg_mepc[14]), .Y(n1269) );
  NAND4X0_LVT U2145 ( .A1(n1272), .A2(n1271), .A3(n1270), .A4(n1269), .Y(
        io_evec[14]) );
  NAND2X0_LVT U2146 ( .A1(n1348), .A2(reg_stvec[15]), .Y(n1276) );
  AOI22X1_LVT U2147 ( .A1(n1356), .A2(reg_dpc[15]), .A3(n500), .A4(
        reg_sepc[15]), .Y(n1275) );
  NAND2X0_LVT U2148 ( .A1(n1333), .A2(reg_mtvec[15]), .Y(n1274) );
  NAND2X0_LVT U2149 ( .A1(n502), .A2(reg_mepc[15]), .Y(n1273) );
  NAND4X0_LVT U2150 ( .A1(n1276), .A2(n1275), .A3(n1274), .A4(n1273), .Y(
        io_evec[15]) );
  NAND2X0_LVT U2151 ( .A1(n1348), .A2(reg_stvec[16]), .Y(n1280) );
  AOI22X1_LVT U2152 ( .A1(n1356), .A2(reg_dpc[16]), .A3(n1355), .A4(
        reg_sepc[16]), .Y(n1279) );
  NAND2X0_LVT U2153 ( .A1(n1333), .A2(reg_mtvec[16]), .Y(n1278) );
  NAND2X0_LVT U2154 ( .A1(n502), .A2(reg_mepc[16]), .Y(n1277) );
  NAND4X0_LVT U2155 ( .A1(n1280), .A2(n1279), .A3(n1278), .A4(n1277), .Y(
        io_evec[16]) );
  NAND2X0_LVT U2156 ( .A1(n1348), .A2(reg_stvec[17]), .Y(n1284) );
  AOI22X1_LVT U2157 ( .A1(n1356), .A2(reg_dpc[17]), .A3(n1355), .A4(
        reg_sepc[17]), .Y(n1283) );
  NAND2X0_LVT U2158 ( .A1(n1333), .A2(reg_mtvec[17]), .Y(n1282) );
  NAND2X0_LVT U2159 ( .A1(n502), .A2(reg_mepc[17]), .Y(n1281) );
  NAND4X0_LVT U2160 ( .A1(n1284), .A2(n1283), .A3(n1282), .A4(n1281), .Y(
        io_evec[17]) );
  NAND2X0_LVT U2161 ( .A1(n1348), .A2(reg_stvec[18]), .Y(n1288) );
  AOI22X1_LVT U2162 ( .A1(n1356), .A2(reg_dpc[18]), .A3(n500), .A4(
        reg_sepc[18]), .Y(n1287) );
  NAND2X0_LVT U2163 ( .A1(n1333), .A2(reg_mtvec[18]), .Y(n1286) );
  NAND2X0_LVT U2164 ( .A1(n502), .A2(reg_mepc[18]), .Y(n1285) );
  NAND4X0_LVT U2165 ( .A1(n1288), .A2(n1287), .A3(n1286), .A4(n1285), .Y(
        io_evec[18]) );
  NAND2X0_LVT U2166 ( .A1(n1348), .A2(reg_stvec[19]), .Y(n1292) );
  AOI22X1_LVT U2167 ( .A1(n1356), .A2(reg_dpc[19]), .A3(n500), .A4(
        reg_sepc[19]), .Y(n1291) );
  NAND2X0_LVT U2168 ( .A1(n1333), .A2(reg_mtvec[19]), .Y(n1290) );
  NAND2X0_LVT U2169 ( .A1(n502), .A2(reg_mepc[19]), .Y(n1289) );
  NAND4X0_LVT U2170 ( .A1(n1292), .A2(n1291), .A3(n1290), .A4(n1289), .Y(
        io_evec[19]) );
  NAND2X0_LVT U2171 ( .A1(n1348), .A2(reg_stvec[20]), .Y(n1296) );
  AOI22X1_LVT U2172 ( .A1(n1356), .A2(reg_dpc[20]), .A3(n1355), .A4(
        reg_sepc[20]), .Y(n1295) );
  NAND2X0_LVT U2173 ( .A1(n1333), .A2(reg_mtvec[20]), .Y(n1294) );
  NAND2X0_LVT U2174 ( .A1(n502), .A2(reg_mepc[20]), .Y(n1293) );
  NAND4X0_LVT U2175 ( .A1(n1296), .A2(n1295), .A3(n1294), .A4(n1293), .Y(
        io_evec[20]) );
  NAND2X0_LVT U2176 ( .A1(n1348), .A2(reg_stvec[21]), .Y(n1300) );
  AOI22X1_LVT U2177 ( .A1(n1356), .A2(reg_dpc[21]), .A3(n500), .A4(
        reg_sepc[21]), .Y(n1299) );
  NAND2X0_LVT U2178 ( .A1(n1333), .A2(reg_mtvec[21]), .Y(n1298) );
  NAND2X0_LVT U2179 ( .A1(n502), .A2(reg_mepc[21]), .Y(n1297) );
  NAND4X0_LVT U2180 ( .A1(n1300), .A2(n1299), .A3(n1298), .A4(n1297), .Y(
        io_evec[21]) );
  NAND2X0_LVT U2181 ( .A1(n499), .A2(reg_stvec[22]), .Y(n1304) );
  AOI22X1_LVT U2182 ( .A1(n1356), .A2(reg_dpc[22]), .A3(n1355), .A4(
        reg_sepc[22]), .Y(n1303) );
  NAND2X0_LVT U2183 ( .A1(n1333), .A2(reg_mtvec[22]), .Y(n1302) );
  NAND2X0_LVT U2184 ( .A1(n502), .A2(reg_mepc[22]), .Y(n1301) );
  NAND4X0_LVT U2185 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), .Y(
        io_evec[22]) );
  NAND2X0_LVT U2186 ( .A1(n499), .A2(reg_stvec[23]), .Y(n1308) );
  AOI22X1_LVT U2187 ( .A1(n1356), .A2(reg_dpc[23]), .A3(n500), .A4(
        reg_sepc[23]), .Y(n1307) );
  NAND2X0_LVT U2188 ( .A1(n1333), .A2(reg_mtvec[23]), .Y(n1306) );
  NAND2X0_LVT U2189 ( .A1(n502), .A2(reg_mepc[23]), .Y(n1305) );
  NAND4X0_LVT U2190 ( .A1(n1308), .A2(n1307), .A3(n1306), .A4(n1305), .Y(
        io_evec[23]) );
  NAND2X0_LVT U2191 ( .A1(n499), .A2(reg_stvec[24]), .Y(n1312) );
  AOI22X1_LVT U2192 ( .A1(n1356), .A2(reg_dpc[24]), .A3(n1355), .A4(
        reg_sepc[24]), .Y(n1311) );
  NAND2X0_LVT U2193 ( .A1(n1333), .A2(reg_mtvec[24]), .Y(n1310) );
  NAND2X0_LVT U2194 ( .A1(n502), .A2(reg_mepc[24]), .Y(n1309) );
  NAND4X0_LVT U2195 ( .A1(n1312), .A2(n1311), .A3(n1310), .A4(n1309), .Y(
        io_evec[24]) );
  NAND2X0_LVT U2196 ( .A1(n499), .A2(reg_stvec[25]), .Y(n1316) );
  AOI22X1_LVT U2197 ( .A1(n1356), .A2(reg_dpc[25]), .A3(n500), .A4(
        reg_sepc[25]), .Y(n1315) );
  NAND2X0_LVT U2198 ( .A1(n1333), .A2(reg_mtvec[25]), .Y(n1314) );
  NAND2X0_LVT U2199 ( .A1(n502), .A2(reg_mepc[25]), .Y(n1313) );
  NAND4X0_LVT U2200 ( .A1(n1316), .A2(n1315), .A3(n1314), .A4(n1313), .Y(
        io_evec[25]) );
  NAND2X0_LVT U2201 ( .A1(n499), .A2(reg_stvec[26]), .Y(n1320) );
  AOI22X1_LVT U2202 ( .A1(n1356), .A2(reg_dpc[26]), .A3(n1355), .A4(
        reg_sepc[26]), .Y(n1319) );
  NAND2X0_LVT U2203 ( .A1(n1333), .A2(reg_mtvec[26]), .Y(n1318) );
  NAND2X0_LVT U2204 ( .A1(n502), .A2(reg_mepc[26]), .Y(n1317) );
  NAND4X0_LVT U2205 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .Y(
        io_evec[26]) );
  NAND2X0_LVT U2206 ( .A1(n499), .A2(reg_stvec[27]), .Y(n1324) );
  AOI22X1_LVT U2207 ( .A1(n1356), .A2(reg_dpc[27]), .A3(n1355), .A4(
        reg_sepc[27]), .Y(n1323) );
  NAND2X0_LVT U2208 ( .A1(n1333), .A2(reg_mtvec[27]), .Y(n1322) );
  NAND2X0_LVT U2209 ( .A1(n502), .A2(reg_mepc[27]), .Y(n1321) );
  NAND4X0_LVT U2210 ( .A1(n1324), .A2(n1323), .A3(n1322), .A4(n1321), .Y(
        io_evec[27]) );
  NAND2X0_LVT U2211 ( .A1(n499), .A2(reg_stvec[28]), .Y(n1328) );
  AOI22X1_LVT U2212 ( .A1(n1356), .A2(reg_dpc[28]), .A3(n500), .A4(
        reg_sepc[28]), .Y(n1327) );
  NAND2X0_LVT U2213 ( .A1(n1333), .A2(reg_mtvec[28]), .Y(n1326) );
  NAND2X0_LVT U2214 ( .A1(n502), .A2(reg_mepc[28]), .Y(n1325) );
  NAND4X0_LVT U2215 ( .A1(n1328), .A2(n1327), .A3(n1326), .A4(n1325), .Y(
        io_evec[28]) );
  NAND2X0_LVT U2216 ( .A1(n499), .A2(reg_stvec[29]), .Y(n1332) );
  AOI22X1_LVT U2217 ( .A1(n1356), .A2(reg_dpc[29]), .A3(n1355), .A4(
        reg_sepc[29]), .Y(n1331) );
  NAND2X0_LVT U2218 ( .A1(n1333), .A2(reg_mtvec[29]), .Y(n1330) );
  NAND2X0_LVT U2219 ( .A1(n502), .A2(reg_mepc[29]), .Y(n1329) );
  NAND4X0_LVT U2220 ( .A1(n1332), .A2(n1331), .A3(n1330), .A4(n1329), .Y(
        io_evec[29]) );
  NAND2X0_LVT U2221 ( .A1(n499), .A2(reg_stvec[31]), .Y(n1337) );
  AOI22X1_LVT U2222 ( .A1(n1356), .A2(reg_dpc[31]), .A3(n1355), .A4(
        reg_sepc[31]), .Y(n1336) );
  NAND2X0_LVT U2223 ( .A1(n1333), .A2(reg_mtvec[31]), .Y(n1335) );
  NAND2X0_LVT U2224 ( .A1(n502), .A2(reg_mepc[31]), .Y(n1334) );
  NAND4X0_LVT U2225 ( .A1(n1337), .A2(n1336), .A3(n1335), .A4(n1334), .Y(
        io_evec[31]) );
  NAND2X0_LVT U2226 ( .A1(n499), .A2(reg_stvec[32]), .Y(n1340) );
  AOI22X1_LVT U2227 ( .A1(n1356), .A2(reg_dpc[32]), .A3(n500), .A4(
        reg_sepc[32]), .Y(n1339) );
  NAND2X0_LVT U2228 ( .A1(n502), .A2(reg_mepc[32]), .Y(n1338) );
  NAND3X0_LVT U2229 ( .A1(n1340), .A2(n1339), .A3(n1338), .Y(io_evec[32]) );
  NAND2X0_LVT U2230 ( .A1(n499), .A2(reg_stvec[33]), .Y(n1343) );
  AOI22X1_LVT U2231 ( .A1(n1356), .A2(reg_dpc[33]), .A3(n1355), .A4(
        reg_sepc[33]), .Y(n1342) );
  NAND2X0_LVT U2232 ( .A1(n502), .A2(reg_mepc[33]), .Y(n1341) );
  NAND3X0_LVT U2233 ( .A1(n1343), .A2(n1342), .A3(n1341), .Y(io_evec[33]) );
  NAND2X0_LVT U2234 ( .A1(n499), .A2(reg_stvec[35]), .Y(n1347) );
  AOI22X1_LVT U2235 ( .A1(n1356), .A2(reg_dpc[35]), .A3(n1355), .A4(
        reg_sepc[35]), .Y(n1345) );
  NAND2X0_LVT U2236 ( .A1(n502), .A2(reg_mepc[35]), .Y(n1344) );
  NAND3X0_LVT U2237 ( .A1(n1347), .A2(n1345), .A3(n1344), .Y(io_evec[35]) );
  NAND2X0_LVT U2238 ( .A1(n499), .A2(reg_stvec[37]), .Y(n1351) );
  AOI22X1_LVT U2239 ( .A1(n1356), .A2(reg_dpc[37]), .A3(n1355), .A4(
        reg_sepc[37]), .Y(n1350) );
  NAND2X0_LVT U2240 ( .A1(n502), .A2(reg_mepc[37]), .Y(n1349) );
  NAND3X0_LVT U2241 ( .A1(n1351), .A2(n1350), .A3(n1349), .Y(io_evec[37]) );
  OR2X1_LVT U2242 ( .A1(n465), .A2(n1352), .Y(n1357) );
  AOI22X1_LVT U2243 ( .A1(n1356), .A2(reg_dpc[38]), .A3(n500), .A4(
        reg_sepc[38]), .Y(n1354) );
  NAND2X0_LVT U2244 ( .A1(n502), .A2(reg_mepc[38]), .Y(n1353) );
  NAND3X0_LVT U2245 ( .A1(n1357), .A2(n1354), .A3(n1353), .Y(io_evec[38]) );
  NAND2X0_LVT U2246 ( .A1(n490), .A2(n1924), .Y(n1362) );
  OR2X1_LVT U2247 ( .A1(n447), .A2(n490), .Y(n1360) );
  AO22X1_LVT U2248 ( .A1(n1407), .A2(n1925), .A3(n1924), .A4(n1417), .Y(n1358)
         );
  NAND2X0_LVT U2249 ( .A1(n1358), .A2(io_decode_0_csr[8]), .Y(n1359) );
  MUX21X1_LVT U2250 ( .A1(n1360), .A2(n1359), .S0(n1406), .Y(n1361) );
  AO21X1_LVT U2251 ( .A1(n1362), .A2(n1361), .A3(io_status_prv[1]), .Y(n1366)
         );
  INVX1_LVT U2252 ( .A(io_decode_0_csr[9]), .Y(n1383) );
  NAND2X0_LVT U2253 ( .A1(n429), .A2(io_decode_0_csr[8]), .Y(n1364) );
  NOR2X0_LVT U2254 ( .A1(n381), .A2(io_decode_0_csr[9]), .Y(n1363) );
  OA22X1_LVT U2255 ( .A1(io_status_prv[1]), .A2(n1383), .A3(n1364), .A4(n1363), 
        .Y(n1401) );
  NAND2X0_LVT U2256 ( .A1(n490), .A2(io_status_debug_BAR), .Y(n1365) );
  NAND3X0_LVT U2257 ( .A1(n1366), .A2(n1401), .A3(n1365), .Y(
        io_decode_0_system_illegal) );
  OR2X1_LVT U2258 ( .A1(io_decode_0_csr[2]), .A2(n1426), .Y(
        io_decode_0_write_flush) );
  AND2X1_LVT U2259 ( .A1(n490), .A2(io_decode_0_csr[11]), .Y(
        io_decode_0_write_illegal) );
  NAND2X0_LVT U2260 ( .A1(n1923), .A2(n1928), .Y(io_decode_0_fp_illegal) );
  AND3X1_LVT U2261 ( .A1(n1376), .A2(io_decode_0_csr[9]), .A3(
        io_decode_0_csr[8]), .Y(n1368) );
  NAND3X0_LVT U2262 ( .A1(n1384), .A2(io_decode_0_csr[7]), .A3(n490), .Y(n1381) );
  NAND4X0_LVT U2263 ( .A1(n1367), .A2(n1407), .A3(n1430), .A4(n1417), .Y(n1372) );
  NAND3X0_LVT U2264 ( .A1(n1406), .A2(io_decode_0_csr[11]), .A3(n1386), .Y(
        n1370) );
  NAND4X0_LVT U2265 ( .A1(n1379), .A2(io_decode_0_write_illegal), .A3(n1371), 
        .A4(n1406), .Y(n1398) );
  AND3X1_LVT U2266 ( .A1(n1372), .A2(n1404), .A3(n1396), .Y(n1374) );
  OR2X1_LVT U2267 ( .A1(n1392), .A2(n1373), .Y(n1389) );
  NAND3X0_LVT U2268 ( .A1(n1377), .A2(n1376), .A3(n1386), .Y(n1427) );
  NOR2X0_LVT U2269 ( .A1(io_decode_0_csr[8]), .A2(io_decode_0_csr[11]), .Y(
        io_decode_0_fp_csr) );
  NAND4X0_LVT U2270 ( .A1(n1380), .A2(n1379), .A3(io_decode_0_fp_csr), .A4(
        n1386), .Y(n1421) );
  AND2X1_LVT U2271 ( .A1(n1421), .A2(n1381), .Y(n1413) );
  AND2X1_LVT U2272 ( .A1(n1419), .A2(io_decode_0_csr[4]), .Y(n1382) );
  AO22X1_LVT U2273 ( .A1(n1427), .A2(n1390), .A3(n1413), .A4(n1382), .Y(n1387)
         );
  OA21X1_LVT U2274 ( .A1(n1383), .A2(n1427), .A3(n1426), .Y(n1414) );
  OR3X1_LVT U2275 ( .A1(n490), .A2(n1386), .A3(n1385), .Y(n1432) );
  NAND4X0_LVT U2276 ( .A1(n1387), .A2(n1414), .A3(n1417), .A4(n1432), .Y(n1388) );
  AO21X1_LVT U2277 ( .A1(n1389), .A2(n1416), .A3(n1388), .Y(n1440) );
  INVX1_LVT U2278 ( .A(n1390), .Y(n1424) );
  OAI22X1_LVT U2279 ( .A1(read_scounteren[2]), .A2(n1407), .A3(
        read_scounteren[0]), .A4(n1424), .Y(n1391) );
  NAND2X0_LVT U2280 ( .A1(n1391), .A2(n429), .Y(n1395) );
  NOR2X0_LVT U2281 ( .A1(io_decode_0_csr[2]), .A2(n1392), .Y(n1412) );
  NAND2X0_LVT U2282 ( .A1(io_decode_0_csr[1]), .A2(read_mcounteren[2]), .Y(
        n1393) );
  OAI22X1_LVT U2283 ( .A1(io_decode_0_csr[0]), .A2(n1393), .A3(n470), .A4(
        n1424), .Y(n1394) );
  AND3X1_LVT U2284 ( .A1(n1395), .A2(n1412), .A3(n1394), .Y(n1397) );
  OA22X1_LVT U2285 ( .A1(n1398), .A2(n1397), .A3(n447), .A4(n1396), .Y(n1403)
         );
  NAND4X0_LVT U2286 ( .A1(n1405), .A2(n490), .A3(io_decode_0_csr[4]), .A4(
        io_status_debug_BAR), .Y(n1400) );
  NAND2X0_LVT U2287 ( .A1(io_decode_0_fp_csr), .A2(io_decode_0_fp_illegal), 
        .Y(n1399) );
  AND3X1_LVT U2288 ( .A1(n1401), .A2(n1400), .A3(n1399), .Y(n1402) );
  OA21X1_LVT U2289 ( .A1(io_status_prv[1]), .A2(n1403), .A3(n1402), .Y(n1439)
         );
  AND3X1_LVT U2290 ( .A1(n1404), .A2(io_decode_0_csr[1]), .A3(n1432), .Y(n1411) );
  NAND3X0_LVT U2291 ( .A1(n1405), .A2(io_decode_0_csr[7]), .A3(
        io_decode_0_csr[6]), .Y(n1409) );
  NAND4X0_LVT U2292 ( .A1(n1406), .A2(io_decode_0_csr[8]), .A3(
        io_decode_0_csr[9]), .A4(n490), .Y(n1408) );
  OA21X1_LVT U2293 ( .A1(n1409), .A2(n1408), .A3(n1407), .Y(n1410) );
  NAND4X0_LVT U2294 ( .A1(n1415), .A2(n1414), .A3(n1413), .A4(n1412), .Y(n1438) );
  NAND3X0_LVT U2295 ( .A1(n1418), .A2(io_decode_0_csr[9]), .A3(n1417), .Y(
        n1423) );
  NAND2X0_LVT U2296 ( .A1(n1420), .A2(io_decode_0_csr[4]), .Y(n1425) );
  AND4X1_LVT U2297 ( .A1(n1421), .A2(io_decode_0_csr[0]), .A3(n1425), .A4(
        io_decode_0_csr[1]), .Y(n1422) );
  NAND3X0_LVT U2298 ( .A1(n1423), .A2(n1422), .A3(io_decode_0_write_flush), 
        .Y(n1431) );
  AO21X1_LVT U2299 ( .A1(n1426), .A2(n1425), .A3(n1424), .Y(n1428) );
  NAND3X0_LVT U2300 ( .A1(n1428), .A2(io_decode_0_csr[2]), .A3(n1427), .Y(
        n1429) );
  NAND3X0_LVT U2301 ( .A1(n1431), .A2(n1430), .A3(n1429), .Y(n1435) );
  NAND2X0_LVT U2302 ( .A1(n1433), .A2(io_decode_0_csr[4]), .Y(n1434) );
  NAND3X0_LVT U2303 ( .A1(n1436), .A2(n1435), .A3(n1434), .Y(n1437) );
  NAND4X0_LVT U2304 ( .A1(n1440), .A2(n1439), .A3(n1438), .A4(n1437), .Y(
        io_decode_0_read_illegal) );
  NAND2X0_LVT U2305 ( .A1(n1927), .A2(io_status_debug_BAR), .Y(n1444) );
  MUX21X1_LVT U2306 ( .A1(n[1929]), .A2(io_status_prv[1]), .S0(n1444), .Y(
        N1692) );
  MUX21X1_LVT U2307 ( .A1(n[1930]), .A2(io_status_prv[0]), .S0(n1444), .Y(
        N1691) );
  NAND2X0_LVT U2308 ( .A1(n1447), .A2(n1446), .Y(N1890) );
  OA21X1_LVT U2309 ( .A1(io_status_debug), .A2(n457), .A3(n504), .Y(n1464) );
  AND2X1_LVT U2310 ( .A1(n1481), .A2(n1464), .Y(N487) );
  OR2X1_LVT U2311 ( .A1(n376), .A2(N487), .Y(N479) );
  NAND2X0_LVT U2312 ( .A1(n450), .A2(n1448), .Y(net35183) );
  NAND2X0_LVT U2313 ( .A1(n590), .A2(n1449), .Y(N438) );
  OR2X1_LVT U2314 ( .A1(n376), .A2(n1450), .Y(N276) );
  NAND2X0_LVT U2315 ( .A1(n1451), .A2(n1461), .Y(N335) );
  NAND2X0_LVT U2316 ( .A1(io_pc[1]), .A2(n1483), .Y(n1453) );
  NAND3X0_LVT U2317 ( .A1(n1453), .A2(n504), .A3(n1452), .Y(n1454) );
  NAND2X0_LVT U2318 ( .A1(n590), .A2(n1454), .Y(N1558) );
  AND2X1_LVT U2319 ( .A1(n1463), .A2(n440), .Y(N531) );
  OR2X1_LVT U2320 ( .A1(n376), .A2(N531), .Y(N527) );
  AND2X1_LVT U2321 ( .A1(n1463), .A2(n443), .Y(N556) );
  OR2X1_LVT U2322 ( .A1(n376), .A2(N556), .Y(N551) );
  AND2X1_LVT U2323 ( .A1(n1463), .A2(n438), .Y(N568) );
  AND2X1_LVT U2324 ( .A1(n1463), .A2(n437), .Y(N580) );
  OR2X1_LVT U2325 ( .A1(n376), .A2(N580), .Y(N575) );
  AND2X1_LVT U2326 ( .A1(n1463), .A2(n439), .Y(N592) );
  OR2X1_LVT U2327 ( .A1(n376), .A2(N592), .Y(N587) );
  NAND2X0_LVT U2328 ( .A1(n449), .A2(n1461), .Y(net34961) );
  AO21X1_LVT U2329 ( .A1(n1497), .A2(n504), .A3(n376), .Y(n2165) );
  NAND2X0_LVT U2330 ( .A1(n1455), .A2(n1462), .Y(N1269) );
  NAND2X0_LVT U2331 ( .A1(n1456), .A2(n1462), .Y(N1381) );
  OR2X1_LVT U2332 ( .A1(n376), .A2(N568), .Y(N559) );
  AND2X1_LVT U2333 ( .A1(n1463), .A2(n453), .Y(N518) );
  OR2X1_LVT U2334 ( .A1(n376), .A2(N518), .Y(N515) );
  NAND2X0_LVT U2335 ( .A1(n1457), .A2(n1461), .Y(N992) );
  AO21X1_LVT U2336 ( .A1(n1459), .A2(n_T_45[5]), .A3(n1458), .Y(N1496) );
  NAND3X0_LVT U2337 ( .A1(n1461), .A2(n590), .A3(n1460), .Y(N880) );
  NAND2X0_LVT U2338 ( .A1(n448), .A2(n1462), .Y(net34759) );
  AND2X1_LVT U2339 ( .A1(n1463), .A2(n441), .Y(N542) );
  OR2X1_LVT U2340 ( .A1(n376), .A2(N542), .Y(N539) );
  AND2X1_LVT U2341 ( .A1(n1463), .A2(n442), .Y(N604) );
  OR2X1_LVT U2342 ( .A1(n376), .A2(N604), .Y(N595) );
  AND2X1_LVT U2343 ( .A1(n1490), .A2(n1464), .Y(n2163) );
  AND3X1_LVT U2344 ( .A1(io_rw_addr[8]), .A2(n1529), .A3(n1517), .Y(n1522) );
  NAND3X0_LVT U2345 ( .A1(io_rw_addr[9]), .A2(io_rw_addr[8]), .A3(n1516), .Y(
        n1525) );
  NOR3X0_LVT U2346 ( .A1(n1521), .A2(n1525), .A3(io_rw_addr[3]), .Y(n1558) );
  AND4X1_LVT U2347 ( .A1(io_rw_addr[7]), .A2(io_rw_addr[5]), .A3(n1558), .A4(
        n1513), .Y(n1523) );
  NAND3X0_LVT U2348 ( .A1(io_rw_addr[7]), .A2(io_rw_addr[5]), .A3(n1513), .Y(
        n1524) );
  AND3X1_LVT U2350 ( .A1(n1517), .A2(n1528), .A3(n1518), .Y(n1557) );
  NAND3X0_LVT U2351 ( .A1(io_rw_addr[10]), .A2(io_rw_addr[11]), .A3(n1511), 
        .Y(n1530) );
  NAND2X0_LVT U2352 ( .A1(n1674), .A2(n1530), .Y(n1531) );
  AO22X1_LVT U2353 ( .A1(n1493), .A2(reg_dpc[8]), .A3(n1497), .A4(reg_mtvec[8]), .Y(n1533) );
  AO22X1_LVT U2354 ( .A1(n1491), .A2(io_pmp_4_addr[5]), .A3(n1506), .A4(
        reg_sepc[5]), .Y(n1537) );
  AO22X1_LVT U2355 ( .A1(n1494), .A2(io_pmp_6_addr[5]), .A3(n1472), .A4(
        io_pmp_5_addr[5]), .Y(n1536) );
  AO22X1_LVT U2356 ( .A1(n488), .A2(io_ptbr_ppn[5]), .A3(n1473), .A4(
        io_pmp_3_addr[5]), .Y(n1535) );
  AO22X1_LVT U2357 ( .A1(n1492), .A2(io_pmp_2_addr[5]), .A3(n1479), .A4(
        io_pmp_7_addr[5]), .Y(n1534) );
  NAND2X0_LVT U2358 ( .A1(n1503), .A2(reg_mie[5]), .Y(n1694) );
  NAND3X0_LVT U2359 ( .A1(n1505), .A2(n1509), .A3(n_T_61_5_), .Y(n1538) );
  NAND3X0_LVT U2360 ( .A1(n1553), .A2(n1694), .A3(n1538), .Y(n1539) );
  AO22X1_LVT U2361 ( .A1(n1474), .A2(n_T_61_5_), .A3(n1493), .A4(reg_dpc[5]), 
        .Y(n1542) );
  OR3X1_LVT U2362 ( .A1(n1542), .A2(n1541), .A3(n1540), .Y(n1543) );
  AO22X1_LVT U2363 ( .A1(n1488), .A2(io_ptbr_ppn[1]), .A3(n1485), .A4(
        reg_mscratch[1]), .Y(n1546) );
  AO22X1_LVT U2364 ( .A1(n1473), .A2(io_pmp_3_addr[1]), .A3(n1496), .A4(
        io_pmp_1_addr[1]), .Y(n1545) );
  AO22X1_LVT U2365 ( .A1(n1492), .A2(io_pmp_2_addr[1]), .A3(n1480), .A4(
        io_pmp_0_addr[1]), .Y(n1547) );
  AND2X1_LVT U2366 ( .A1(n1474), .A2(n_T_61_1), .Y(n1551) );
  AO22X1_LVT U2367 ( .A1(n1494), .A2(io_pmp_6_addr[1]), .A3(n1466), .A4(
        io_fcsr_rm[1]), .Y(n1550) );
  AO22X1_LVT U2368 ( .A1(n1472), .A2(io_pmp_5_addr[1]), .A3(n1491), .A4(
        io_pmp_4_addr[1]), .Y(n1549) );
  AO22X1_LVT U2369 ( .A1(n1510), .A2(reg_dscratch[1]), .A3(n1479), .A4(
        io_pmp_7_addr[1]), .Y(n1548) );
  NAND3X0_LVT U2370 ( .A1(n1504), .A2(reg_mie[1]), .A3(n1515), .Y(n1692) );
  NAND3X0_LVT U2371 ( .A1(n1505), .A2(n1509), .A3(n_T_61_1), .Y(n1552) );
  AO22X1_LVT U2372 ( .A1(n1502), .A2(reg_mie[1]), .A3(n1465), .A4(
        read_scounteren[1]), .Y(n1554) );
  AND2X1_LVT U2374 ( .A1(io_rw_addr[10]), .A2(io_rw_addr[11]), .Y(n1556) );
  AND4X1_LVT U2375 ( .A1(io_rw_addr[1]), .A2(n1558), .A3(n1557), .A4(n1556), 
        .Y(n1656) );
  AND2X1_LVT U2376 ( .A1(io_rw_addr[0]), .A2(n1656), .Y(n1670) );
  AO22X1_LVT U2377 ( .A1(n1493), .A2(reg_dpc[13]), .A3(n1506), .A4(
        reg_sepc[13]), .Y(n1559) );
  AO22X1_LVT U2378 ( .A1(n1506), .A2(reg_sepc[15]), .A3(read_medeleg_15), .A4(
        n1469), .Y(n1560) );
  AO22X1_LVT U2379 ( .A1(n1492), .A2(io_pmp_2_addr[16]), .A3(n1496), .A4(
        io_pmp_1_addr[16]), .Y(n1563) );
  AO22X1_LVT U2380 ( .A1(n1507), .A2(io_pmp_2_cfg_r), .A3(n1508), .A4(
        reg_sscratch[16]), .Y(n1562) );
  AO22X1_LVT U2381 ( .A1(n1494), .A2(io_pmp_6_addr[16]), .A3(n1497), .A4(
        reg_mtvec[16]), .Y(n1561) );
  AO22X1_LVT U2382 ( .A1(n1472), .A2(io_pmp_5_addr[16]), .A3(n1491), .A4(
        io_pmp_4_addr[16]), .Y(n1567) );
  AO22X1_LVT U2383 ( .A1(n1473), .A2(io_pmp_3_addr[16]), .A3(n1479), .A4(
        io_pmp_7_addr[16]), .Y(n1566) );
  AO22X1_LVT U2384 ( .A1(n1485), .A2(reg_mscratch[16]), .A3(n1480), .A4(
        io_pmp_0_addr[16]), .Y(n1565) );
  AO22X1_LVT U2385 ( .A1(n1490), .A2(io_bp_0_address[16]), .A3(n1489), .A4(
        reg_mepc[16]), .Y(n1564) );
  AO22X1_LVT U2386 ( .A1(n488), .A2(io_ptbr_ppn[16]), .A3(n1506), .A4(
        reg_sepc[16]), .Y(n1568) );
  AO21X1_LVT U2387 ( .A1(n1487), .A2(reg_stvec[16]), .A3(n1568), .Y(n1569) );
  AO22X1_LVT U2388 ( .A1(n1490), .A2(io_bp_0_address[17]), .A3(n1472), .A4(
        io_pmp_5_addr[17]), .Y(n1574) );
  AO22X1_LVT U2389 ( .A1(n1496), .A2(io_pmp_1_addr[17]), .A3(n1497), .A4(
        reg_mtvec[17]), .Y(n1572) );
  AO22X1_LVT U2390 ( .A1(n1479), .A2(io_pmp_7_addr[17]), .A3(n1508), .A4(
        reg_sscratch[17]), .Y(n1571) );
  AO22X1_LVT U2391 ( .A1(n1473), .A2(io_pmp_3_addr[17]), .A3(n1485), .A4(
        reg_mscratch[17]), .Y(n1576) );
  AO22X1_LVT U2392 ( .A1(n1510), .A2(reg_dscratch[17]), .A3(n1506), .A4(
        reg_sepc[17]), .Y(n1575) );
  NAND2X0_LVT U2393 ( .A1(n1487), .A2(reg_stvec[17]), .Y(n1579) );
  AO22X1_LVT U2394 ( .A1(n1488), .A2(io_ptbr_ppn[18]), .A3(n1472), .A4(
        io_pmp_5_addr[18]), .Y(n1582) );
  AO22X1_LVT U2395 ( .A1(n1490), .A2(io_bp_0_address[18]), .A3(n1506), .A4(
        reg_sepc[18]), .Y(n1584) );
  AO22X1_LVT U2396 ( .A1(n1489), .A2(reg_mepc[18]), .A3(n1508), .A4(
        reg_sscratch[18]), .Y(n1583) );
  AO22X1_LVT U2397 ( .A1(n1485), .A2(reg_mscratch[18]), .A3(n1493), .A4(
        reg_dpc[18]), .Y(n1586) );
  AO22X1_LVT U2398 ( .A1(n1492), .A2(io_pmp_2_addr[18]), .A3(n1494), .A4(
        io_pmp_6_addr[18]), .Y(n1585) );
  AO22X1_LVT U2399 ( .A1(n1490), .A2(io_bp_0_address[19]), .A3(n1496), .A4(
        io_pmp_1_addr[19]), .Y(n1587) );
  AO22X1_LVT U2400 ( .A1(n1510), .A2(reg_dscratch[19]), .A3(n1473), .A4(
        io_pmp_3_addr[19]), .Y(n1590) );
  AO22X1_LVT U2401 ( .A1(n1489), .A2(reg_mepc[19]), .A3(n1508), .A4(
        reg_sscratch[19]), .Y(n1589) );
  AO22X1_LVT U2402 ( .A1(n1491), .A2(io_pmp_4_addr[19]), .A3(n1506), .A4(
        reg_sepc[19]), .Y(n1588) );
  AO22X1_LVT U2403 ( .A1(n1490), .A2(io_bp_0_address[20]), .A3(n1480), .A4(
        io_pmp_0_addr[20]), .Y(n1594) );
  AO22X1_LVT U2404 ( .A1(n1494), .A2(io_pmp_6_addr[20]), .A3(n1497), .A4(
        reg_mtvec[20]), .Y(n1593) );
  AO22X1_LVT U2405 ( .A1(n1473), .A2(io_pmp_3_addr[20]), .A3(n1479), .A4(
        io_pmp_7_addr[20]), .Y(n1592) );
  AO22X1_LVT U2406 ( .A1(n1472), .A2(io_pmp_5_addr[20]), .A3(n1491), .A4(
        io_pmp_4_addr[20]), .Y(n1595) );
  AO21X1_LVT U2407 ( .A1(n1496), .A2(io_pmp_1_addr[20]), .A3(n1596), .Y(n1597)
         );
  AO22X1_LVT U2408 ( .A1(n1490), .A2(io_bp_0_address[23]), .A3(n1497), .A4(
        reg_mtvec[23]), .Y(n1601) );
  AO22X1_LVT U2409 ( .A1(n1494), .A2(io_pmp_6_addr[23]), .A3(n1491), .A4(
        io_pmp_4_addr[23]), .Y(n1600) );
  AO22X1_LVT U2410 ( .A1(n1472), .A2(io_pmp_5_addr[23]), .A3(n1479), .A4(
        io_pmp_7_addr[23]), .Y(n1599) );
  AO22X1_LVT U2411 ( .A1(n1485), .A2(reg_mscratch[23]), .A3(n1493), .A4(
        reg_dpc[23]), .Y(n1598) );
  AO22X1_LVT U2412 ( .A1(n1473), .A2(io_pmp_3_addr[23]), .A3(n1496), .A4(
        io_pmp_1_addr[23]), .Y(n1602) );
  AO21X1_LVT U2413 ( .A1(n1487), .A2(reg_stvec[23]), .A3(n1603), .Y(n1604) );
  AO22X1_LVT U2414 ( .A1(n1492), .A2(io_pmp_2_addr[24]), .A3(n1479), .A4(
        io_pmp_7_addr[24]), .Y(n1607) );
  AO22X1_LVT U2415 ( .A1(n1473), .A2(io_pmp_3_addr[24]), .A3(n1496), .A4(
        io_pmp_1_addr[24]), .Y(n1606) );
  AO22X1_LVT U2416 ( .A1(n1480), .A2(io_pmp_0_addr[24]), .A3(n1491), .A4(
        io_pmp_4_addr[24]), .Y(n1611) );
  AO22X1_LVT U2417 ( .A1(n1494), .A2(io_pmp_6_addr[24]), .A3(n1472), .A4(
        io_pmp_5_addr[24]), .Y(n1610) );
  AO22X1_LVT U2418 ( .A1(n1510), .A2(reg_dscratch[24]), .A3(n1506), .A4(
        reg_sepc[24]), .Y(n1609) );
  AO22X1_LVT U2419 ( .A1(n1489), .A2(reg_mepc[24]), .A3(n1508), .A4(
        reg_sscratch[24]), .Y(n1608) );
  AO22X1_LVT U2420 ( .A1(n1490), .A2(io_bp_0_address[24]), .A3(n1485), .A4(
        reg_mscratch[24]), .Y(n1612) );
  AO22X1_LVT U2421 ( .A1(n1494), .A2(io_pmp_6_addr[27]), .A3(n1489), .A4(
        reg_mepc[27]), .Y(n1614) );
  AO22X1_LVT U2422 ( .A1(n1473), .A2(io_pmp_3_addr[27]), .A3(n1472), .A4(
        io_pmp_5_addr[27]), .Y(n1616) );
  AO22X1_LVT U2423 ( .A1(n1492), .A2(io_pmp_2_addr[27]), .A3(n1485), .A4(
        reg_mscratch[27]), .Y(n1615) );
  AO22X1_LVT U2424 ( .A1(n1490), .A2(io_bp_0_address[27]), .A3(n1480), .A4(
        io_pmp_0_addr[27]), .Y(n1619) );
  AO22X1_LVT U2425 ( .A1(n1510), .A2(reg_dscratch[27]), .A3(n1479), .A4(
        io_pmp_7_addr[27]), .Y(n1618) );
  AO22X1_LVT U2426 ( .A1(n1487), .A2(reg_stvec[27]), .A3(n1497), .A4(
        reg_mtvec[27]), .Y(n1617) );
  AO22X1_LVT U2427 ( .A1(n1494), .A2(io_pmp_6_addr[29]), .A3(n1506), .A4(
        reg_sepc[29]), .Y(n1622) );
  AO22X1_LVT U2428 ( .A1(n1510), .A2(reg_dscratch[29]), .A3(n1479), .A4(
        io_pmp_7_addr[29]), .Y(n1621) );
  AO22X1_LVT U2429 ( .A1(n1485), .A2(reg_mscratch[29]), .A3(n1472), .A4(
        io_pmp_5_addr[29]), .Y(n1620) );
  AO22X1_LVT U2430 ( .A1(n1491), .A2(io_pmp_4_addr[29]), .A3(n1508), .A4(
        reg_sscratch[29]), .Y(n1624) );
  AO22X1_LVT U2431 ( .A1(n1490), .A2(io_bp_0_address[29]), .A3(n1497), .A4(
        reg_mtvec[29]), .Y(n1623) );
  AO21X1_LVT U2432 ( .A1(n1492), .A2(io_pmp_2_addr[29]), .A3(n1670), .Y(n1626)
         );
  AO22X1_LVT U2433 ( .A1(n1473), .A2(io_pmp_3_addr[29]), .A3(n1496), .A4(
        io_pmp_1_addr[29]), .Y(n1625) );
  AO22X1_LVT U2434 ( .A1(n1508), .A2(reg_sscratch[30]), .A3(n1497), .A4(
        reg_mtvec[30]), .Y(n1628) );
  AO22X1_LVT U2435 ( .A1(n1507), .A2(io_pmp_4_cfg_r), .A3(n1508), .A4(
        reg_sscratch[32]), .Y(n1632) );
  OR4X1_LVT U2436 ( .A1(n1632), .A2(n1631), .A3(n1630), .A4(n1629), .Y(n1633)
         );
  AO22X1_LVT U2437 ( .A1(n1485), .A2(reg_mscratch[34]), .A3(n1507), .A4(
        io_pmp_4_cfg_x), .Y(n1637) );
  OR4X1_LVT U2438 ( .A1(n1637), .A2(n1636), .A3(n1635), .A4(n1634), .Y(n1638)
         );
  AO22X1_LVT U2439 ( .A1(n1489), .A2(reg_mepc[36]), .A3(n1485), .A4(
        reg_mscratch[36]), .Y(n1642) );
  AO22X1_LVT U2440 ( .A1(n1490), .A2(io_bp_0_address[36]), .A3(n1510), .A4(
        reg_dscratch[36]), .Y(n1641) );
  AO22X1_LVT U2441 ( .A1(n1493), .A2(reg_dpc[36]), .A3(n1508), .A4(
        reg_sscratch[36]), .Y(n1639) );
  OR4X1_LVT U2442 ( .A1(n1642), .A2(n1641), .A3(n1640), .A4(n1639), .Y(n1643)
         );
  AO22X1_LVT U2443 ( .A1(n1510), .A2(reg_dscratch[37]), .A3(n1489), .A4(
        reg_mepc[37]), .Y(n1647) );
  AO22X1_LVT U2444 ( .A1(n1493), .A2(reg_dpc[37]), .A3(n1506), .A4(
        reg_sepc[37]), .Y(n1646) );
  OR4X1_LVT U2445 ( .A1(n1647), .A2(n1646), .A3(n1645), .A4(n1644), .Y(n1648)
         );
  AO22X1_LVT U2446 ( .A1(n1487), .A2(reg_stvec[38]), .A3(n1490), .A4(
        io_bp_0_address[38]), .Y(n1650) );
  AO22X1_LVT U2447 ( .A1(n1489), .A2(reg_mepc[39]), .A3(n1506), .A4(
        reg_sepc[39]), .Y(n1649) );
  AND2X1_LVT U2448 ( .A1(n1485), .A2(n504), .Y(N1033) );
  AO22X1_LVT U2449 ( .A1(n1479), .A2(io_pmp_7_addr[0]), .A3(n1484), .A4(
        read_mcounteren[0]), .Y(n1653) );
  AO22X1_LVT U2450 ( .A1(n1508), .A2(reg_sscratch[0]), .A3(n1496), .A4(
        io_pmp_1_addr[0]), .Y(n1652) );
  AO22X1_LVT U2451 ( .A1(n1473), .A2(io_pmp_3_addr[0]), .A3(n1494), .A4(
        io_pmp_6_addr[0]), .Y(n1651) );
  AO22X1_LVT U2452 ( .A1(n1485), .A2(reg_mscratch[0]), .A3(read_medeleg_0), 
        .A4(n1469), .Y(n1654) );
  AO22X1_LVT U2453 ( .A1(n1472), .A2(io_pmp_5_addr[0]), .A3(n1491), .A4(
        io_pmp_4_addr[0]), .Y(n1657) );
  AO22X1_LVT U2454 ( .A1(n1487), .A2(n428), .A3(n1492), .A4(io_pmp_2_addr[0]), 
        .Y(n1655) );
  AO22X1_LVT U2455 ( .A1(n1480), .A2(io_pmp_0_addr[2]), .A3(n1491), .A4(
        io_pmp_4_addr[2]), .Y(n1659) );
  AO22X1_LVT U2456 ( .A1(n1473), .A2(io_pmp_3_addr[2]), .A3(n1508), .A4(
        reg_sscratch[2]), .Y(n1658) );
  AO22X1_LVT U2457 ( .A1(n1494), .A2(io_pmp_6_addr[2]), .A3(n1506), .A4(
        reg_sepc[2]), .Y(n1660) );
  AO22X1_LVT U2458 ( .A1(n1479), .A2(io_pmp_7_addr[2]), .A3(reg_mtvec[2]), 
        .A4(n1470), .Y(n1668) );
  AO22X1_LVT U2459 ( .A1(n1490), .A2(io_bp_0_address[2]), .A3(n1489), .A4(
        reg_mepc[2]), .Y(n1665) );
  AO22X1_LVT U2460 ( .A1(n488), .A2(io_ptbr_ppn[2]), .A3(n1472), .A4(
        io_pmp_5_addr[2]), .Y(n1662) );
  AO22X1_LVT U2461 ( .A1(n1507), .A2(io_pmp_0_cfg_x), .A3(read_medeleg[2]), 
        .A4(n1469), .Y(n1661) );
  OR3X1_LVT U2462 ( .A1(n1663), .A2(n1662), .A3(n1661), .Y(n1664) );
  OR3X1_LVT U2463 ( .A1(n1666), .A2(n1665), .A3(n1664), .Y(n1667) );
  AO22X1_LVT U2464 ( .A1(n1485), .A2(reg_mscratch[63]), .A3(n1508), .A4(
        reg_sscratch[63]), .Y(n1672) );
  AND2X1_LVT U2465 ( .A1(n1508), .A2(n504), .Y(N1422) );
  NAND2X0_LVT U2466 ( .A1(n488), .A2(n504), .Y(n1673) );
  AOI22X1_LVT U2467 ( .A1(n1507), .A2(io_pmp_5_cfg_r), .A3(n1508), .A4(
        reg_sscratch[40]), .Y(n1675) );
  AOI22X1_LVT U2468 ( .A1(n1510), .A2(reg_dscratch[41]), .A3(n1507), .A4(
        io_pmp_5_cfg_w), .Y(n1676) );
  AOI22X1_LVT U2469 ( .A1(n1510), .A2(reg_dscratch[42]), .A3(n1485), .A4(
        reg_mscratch[42]), .Y(n1677) );
  AOI22X1_LVT U2470 ( .A1(n1510), .A2(reg_dscratch[43]), .A3(n1485), .A4(
        reg_mscratch[43]), .Y(n1678) );
  AOI22X1_LVT U2471 ( .A1(n1510), .A2(reg_dscratch[47]), .A3(n1508), .A4(
        reg_sscratch[47]), .Y(n1680) );
  AOI22X1_LVT U2472 ( .A1(n1510), .A2(reg_dscratch[48]), .A3(n1485), .A4(
        reg_mscratch[48]), .Y(n1681) );
  AOI22X1_LVT U2473 ( .A1(n1510), .A2(reg_dscratch[49]), .A3(n1508), .A4(
        reg_sscratch[49]), .Y(n1682) );
  AOI22X1_LVT U2474 ( .A1(n1485), .A2(reg_mscratch[50]), .A3(n1507), .A4(
        io_pmp_6_cfg_x), .Y(n1683) );
  AOI22X1_LVT U2475 ( .A1(n1510), .A2(reg_dscratch[51]), .A3(n1485), .A4(
        reg_mscratch[51]), .Y(n1684) );
  AOI22X1_LVT U2476 ( .A1(n1510), .A2(reg_dscratch[52]), .A3(n1508), .A4(
        reg_sscratch[52]), .Y(n1685) );
  AOI22X1_LVT U2477 ( .A1(n1507), .A2(io_pmp_7_cfg_r), .A3(n1508), .A4(
        reg_sscratch[56]), .Y(n1686) );
  AOI22X1_LVT U2478 ( .A1(n1485), .A2(reg_mscratch[57]), .A3(n1508), .A4(
        reg_sscratch[57]), .Y(n1687) );
  AOI22X1_LVT U2479 ( .A1(n1485), .A2(reg_mscratch[58]), .A3(n1508), .A4(
        reg_sscratch[58]), .Y(n1688) );
  AND2X1_LVT U2480 ( .A1(n504), .A2(n1691), .Y(N459) );
  AND2X1_LVT U2481 ( .A1(n504), .A2(n1469), .Y(N460) );
  AND2X1_LVT U2482 ( .A1(n1510), .A2(n504), .Y(N475) );
  OA21X1_LVT U2483 ( .A1(io_rw_addr[9]), .A2(read_mideleg_1), .A3(wdata[1]), 
        .Y(n1693) );
  OA21X1_LVT U2484 ( .A1(io_rw_addr[9]), .A2(read_mideleg_5), .A3(wdata[5]), 
        .Y(n1695) );
  AND2X1_LVT U2485 ( .A1(n1504), .A2(n504), .Y(N670) );
  AO22X1_LVT U2486 ( .A1(n1477), .A2(wdata[5]), .A3(n1696), .A4(wdata[0]), .Y(
        n_GEN_155[0]) );
  AO22X1_LVT U2487 ( .A1(n1477), .A2(wdata[6]), .A3(n1696), .A4(wdata[1]), .Y(
        n_GEN_155[1]) );
  AO22X1_LVT U2488 ( .A1(n505), .A2(wdata[0]), .A3(n430), .A4(io_pmp_0_addr[0]), .Y(n_GEN_258[0]) );
  AO22X1_LVT U2489 ( .A1(n505), .A2(wdata[10]), .A3(n430), .A4(
        io_pmp_0_addr[10]), .Y(n_GEN_258[10]) );
  AO22X1_LVT U2490 ( .A1(n505), .A2(wdata[12]), .A3(n430), .A4(
        io_pmp_0_addr[12]), .Y(n_GEN_258[12]) );
  AO22X1_LVT U2491 ( .A1(n505), .A2(wdata[13]), .A3(n430), .A4(
        io_pmp_0_addr[13]), .Y(n_GEN_258[13]) );
  AO22X1_LVT U2492 ( .A1(n505), .A2(wdata[14]), .A3(n430), .A4(
        io_pmp_0_addr[14]), .Y(n_GEN_258[14]) );
  AO22X1_LVT U2493 ( .A1(n505), .A2(wdata[15]), .A3(n430), .A4(
        io_pmp_0_addr[15]), .Y(n_GEN_258[15]) );
  AO22X1_LVT U2494 ( .A1(n505), .A2(wdata[16]), .A3(n430), .A4(
        io_pmp_0_addr[16]), .Y(n_GEN_258[16]) );
  AO22X1_LVT U2495 ( .A1(n505), .A2(wdata[17]), .A3(n430), .A4(
        io_pmp_0_addr[17]), .Y(n_GEN_258[17]) );
  AO22X1_LVT U2496 ( .A1(n505), .A2(wdata[18]), .A3(n430), .A4(
        io_pmp_0_addr[18]), .Y(n_GEN_258[18]) );
  AO22X1_LVT U2497 ( .A1(n505), .A2(wdata[19]), .A3(n430), .A4(
        io_pmp_0_addr[19]), .Y(n_GEN_258[19]) );
  AO22X1_LVT U2498 ( .A1(n505), .A2(wdata[1]), .A3(n430), .A4(io_pmp_0_addr[1]), .Y(n_GEN_258[1]) );
  AO22X1_LVT U2499 ( .A1(n505), .A2(wdata[20]), .A3(n430), .A4(
        io_pmp_0_addr[20]), .Y(n_GEN_258[20]) );
  AO22X1_LVT U2500 ( .A1(n505), .A2(wdata[21]), .A3(n430), .A4(
        io_pmp_0_addr[21]), .Y(n_GEN_258[21]) );
  AO22X1_LVT U2501 ( .A1(n505), .A2(wdata[22]), .A3(n430), .A4(
        io_pmp_0_addr[22]), .Y(n_GEN_258[22]) );
  AO22X1_LVT U2502 ( .A1(n505), .A2(wdata[23]), .A3(n430), .A4(
        io_pmp_0_addr[23]), .Y(n_GEN_258[23]) );
  AO22X1_LVT U2503 ( .A1(n505), .A2(wdata[24]), .A3(n430), .A4(
        io_pmp_0_addr[24]), .Y(n_GEN_258[24]) );
  AO22X1_LVT U2504 ( .A1(n505), .A2(wdata[25]), .A3(n430), .A4(
        io_pmp_0_addr[25]), .Y(n_GEN_258[25]) );
  AO22X1_LVT U2505 ( .A1(n505), .A2(wdata[26]), .A3(n430), .A4(
        io_pmp_0_addr[26]), .Y(n_GEN_258[26]) );
  AO22X1_LVT U2506 ( .A1(n505), .A2(wdata[27]), .A3(n430), .A4(
        io_pmp_0_addr[27]), .Y(n_GEN_258[27]) );
  AO22X1_LVT U2507 ( .A1(n505), .A2(wdata[28]), .A3(n430), .A4(
        io_pmp_0_addr[28]), .Y(n_GEN_258[28]) );
  AO22X1_LVT U2508 ( .A1(n505), .A2(wdata[29]), .A3(n430), .A4(
        io_pmp_0_addr[29]), .Y(n_GEN_258[29]) );
  AO22X1_LVT U2509 ( .A1(n505), .A2(wdata[2]), .A3(n430), .A4(io_pmp_0_addr[2]), .Y(n_GEN_258[2]) );
  AO22X1_LVT U2510 ( .A1(n505), .A2(wdata[4]), .A3(n430), .A4(io_pmp_0_addr[4]), .Y(n_GEN_258[4]) );
  AO22X1_LVT U2511 ( .A1(n505), .A2(wdata[5]), .A3(n430), .A4(io_pmp_0_addr[5]), .Y(n_GEN_258[5]) );
  AO22X1_LVT U2512 ( .A1(n505), .A2(wdata[6]), .A3(n430), .A4(io_pmp_0_addr[6]), .Y(n_GEN_258[6]) );
  AO22X1_LVT U2513 ( .A1(n505), .A2(wdata[8]), .A3(n430), .A4(io_pmp_0_addr[8]), .Y(n_GEN_258[8]) );
  AO22X1_LVT U2514 ( .A1(n506), .A2(wdata[0]), .A3(n431), .A4(io_pmp_1_addr[0]), .Y(n_GEN_265[0]) );
  AO22X1_LVT U2515 ( .A1(n506), .A2(wdata[10]), .A3(n431), .A4(
        io_pmp_1_addr[10]), .Y(n_GEN_265[10]) );
  AO22X1_LVT U2516 ( .A1(n506), .A2(wdata[12]), .A3(n431), .A4(
        io_pmp_1_addr[12]), .Y(n_GEN_265[12]) );
  AO22X1_LVT U2517 ( .A1(n506), .A2(wdata[13]), .A3(n431), .A4(
        io_pmp_1_addr[13]), .Y(n_GEN_265[13]) );
  AO22X1_LVT U2518 ( .A1(n506), .A2(wdata[14]), .A3(n431), .A4(
        io_pmp_1_addr[14]), .Y(n_GEN_265[14]) );
  AO22X1_LVT U2519 ( .A1(n506), .A2(wdata[15]), .A3(n431), .A4(
        io_pmp_1_addr[15]), .Y(n_GEN_265[15]) );
  AO22X1_LVT U2520 ( .A1(n506), .A2(wdata[16]), .A3(n431), .A4(
        io_pmp_1_addr[16]), .Y(n_GEN_265[16]) );
  AO22X1_LVT U2521 ( .A1(n506), .A2(wdata[17]), .A3(n431), .A4(
        io_pmp_1_addr[17]), .Y(n_GEN_265[17]) );
  AO22X1_LVT U2522 ( .A1(n506), .A2(wdata[18]), .A3(n431), .A4(
        io_pmp_1_addr[18]), .Y(n_GEN_265[18]) );
  AO22X1_LVT U2523 ( .A1(n506), .A2(wdata[19]), .A3(n431), .A4(
        io_pmp_1_addr[19]), .Y(n_GEN_265[19]) );
  AO22X1_LVT U2524 ( .A1(n506), .A2(wdata[1]), .A3(n431), .A4(io_pmp_1_addr[1]), .Y(n_GEN_265[1]) );
  AO22X1_LVT U2525 ( .A1(n506), .A2(wdata[20]), .A3(n431), .A4(
        io_pmp_1_addr[20]), .Y(n_GEN_265[20]) );
  AO22X1_LVT U2526 ( .A1(n506), .A2(wdata[21]), .A3(n431), .A4(
        io_pmp_1_addr[21]), .Y(n_GEN_265[21]) );
  AO22X1_LVT U2527 ( .A1(n506), .A2(wdata[22]), .A3(n431), .A4(
        io_pmp_1_addr[22]), .Y(n_GEN_265[22]) );
  AO22X1_LVT U2528 ( .A1(n506), .A2(wdata[23]), .A3(n431), .A4(
        io_pmp_1_addr[23]), .Y(n_GEN_265[23]) );
  AO22X1_LVT U2529 ( .A1(n506), .A2(wdata[24]), .A3(n431), .A4(
        io_pmp_1_addr[24]), .Y(n_GEN_265[24]) );
  AO22X1_LVT U2530 ( .A1(n506), .A2(wdata[25]), .A3(n431), .A4(
        io_pmp_1_addr[25]), .Y(n_GEN_265[25]) );
  AO22X1_LVT U2531 ( .A1(n506), .A2(wdata[26]), .A3(n431), .A4(
        io_pmp_1_addr[26]), .Y(n_GEN_265[26]) );
  AO22X1_LVT U2532 ( .A1(n506), .A2(wdata[27]), .A3(n431), .A4(
        io_pmp_1_addr[27]), .Y(n_GEN_265[27]) );
  AO22X1_LVT U2533 ( .A1(n506), .A2(wdata[28]), .A3(n431), .A4(
        io_pmp_1_addr[28]), .Y(n_GEN_265[28]) );
  AO22X1_LVT U2534 ( .A1(n506), .A2(wdata[29]), .A3(n431), .A4(
        io_pmp_1_addr[29]), .Y(n_GEN_265[29]) );
  AO22X1_LVT U2535 ( .A1(n506), .A2(wdata[2]), .A3(n431), .A4(io_pmp_1_addr[2]), .Y(n_GEN_265[2]) );
  AO22X1_LVT U2536 ( .A1(n506), .A2(wdata[4]), .A3(n431), .A4(io_pmp_1_addr[4]), .Y(n_GEN_265[4]) );
  AO22X1_LVT U2537 ( .A1(n506), .A2(wdata[5]), .A3(n431), .A4(io_pmp_1_addr[5]), .Y(n_GEN_265[5]) );
  AO22X1_LVT U2538 ( .A1(n506), .A2(wdata[6]), .A3(n431), .A4(io_pmp_1_addr[6]), .Y(n_GEN_265[6]) );
  AO22X1_LVT U2539 ( .A1(n506), .A2(wdata[8]), .A3(n431), .A4(io_pmp_1_addr[8]), .Y(n_GEN_265[8]) );
  AO22X1_LVT U2540 ( .A1(n507), .A2(wdata[0]), .A3(n432), .A4(io_pmp_2_addr[0]), .Y(n_GEN_272[0]) );
  AO22X1_LVT U2541 ( .A1(n507), .A2(wdata[10]), .A3(n432), .A4(
        io_pmp_2_addr[10]), .Y(n_GEN_272[10]) );
  AO22X1_LVT U2542 ( .A1(n507), .A2(wdata[12]), .A3(n432), .A4(
        io_pmp_2_addr[12]), .Y(n_GEN_272[12]) );
  AO22X1_LVT U2543 ( .A1(n507), .A2(wdata[13]), .A3(n432), .A4(
        io_pmp_2_addr[13]), .Y(n_GEN_272[13]) );
  AO22X1_LVT U2544 ( .A1(n507), .A2(wdata[14]), .A3(n432), .A4(
        io_pmp_2_addr[14]), .Y(n_GEN_272[14]) );
  AO22X1_LVT U2545 ( .A1(n507), .A2(wdata[15]), .A3(n432), .A4(
        io_pmp_2_addr[15]), .Y(n_GEN_272[15]) );
  AO22X1_LVT U2546 ( .A1(n507), .A2(wdata[16]), .A3(n432), .A4(
        io_pmp_2_addr[16]), .Y(n_GEN_272[16]) );
  AO22X1_LVT U2547 ( .A1(n507), .A2(wdata[17]), .A3(n432), .A4(
        io_pmp_2_addr[17]), .Y(n_GEN_272[17]) );
  AO22X1_LVT U2548 ( .A1(n507), .A2(wdata[18]), .A3(n432), .A4(
        io_pmp_2_addr[18]), .Y(n_GEN_272[18]) );
  AO22X1_LVT U2549 ( .A1(n507), .A2(wdata[19]), .A3(n432), .A4(
        io_pmp_2_addr[19]), .Y(n_GEN_272[19]) );
  AO22X1_LVT U2550 ( .A1(n507), .A2(wdata[1]), .A3(n432), .A4(io_pmp_2_addr[1]), .Y(n_GEN_272[1]) );
  AO22X1_LVT U2551 ( .A1(n507), .A2(wdata[20]), .A3(n432), .A4(
        io_pmp_2_addr[20]), .Y(n_GEN_272[20]) );
  AO22X1_LVT U2552 ( .A1(n507), .A2(wdata[21]), .A3(n432), .A4(
        io_pmp_2_addr[21]), .Y(n_GEN_272[21]) );
  AO22X1_LVT U2553 ( .A1(n507), .A2(wdata[22]), .A3(n432), .A4(
        io_pmp_2_addr[22]), .Y(n_GEN_272[22]) );
  AO22X1_LVT U2554 ( .A1(n507), .A2(wdata[23]), .A3(n432), .A4(
        io_pmp_2_addr[23]), .Y(n_GEN_272[23]) );
  AO22X1_LVT U2555 ( .A1(n507), .A2(wdata[24]), .A3(n432), .A4(
        io_pmp_2_addr[24]), .Y(n_GEN_272[24]) );
  AO22X1_LVT U2556 ( .A1(n507), .A2(wdata[25]), .A3(n432), .A4(
        io_pmp_2_addr[25]), .Y(n_GEN_272[25]) );
  AO22X1_LVT U2557 ( .A1(n507), .A2(wdata[26]), .A3(n432), .A4(
        io_pmp_2_addr[26]), .Y(n_GEN_272[26]) );
  AO22X1_LVT U2558 ( .A1(n507), .A2(wdata[27]), .A3(n432), .A4(
        io_pmp_2_addr[27]), .Y(n_GEN_272[27]) );
  AO22X1_LVT U2559 ( .A1(n507), .A2(wdata[28]), .A3(n432), .A4(
        io_pmp_2_addr[28]), .Y(n_GEN_272[28]) );
  AO22X1_LVT U2560 ( .A1(n507), .A2(wdata[29]), .A3(n432), .A4(
        io_pmp_2_addr[29]), .Y(n_GEN_272[29]) );
  AO22X1_LVT U2561 ( .A1(n507), .A2(wdata[2]), .A3(n432), .A4(io_pmp_2_addr[2]), .Y(n_GEN_272[2]) );
  AO22X1_LVT U2562 ( .A1(n507), .A2(wdata[4]), .A3(n432), .A4(io_pmp_2_addr[4]), .Y(n_GEN_272[4]) );
  AO22X1_LVT U2563 ( .A1(n507), .A2(wdata[5]), .A3(n432), .A4(io_pmp_2_addr[5]), .Y(n_GEN_272[5]) );
  AO22X1_LVT U2564 ( .A1(n507), .A2(wdata[6]), .A3(n432), .A4(io_pmp_2_addr[6]), .Y(n_GEN_272[6]) );
  AO22X1_LVT U2565 ( .A1(n507), .A2(wdata[8]), .A3(n432), .A4(io_pmp_2_addr[8]), .Y(n_GEN_272[8]) );
  AO22X1_LVT U2566 ( .A1(n508), .A2(wdata[0]), .A3(n436), .A4(io_pmp_3_addr[0]), .Y(n_GEN_279[0]) );
  AO22X1_LVT U2567 ( .A1(n508), .A2(wdata[10]), .A3(n436), .A4(
        io_pmp_3_addr[10]), .Y(n_GEN_279[10]) );
  AO22X1_LVT U2568 ( .A1(n508), .A2(wdata[12]), .A3(n436), .A4(
        io_pmp_3_addr[12]), .Y(n_GEN_279[12]) );
  AO22X1_LVT U2569 ( .A1(n508), .A2(wdata[13]), .A3(n436), .A4(
        io_pmp_3_addr[13]), .Y(n_GEN_279[13]) );
  AO22X1_LVT U2570 ( .A1(n508), .A2(wdata[14]), .A3(n436), .A4(
        io_pmp_3_addr[14]), .Y(n_GEN_279[14]) );
  AO22X1_LVT U2571 ( .A1(n508), .A2(wdata[15]), .A3(n436), .A4(
        io_pmp_3_addr[15]), .Y(n_GEN_279[15]) );
  AO22X1_LVT U2572 ( .A1(n508), .A2(wdata[16]), .A3(n436), .A4(
        io_pmp_3_addr[16]), .Y(n_GEN_279[16]) );
  AO22X1_LVT U2573 ( .A1(n508), .A2(wdata[17]), .A3(n436), .A4(
        io_pmp_3_addr[17]), .Y(n_GEN_279[17]) );
  AO22X1_LVT U2574 ( .A1(n508), .A2(wdata[18]), .A3(n436), .A4(
        io_pmp_3_addr[18]), .Y(n_GEN_279[18]) );
  AO22X1_LVT U2575 ( .A1(n508), .A2(wdata[19]), .A3(n436), .A4(
        io_pmp_3_addr[19]), .Y(n_GEN_279[19]) );
  AO22X1_LVT U2576 ( .A1(n508), .A2(wdata[1]), .A3(n436), .A4(io_pmp_3_addr[1]), .Y(n_GEN_279[1]) );
  AO22X1_LVT U2577 ( .A1(n508), .A2(wdata[20]), .A3(n436), .A4(
        io_pmp_3_addr[20]), .Y(n_GEN_279[20]) );
  AO22X1_LVT U2578 ( .A1(n508), .A2(wdata[21]), .A3(n436), .A4(
        io_pmp_3_addr[21]), .Y(n_GEN_279[21]) );
  AO22X1_LVT U2579 ( .A1(n508), .A2(wdata[22]), .A3(n436), .A4(
        io_pmp_3_addr[22]), .Y(n_GEN_279[22]) );
  AO22X1_LVT U2580 ( .A1(n508), .A2(wdata[23]), .A3(n436), .A4(
        io_pmp_3_addr[23]), .Y(n_GEN_279[23]) );
  AO22X1_LVT U2581 ( .A1(n508), .A2(wdata[24]), .A3(n436), .A4(
        io_pmp_3_addr[24]), .Y(n_GEN_279[24]) );
  AO22X1_LVT U2582 ( .A1(n508), .A2(wdata[25]), .A3(n436), .A4(
        io_pmp_3_addr[25]), .Y(n_GEN_279[25]) );
  AO22X1_LVT U2583 ( .A1(n508), .A2(wdata[26]), .A3(n436), .A4(
        io_pmp_3_addr[26]), .Y(n_GEN_279[26]) );
  AO22X1_LVT U2584 ( .A1(n508), .A2(wdata[27]), .A3(n436), .A4(
        io_pmp_3_addr[27]), .Y(n_GEN_279[27]) );
  AO22X1_LVT U2585 ( .A1(n508), .A2(wdata[28]), .A3(n436), .A4(
        io_pmp_3_addr[28]), .Y(n_GEN_279[28]) );
  AO22X1_LVT U2586 ( .A1(n508), .A2(wdata[29]), .A3(n436), .A4(
        io_pmp_3_addr[29]), .Y(n_GEN_279[29]) );
  AO22X1_LVT U2587 ( .A1(n508), .A2(wdata[2]), .A3(n436), .A4(io_pmp_3_addr[2]), .Y(n_GEN_279[2]) );
  AO22X1_LVT U2588 ( .A1(n508), .A2(wdata[4]), .A3(n436), .A4(io_pmp_3_addr[4]), .Y(n_GEN_279[4]) );
  AO22X1_LVT U2589 ( .A1(n508), .A2(wdata[5]), .A3(n436), .A4(io_pmp_3_addr[5]), .Y(n_GEN_279[5]) );
  AO22X1_LVT U2590 ( .A1(n508), .A2(wdata[6]), .A3(n436), .A4(io_pmp_3_addr[6]), .Y(n_GEN_279[6]) );
  AO22X1_LVT U2591 ( .A1(n508), .A2(wdata[8]), .A3(n436), .A4(io_pmp_3_addr[8]), .Y(n_GEN_279[8]) );
  AO22X1_LVT U2592 ( .A1(n509), .A2(wdata[0]), .A3(n433), .A4(io_pmp_4_addr[0]), .Y(n_GEN_286[0]) );
  AO22X1_LVT U2593 ( .A1(n509), .A2(wdata[10]), .A3(n433), .A4(
        io_pmp_4_addr[10]), .Y(n_GEN_286[10]) );
  AO22X1_LVT U2594 ( .A1(n509), .A2(wdata[12]), .A3(n433), .A4(
        io_pmp_4_addr[12]), .Y(n_GEN_286[12]) );
  AO22X1_LVT U2595 ( .A1(n509), .A2(wdata[13]), .A3(n433), .A4(
        io_pmp_4_addr[13]), .Y(n_GEN_286[13]) );
  AO22X1_LVT U2596 ( .A1(n509), .A2(wdata[14]), .A3(n433), .A4(
        io_pmp_4_addr[14]), .Y(n_GEN_286[14]) );
  AO22X1_LVT U2597 ( .A1(n509), .A2(wdata[15]), .A3(n433), .A4(
        io_pmp_4_addr[15]), .Y(n_GEN_286[15]) );
  AO22X1_LVT U2598 ( .A1(n509), .A2(wdata[16]), .A3(n433), .A4(
        io_pmp_4_addr[16]), .Y(n_GEN_286[16]) );
  AO22X1_LVT U2599 ( .A1(n509), .A2(wdata[17]), .A3(n433), .A4(
        io_pmp_4_addr[17]), .Y(n_GEN_286[17]) );
  AO22X1_LVT U2600 ( .A1(n509), .A2(wdata[18]), .A3(n433), .A4(
        io_pmp_4_addr[18]), .Y(n_GEN_286[18]) );
  AO22X1_LVT U2601 ( .A1(n509), .A2(wdata[19]), .A3(n433), .A4(
        io_pmp_4_addr[19]), .Y(n_GEN_286[19]) );
  AO22X1_LVT U2602 ( .A1(n509), .A2(wdata[1]), .A3(n433), .A4(io_pmp_4_addr[1]), .Y(n_GEN_286[1]) );
  AO22X1_LVT U2603 ( .A1(n509), .A2(wdata[20]), .A3(n433), .A4(
        io_pmp_4_addr[20]), .Y(n_GEN_286[20]) );
  AO22X1_LVT U2604 ( .A1(n509), .A2(wdata[21]), .A3(n433), .A4(
        io_pmp_4_addr[21]), .Y(n_GEN_286[21]) );
  AO22X1_LVT U2605 ( .A1(n509), .A2(wdata[22]), .A3(n433), .A4(
        io_pmp_4_addr[22]), .Y(n_GEN_286[22]) );
  AO22X1_LVT U2606 ( .A1(n509), .A2(wdata[23]), .A3(n433), .A4(
        io_pmp_4_addr[23]), .Y(n_GEN_286[23]) );
  AO22X1_LVT U2607 ( .A1(n509), .A2(wdata[24]), .A3(n433), .A4(
        io_pmp_4_addr[24]), .Y(n_GEN_286[24]) );
  AO22X1_LVT U2608 ( .A1(n509), .A2(wdata[25]), .A3(n433), .A4(
        io_pmp_4_addr[25]), .Y(n_GEN_286[25]) );
  AO22X1_LVT U2609 ( .A1(n509), .A2(wdata[26]), .A3(n433), .A4(
        io_pmp_4_addr[26]), .Y(n_GEN_286[26]) );
  AO22X1_LVT U2610 ( .A1(n509), .A2(wdata[27]), .A3(n433), .A4(
        io_pmp_4_addr[27]), .Y(n_GEN_286[27]) );
  AO22X1_LVT U2611 ( .A1(n509), .A2(wdata[28]), .A3(n433), .A4(
        io_pmp_4_addr[28]), .Y(n_GEN_286[28]) );
  AO22X1_LVT U2612 ( .A1(n509), .A2(wdata[29]), .A3(n433), .A4(
        io_pmp_4_addr[29]), .Y(n_GEN_286[29]) );
  AO22X1_LVT U2613 ( .A1(n509), .A2(wdata[2]), .A3(n433), .A4(io_pmp_4_addr[2]), .Y(n_GEN_286[2]) );
  AO22X1_LVT U2614 ( .A1(n509), .A2(wdata[4]), .A3(n433), .A4(io_pmp_4_addr[4]), .Y(n_GEN_286[4]) );
  AO22X1_LVT U2615 ( .A1(n509), .A2(wdata[5]), .A3(n433), .A4(io_pmp_4_addr[5]), .Y(n_GEN_286[5]) );
  AO22X1_LVT U2616 ( .A1(n509), .A2(wdata[6]), .A3(n433), .A4(io_pmp_4_addr[6]), .Y(n_GEN_286[6]) );
  AO22X1_LVT U2617 ( .A1(n509), .A2(wdata[8]), .A3(n433), .A4(io_pmp_4_addr[8]), .Y(n_GEN_286[8]) );
  AO22X1_LVT U2618 ( .A1(n510), .A2(wdata[0]), .A3(n434), .A4(io_pmp_5_addr[0]), .Y(n_GEN_293[0]) );
  AO22X1_LVT U2619 ( .A1(n510), .A2(wdata[10]), .A3(n434), .A4(
        io_pmp_5_addr[10]), .Y(n_GEN_293[10]) );
  AO22X1_LVT U2620 ( .A1(n510), .A2(wdata[12]), .A3(n434), .A4(
        io_pmp_5_addr[12]), .Y(n_GEN_293[12]) );
  AO22X1_LVT U2621 ( .A1(n510), .A2(wdata[13]), .A3(n434), .A4(
        io_pmp_5_addr[13]), .Y(n_GEN_293[13]) );
  AO22X1_LVT U2622 ( .A1(n510), .A2(wdata[14]), .A3(n434), .A4(
        io_pmp_5_addr[14]), .Y(n_GEN_293[14]) );
  AO22X1_LVT U2623 ( .A1(n510), .A2(wdata[15]), .A3(n434), .A4(
        io_pmp_5_addr[15]), .Y(n_GEN_293[15]) );
  AO22X1_LVT U2624 ( .A1(n510), .A2(wdata[16]), .A3(n434), .A4(
        io_pmp_5_addr[16]), .Y(n_GEN_293[16]) );
  AO22X1_LVT U2625 ( .A1(n510), .A2(wdata[17]), .A3(n434), .A4(
        io_pmp_5_addr[17]), .Y(n_GEN_293[17]) );
  AO22X1_LVT U2626 ( .A1(n510), .A2(wdata[18]), .A3(n434), .A4(
        io_pmp_5_addr[18]), .Y(n_GEN_293[18]) );
  AO22X1_LVT U2627 ( .A1(n510), .A2(wdata[19]), .A3(n434), .A4(
        io_pmp_5_addr[19]), .Y(n_GEN_293[19]) );
  AO22X1_LVT U2628 ( .A1(n510), .A2(wdata[1]), .A3(n434), .A4(io_pmp_5_addr[1]), .Y(n_GEN_293[1]) );
  AO22X1_LVT U2629 ( .A1(n510), .A2(wdata[20]), .A3(n434), .A4(
        io_pmp_5_addr[20]), .Y(n_GEN_293[20]) );
  AO22X1_LVT U2630 ( .A1(n510), .A2(wdata[21]), .A3(n434), .A4(
        io_pmp_5_addr[21]), .Y(n_GEN_293[21]) );
  AO22X1_LVT U2631 ( .A1(n510), .A2(wdata[22]), .A3(n434), .A4(
        io_pmp_5_addr[22]), .Y(n_GEN_293[22]) );
  AO22X1_LVT U2632 ( .A1(n510), .A2(wdata[23]), .A3(n434), .A4(
        io_pmp_5_addr[23]), .Y(n_GEN_293[23]) );
  AO22X1_LVT U2633 ( .A1(n510), .A2(wdata[24]), .A3(n434), .A4(
        io_pmp_5_addr[24]), .Y(n_GEN_293[24]) );
  AO22X1_LVT U2634 ( .A1(n510), .A2(wdata[25]), .A3(n434), .A4(
        io_pmp_5_addr[25]), .Y(n_GEN_293[25]) );
  AO22X1_LVT U2635 ( .A1(n510), .A2(wdata[26]), .A3(n434), .A4(
        io_pmp_5_addr[26]), .Y(n_GEN_293[26]) );
  AO22X1_LVT U2636 ( .A1(n510), .A2(wdata[27]), .A3(n434), .A4(
        io_pmp_5_addr[27]), .Y(n_GEN_293[27]) );
  AO22X1_LVT U2637 ( .A1(n510), .A2(wdata[28]), .A3(n434), .A4(
        io_pmp_5_addr[28]), .Y(n_GEN_293[28]) );
  AO22X1_LVT U2638 ( .A1(n510), .A2(wdata[29]), .A3(n434), .A4(
        io_pmp_5_addr[29]), .Y(n_GEN_293[29]) );
  AO22X1_LVT U2639 ( .A1(n510), .A2(wdata[2]), .A3(n434), .A4(io_pmp_5_addr[2]), .Y(n_GEN_293[2]) );
  AO22X1_LVT U2640 ( .A1(n510), .A2(wdata[4]), .A3(n434), .A4(io_pmp_5_addr[4]), .Y(n_GEN_293[4]) );
  AO22X1_LVT U2641 ( .A1(n510), .A2(wdata[5]), .A3(n434), .A4(io_pmp_5_addr[5]), .Y(n_GEN_293[5]) );
  AO22X1_LVT U2642 ( .A1(n510), .A2(wdata[6]), .A3(n434), .A4(io_pmp_5_addr[6]), .Y(n_GEN_293[6]) );
  AO22X1_LVT U2643 ( .A1(n510), .A2(wdata[8]), .A3(n434), .A4(io_pmp_5_addr[8]), .Y(n_GEN_293[8]) );
  AO22X1_LVT U2644 ( .A1(n511), .A2(wdata[0]), .A3(n435), .A4(io_pmp_6_addr[0]), .Y(n_GEN_300[0]) );
  AO22X1_LVT U2645 ( .A1(n511), .A2(wdata[10]), .A3(n435), .A4(
        io_pmp_6_addr[10]), .Y(n_GEN_300[10]) );
  AO22X1_LVT U2646 ( .A1(n511), .A2(wdata[12]), .A3(n435), .A4(
        io_pmp_6_addr[12]), .Y(n_GEN_300[12]) );
  AO22X1_LVT U2647 ( .A1(n511), .A2(wdata[13]), .A3(n435), .A4(
        io_pmp_6_addr[13]), .Y(n_GEN_300[13]) );
  AO22X1_LVT U2648 ( .A1(n511), .A2(wdata[14]), .A3(n435), .A4(
        io_pmp_6_addr[14]), .Y(n_GEN_300[14]) );
  AO22X1_LVT U2649 ( .A1(n511), .A2(wdata[15]), .A3(n435), .A4(
        io_pmp_6_addr[15]), .Y(n_GEN_300[15]) );
  AO22X1_LVT U2650 ( .A1(n511), .A2(wdata[16]), .A3(n435), .A4(
        io_pmp_6_addr[16]), .Y(n_GEN_300[16]) );
  AO22X1_LVT U2651 ( .A1(n511), .A2(wdata[17]), .A3(n435), .A4(
        io_pmp_6_addr[17]), .Y(n_GEN_300[17]) );
  AO22X1_LVT U2652 ( .A1(n511), .A2(wdata[18]), .A3(n435), .A4(
        io_pmp_6_addr[18]), .Y(n_GEN_300[18]) );
  AO22X1_LVT U2653 ( .A1(n511), .A2(wdata[19]), .A3(n435), .A4(
        io_pmp_6_addr[19]), .Y(n_GEN_300[19]) );
  AO22X1_LVT U2654 ( .A1(n511), .A2(wdata[1]), .A3(n435), .A4(io_pmp_6_addr[1]), .Y(n_GEN_300[1]) );
  AO22X1_LVT U2655 ( .A1(n511), .A2(wdata[20]), .A3(n435), .A4(
        io_pmp_6_addr[20]), .Y(n_GEN_300[20]) );
  AO22X1_LVT U2656 ( .A1(n511), .A2(wdata[21]), .A3(n435), .A4(
        io_pmp_6_addr[21]), .Y(n_GEN_300[21]) );
  AO22X1_LVT U2657 ( .A1(n511), .A2(wdata[22]), .A3(n435), .A4(
        io_pmp_6_addr[22]), .Y(n_GEN_300[22]) );
  AO22X1_LVT U2658 ( .A1(n511), .A2(wdata[23]), .A3(n435), .A4(
        io_pmp_6_addr[23]), .Y(n_GEN_300[23]) );
  AO22X1_LVT U2659 ( .A1(n511), .A2(wdata[24]), .A3(n435), .A4(
        io_pmp_6_addr[24]), .Y(n_GEN_300[24]) );
  AO22X1_LVT U2660 ( .A1(n511), .A2(wdata[25]), .A3(n435), .A4(
        io_pmp_6_addr[25]), .Y(n_GEN_300[25]) );
  AO22X1_LVT U2661 ( .A1(n511), .A2(wdata[26]), .A3(n435), .A4(
        io_pmp_6_addr[26]), .Y(n_GEN_300[26]) );
  AO22X1_LVT U2662 ( .A1(n511), .A2(wdata[27]), .A3(n435), .A4(
        io_pmp_6_addr[27]), .Y(n_GEN_300[27]) );
  AO22X1_LVT U2663 ( .A1(n511), .A2(wdata[28]), .A3(n435), .A4(
        io_pmp_6_addr[28]), .Y(n_GEN_300[28]) );
  AO22X1_LVT U2664 ( .A1(n511), .A2(wdata[29]), .A3(n435), .A4(
        io_pmp_6_addr[29]), .Y(n_GEN_300[29]) );
  AO22X1_LVT U2665 ( .A1(n511), .A2(wdata[2]), .A3(n435), .A4(io_pmp_6_addr[2]), .Y(n_GEN_300[2]) );
  AO22X1_LVT U2666 ( .A1(n511), .A2(wdata[4]), .A3(n435), .A4(io_pmp_6_addr[4]), .Y(n_GEN_300[4]) );
  AO22X1_LVT U2667 ( .A1(n511), .A2(wdata[5]), .A3(n435), .A4(io_pmp_6_addr[5]), .Y(n_GEN_300[5]) );
  AO22X1_LVT U2668 ( .A1(n511), .A2(wdata[6]), .A3(n435), .A4(io_pmp_6_addr[6]), .Y(n_GEN_300[6]) );
  AO22X1_LVT U2669 ( .A1(n511), .A2(wdata[8]), .A3(n435), .A4(io_pmp_6_addr[8]), .Y(n_GEN_300[8]) );
  AO22X1_LVT U2670 ( .A1(n512), .A2(wdata[0]), .A3(n386), .A4(io_pmp_7_addr[0]), .Y(n_GEN_307[0]) );
  AO22X1_LVT U2671 ( .A1(n512), .A2(wdata[10]), .A3(n386), .A4(
        io_pmp_7_addr[10]), .Y(n_GEN_307[10]) );
  AO22X1_LVT U2672 ( .A1(n512), .A2(wdata[12]), .A3(n386), .A4(
        io_pmp_7_addr[12]), .Y(n_GEN_307[12]) );
  AO22X1_LVT U2673 ( .A1(n512), .A2(wdata[13]), .A3(n386), .A4(
        io_pmp_7_addr[13]), .Y(n_GEN_307[13]) );
  AO22X1_LVT U2674 ( .A1(n512), .A2(wdata[14]), .A3(n386), .A4(
        io_pmp_7_addr[14]), .Y(n_GEN_307[14]) );
  AO22X1_LVT U2675 ( .A1(n512), .A2(wdata[15]), .A3(n386), .A4(
        io_pmp_7_addr[15]), .Y(n_GEN_307[15]) );
  AO22X1_LVT U2676 ( .A1(n512), .A2(wdata[16]), .A3(n386), .A4(
        io_pmp_7_addr[16]), .Y(n_GEN_307[16]) );
  AO22X1_LVT U2677 ( .A1(n512), .A2(wdata[17]), .A3(n386), .A4(
        io_pmp_7_addr[17]), .Y(n_GEN_307[17]) );
  AO22X1_LVT U2678 ( .A1(n512), .A2(wdata[18]), .A3(n386), .A4(
        io_pmp_7_addr[18]), .Y(n_GEN_307[18]) );
  AO22X1_LVT U2679 ( .A1(n512), .A2(wdata[19]), .A3(n386), .A4(
        io_pmp_7_addr[19]), .Y(n_GEN_307[19]) );
  AO22X1_LVT U2680 ( .A1(n512), .A2(wdata[1]), .A3(n386), .A4(io_pmp_7_addr[1]), .Y(n_GEN_307[1]) );
  AO22X1_LVT U2681 ( .A1(n512), .A2(wdata[20]), .A3(n386), .A4(
        io_pmp_7_addr[20]), .Y(n_GEN_307[20]) );
  AO22X1_LVT U2682 ( .A1(n512), .A2(wdata[21]), .A3(n386), .A4(
        io_pmp_7_addr[21]), .Y(n_GEN_307[21]) );
  AO22X1_LVT U2683 ( .A1(n512), .A2(wdata[22]), .A3(n386), .A4(
        io_pmp_7_addr[22]), .Y(n_GEN_307[22]) );
  AO22X1_LVT U2684 ( .A1(n512), .A2(wdata[23]), .A3(n386), .A4(
        io_pmp_7_addr[23]), .Y(n_GEN_307[23]) );
  AO22X1_LVT U2685 ( .A1(n512), .A2(wdata[24]), .A3(n386), .A4(
        io_pmp_7_addr[24]), .Y(n_GEN_307[24]) );
  AO22X1_LVT U2686 ( .A1(n512), .A2(wdata[25]), .A3(n386), .A4(
        io_pmp_7_addr[25]), .Y(n_GEN_307[25]) );
  AO22X1_LVT U2687 ( .A1(n512), .A2(wdata[26]), .A3(n386), .A4(
        io_pmp_7_addr[26]), .Y(n_GEN_307[26]) );
  AO22X1_LVT U2688 ( .A1(n512), .A2(wdata[27]), .A3(n386), .A4(
        io_pmp_7_addr[27]), .Y(n_GEN_307[27]) );
  AO22X1_LVT U2689 ( .A1(n512), .A2(wdata[28]), .A3(n386), .A4(
        io_pmp_7_addr[28]), .Y(n_GEN_307[28]) );
  AO22X1_LVT U2690 ( .A1(n512), .A2(wdata[29]), .A3(n386), .A4(
        io_pmp_7_addr[29]), .Y(n_GEN_307[29]) );
  AO22X1_LVT U2691 ( .A1(n512), .A2(wdata[2]), .A3(n386), .A4(io_pmp_7_addr[2]), .Y(n_GEN_307[2]) );
  AO22X1_LVT U2692 ( .A1(n512), .A2(wdata[4]), .A3(n386), .A4(io_pmp_7_addr[4]), .Y(n_GEN_307[4]) );
  AO22X1_LVT U2693 ( .A1(n512), .A2(wdata[5]), .A3(n386), .A4(io_pmp_7_addr[5]), .Y(n_GEN_307[5]) );
  AO22X1_LVT U2694 ( .A1(n512), .A2(wdata[6]), .A3(n386), .A4(io_pmp_7_addr[6]), .Y(n_GEN_307[6]) );
  AO22X1_LVT U2695 ( .A1(n512), .A2(wdata[8]), .A3(n386), .A4(io_pmp_7_addr[8]), .Y(n_GEN_307[8]) );
  AND2X1_LVT U2696 ( .A1(n1698), .A2(io_pmp_0_addr[8]), .Y(io_pmp_0_mask[11])
         );
  AND2X1_LVT U2697 ( .A1(n1699), .A2(io_pmp_0_addr[10]), .Y(io_pmp_0_mask[13])
         );
  AND2X1_LVT U2698 ( .A1(n1700), .A2(io_pmp_0_addr[12]), .Y(io_pmp_0_mask[15])
         );
  AND2X1_LVT U2699 ( .A1(n1701), .A2(io_pmp_0_addr[13]), .Y(io_pmp_0_mask[16])
         );
  AND2X1_LVT U2700 ( .A1(n1702), .A2(io_pmp_0_addr[14]), .Y(io_pmp_0_mask[17])
         );
  AND2X1_LVT U2701 ( .A1(n1703), .A2(io_pmp_0_addr[15]), .Y(io_pmp_0_mask[18])
         );
  AND2X1_LVT U2702 ( .A1(n1704), .A2(io_pmp_0_addr[16]), .Y(io_pmp_0_mask[19])
         );
  AND2X1_LVT U2703 ( .A1(n1705), .A2(io_pmp_0_addr[17]), .Y(io_pmp_0_mask[20])
         );
  AND2X1_LVT U2704 ( .A1(n1706), .A2(io_pmp_0_addr[18]), .Y(io_pmp_0_mask[21])
         );
  AND2X1_LVT U2705 ( .A1(n1707), .A2(io_pmp_0_addr[19]), .Y(io_pmp_0_mask[22])
         );
  AND2X1_LVT U2706 ( .A1(n1708), .A2(io_pmp_0_addr[20]), .Y(io_pmp_0_mask[23])
         );
  AND2X1_LVT U2707 ( .A1(n1709), .A2(io_pmp_0_addr[21]), .Y(io_pmp_0_mask[24])
         );
  AND2X1_LVT U2708 ( .A1(n1710), .A2(io_pmp_0_addr[22]), .Y(io_pmp_0_mask[25])
         );
  AND2X1_LVT U2709 ( .A1(n1711), .A2(io_pmp_0_addr[23]), .Y(io_pmp_0_mask[26])
         );
  AND2X1_LVT U2710 ( .A1(n1712), .A2(io_pmp_0_addr[24]), .Y(io_pmp_0_mask[27])
         );
  AND2X1_LVT U2711 ( .A1(n1713), .A2(io_pmp_0_addr[25]), .Y(io_pmp_0_mask[28])
         );
  AND2X1_LVT U2712 ( .A1(n1714), .A2(io_pmp_0_addr[26]), .Y(io_pmp_0_mask[29])
         );
  AND2X1_LVT U2713 ( .A1(n1715), .A2(io_pmp_0_addr[27]), .Y(io_pmp_0_mask[30])
         );
  AND2X1_LVT U2714 ( .A1(n1716), .A2(io_pmp_0_addr[28]), .Y(io_pmp_0_mask[31])
         );
  AND2X1_LVT U2715 ( .A1(n1717), .A2(io_pmp_0_addr[0]), .Y(io_pmp_0_mask[3])
         );
  AND2X1_LVT U2716 ( .A1(n1718), .A2(io_pmp_0_addr[1]), .Y(io_pmp_0_mask[4])
         );
  AND2X1_LVT U2717 ( .A1(n1719), .A2(io_pmp_0_addr[2]), .Y(io_pmp_0_mask[5])
         );
  AND2X1_LVT U2718 ( .A1(n1720), .A2(io_pmp_0_addr[4]), .Y(io_pmp_0_mask[7])
         );
  AND2X1_LVT U2719 ( .A1(n1721), .A2(io_pmp_0_addr[5]), .Y(io_pmp_0_mask[8])
         );
  AND2X1_LVT U2720 ( .A1(n1722), .A2(io_pmp_0_addr[6]), .Y(io_pmp_0_mask[9])
         );
  AND2X1_LVT U2721 ( .A1(n1723), .A2(io_pmp_1_addr[8]), .Y(io_pmp_1_mask[11])
         );
  AND2X1_LVT U2722 ( .A1(n1724), .A2(io_pmp_1_addr[10]), .Y(io_pmp_1_mask[13])
         );
  AND2X1_LVT U2723 ( .A1(n1725), .A2(io_pmp_1_addr[12]), .Y(io_pmp_1_mask[15])
         );
  AND2X1_LVT U2724 ( .A1(n1726), .A2(io_pmp_1_addr[13]), .Y(io_pmp_1_mask[16])
         );
  AND2X1_LVT U2725 ( .A1(n1727), .A2(io_pmp_1_addr[14]), .Y(io_pmp_1_mask[17])
         );
  AND2X1_LVT U2726 ( .A1(n1728), .A2(io_pmp_1_addr[15]), .Y(io_pmp_1_mask[18])
         );
  AND2X1_LVT U2727 ( .A1(n1729), .A2(io_pmp_1_addr[16]), .Y(io_pmp_1_mask[19])
         );
  AND2X1_LVT U2728 ( .A1(n1730), .A2(io_pmp_1_addr[17]), .Y(io_pmp_1_mask[20])
         );
  AND2X1_LVT U2729 ( .A1(n1731), .A2(io_pmp_1_addr[18]), .Y(io_pmp_1_mask[21])
         );
  AND2X1_LVT U2730 ( .A1(n1732), .A2(io_pmp_1_addr[19]), .Y(io_pmp_1_mask[22])
         );
  AND2X1_LVT U2731 ( .A1(n1733), .A2(io_pmp_1_addr[20]), .Y(io_pmp_1_mask[23])
         );
  AND2X1_LVT U2732 ( .A1(n1734), .A2(io_pmp_1_addr[21]), .Y(io_pmp_1_mask[24])
         );
  AND2X1_LVT U2733 ( .A1(n1735), .A2(io_pmp_1_addr[22]), .Y(io_pmp_1_mask[25])
         );
  AND2X1_LVT U2734 ( .A1(n1736), .A2(io_pmp_1_addr[23]), .Y(io_pmp_1_mask[26])
         );
  AND2X1_LVT U2735 ( .A1(n1737), .A2(io_pmp_1_addr[24]), .Y(io_pmp_1_mask[27])
         );
  AND2X1_LVT U2736 ( .A1(n1738), .A2(io_pmp_1_addr[25]), .Y(io_pmp_1_mask[28])
         );
  AND2X1_LVT U2737 ( .A1(n1739), .A2(io_pmp_1_addr[26]), .Y(io_pmp_1_mask[29])
         );
  AND2X1_LVT U2738 ( .A1(n1740), .A2(io_pmp_1_addr[27]), .Y(io_pmp_1_mask[30])
         );
  AND2X1_LVT U2739 ( .A1(n1741), .A2(io_pmp_1_addr[28]), .Y(io_pmp_1_mask[31])
         );
  AND2X1_LVT U2740 ( .A1(n1742), .A2(io_pmp_1_addr[0]), .Y(io_pmp_1_mask[3])
         );
  AND2X1_LVT U2741 ( .A1(n1743), .A2(io_pmp_1_addr[1]), .Y(io_pmp_1_mask[4])
         );
  AND2X1_LVT U2742 ( .A1(n1744), .A2(io_pmp_1_addr[2]), .Y(io_pmp_1_mask[5])
         );
  AND2X1_LVT U2743 ( .A1(n1745), .A2(io_pmp_1_addr[4]), .Y(io_pmp_1_mask[7])
         );
  AND2X1_LVT U2744 ( .A1(n1746), .A2(io_pmp_1_addr[5]), .Y(io_pmp_1_mask[8])
         );
  AND2X1_LVT U2745 ( .A1(n1747), .A2(io_pmp_1_addr[6]), .Y(io_pmp_1_mask[9])
         );
  AND2X1_LVT U2746 ( .A1(n1748), .A2(io_pmp_2_addr[8]), .Y(io_pmp_2_mask[11])
         );
  AND2X1_LVT U2747 ( .A1(n1749), .A2(io_pmp_2_addr[10]), .Y(io_pmp_2_mask[13])
         );
  AND2X1_LVT U2748 ( .A1(n1750), .A2(io_pmp_2_addr[12]), .Y(io_pmp_2_mask[15])
         );
  AND2X1_LVT U2749 ( .A1(n1751), .A2(io_pmp_2_addr[13]), .Y(io_pmp_2_mask[16])
         );
  AND2X1_LVT U2750 ( .A1(n1752), .A2(io_pmp_2_addr[14]), .Y(io_pmp_2_mask[17])
         );
  AND2X1_LVT U2751 ( .A1(n1753), .A2(io_pmp_2_addr[15]), .Y(io_pmp_2_mask[18])
         );
  AND2X1_LVT U2752 ( .A1(n1754), .A2(io_pmp_2_addr[16]), .Y(io_pmp_2_mask[19])
         );
  AND2X1_LVT U2753 ( .A1(n1755), .A2(io_pmp_2_addr[17]), .Y(io_pmp_2_mask[20])
         );
  AND2X1_LVT U2754 ( .A1(n1756), .A2(io_pmp_2_addr[18]), .Y(io_pmp_2_mask[21])
         );
  AND2X1_LVT U2755 ( .A1(n1757), .A2(io_pmp_2_addr[19]), .Y(io_pmp_2_mask[22])
         );
  AND2X1_LVT U2756 ( .A1(n1758), .A2(io_pmp_2_addr[20]), .Y(io_pmp_2_mask[23])
         );
  AND2X1_LVT U2757 ( .A1(n1759), .A2(io_pmp_2_addr[21]), .Y(io_pmp_2_mask[24])
         );
  AND2X1_LVT U2758 ( .A1(n1760), .A2(io_pmp_2_addr[22]), .Y(io_pmp_2_mask[25])
         );
  AND2X1_LVT U2759 ( .A1(n1761), .A2(io_pmp_2_addr[23]), .Y(io_pmp_2_mask[26])
         );
  AND2X1_LVT U2760 ( .A1(n1762), .A2(io_pmp_2_addr[24]), .Y(io_pmp_2_mask[27])
         );
  AND2X1_LVT U2761 ( .A1(n1763), .A2(io_pmp_2_addr[25]), .Y(io_pmp_2_mask[28])
         );
  AND2X1_LVT U2762 ( .A1(n1764), .A2(io_pmp_2_addr[26]), .Y(io_pmp_2_mask[29])
         );
  AND2X1_LVT U2763 ( .A1(n1765), .A2(io_pmp_2_addr[27]), .Y(io_pmp_2_mask[30])
         );
  AND2X1_LVT U2764 ( .A1(n1766), .A2(io_pmp_2_addr[28]), .Y(io_pmp_2_mask[31])
         );
  AND2X1_LVT U2765 ( .A1(n1767), .A2(io_pmp_2_addr[0]), .Y(io_pmp_2_mask[3])
         );
  AND2X1_LVT U2766 ( .A1(n1768), .A2(io_pmp_2_addr[1]), .Y(io_pmp_2_mask[4])
         );
  AND2X1_LVT U2767 ( .A1(n1769), .A2(io_pmp_2_addr[2]), .Y(io_pmp_2_mask[5])
         );
  AND2X1_LVT U2768 ( .A1(n1770), .A2(io_pmp_2_addr[4]), .Y(io_pmp_2_mask[7])
         );
  AND2X1_LVT U2769 ( .A1(n1771), .A2(io_pmp_2_addr[5]), .Y(io_pmp_2_mask[8])
         );
  AND2X1_LVT U2770 ( .A1(n1772), .A2(io_pmp_2_addr[6]), .Y(io_pmp_2_mask[9])
         );
  AND2X1_LVT U2771 ( .A1(n1773), .A2(io_pmp_3_addr[8]), .Y(io_pmp_3_mask[11])
         );
  AND2X1_LVT U2772 ( .A1(n1774), .A2(io_pmp_3_addr[10]), .Y(io_pmp_3_mask[13])
         );
  AND2X1_LVT U2773 ( .A1(n1775), .A2(io_pmp_3_addr[12]), .Y(io_pmp_3_mask[15])
         );
  AND2X1_LVT U2774 ( .A1(n1776), .A2(io_pmp_3_addr[13]), .Y(io_pmp_3_mask[16])
         );
  AND2X1_LVT U2775 ( .A1(n1777), .A2(io_pmp_3_addr[14]), .Y(io_pmp_3_mask[17])
         );
  AND2X1_LVT U2776 ( .A1(n1778), .A2(io_pmp_3_addr[15]), .Y(io_pmp_3_mask[18])
         );
  AND2X1_LVT U2777 ( .A1(n1779), .A2(io_pmp_3_addr[16]), .Y(io_pmp_3_mask[19])
         );
  AND2X1_LVT U2778 ( .A1(n1780), .A2(io_pmp_3_addr[17]), .Y(io_pmp_3_mask[20])
         );
  AND2X1_LVT U2779 ( .A1(n1781), .A2(io_pmp_3_addr[18]), .Y(io_pmp_3_mask[21])
         );
  AND2X1_LVT U2780 ( .A1(n1782), .A2(io_pmp_3_addr[19]), .Y(io_pmp_3_mask[22])
         );
  AND2X1_LVT U2781 ( .A1(n1783), .A2(io_pmp_3_addr[20]), .Y(io_pmp_3_mask[23])
         );
  AND2X1_LVT U2782 ( .A1(n1784), .A2(io_pmp_3_addr[21]), .Y(io_pmp_3_mask[24])
         );
  AND2X1_LVT U2783 ( .A1(n1785), .A2(io_pmp_3_addr[22]), .Y(io_pmp_3_mask[25])
         );
  AND2X1_LVT U2784 ( .A1(n1786), .A2(io_pmp_3_addr[23]), .Y(io_pmp_3_mask[26])
         );
  AND2X1_LVT U2785 ( .A1(n1787), .A2(io_pmp_3_addr[24]), .Y(io_pmp_3_mask[27])
         );
  AND2X1_LVT U2786 ( .A1(n1788), .A2(io_pmp_3_addr[25]), .Y(io_pmp_3_mask[28])
         );
  AND2X1_LVT U2787 ( .A1(n1789), .A2(io_pmp_3_addr[26]), .Y(io_pmp_3_mask[29])
         );
  AND2X1_LVT U2788 ( .A1(n1790), .A2(io_pmp_3_addr[27]), .Y(io_pmp_3_mask[30])
         );
  AND2X1_LVT U2789 ( .A1(n1791), .A2(io_pmp_3_addr[28]), .Y(io_pmp_3_mask[31])
         );
  AND2X1_LVT U2790 ( .A1(n1792), .A2(io_pmp_3_addr[0]), .Y(io_pmp_3_mask[3])
         );
  AND2X1_LVT U2791 ( .A1(n1793), .A2(io_pmp_3_addr[1]), .Y(io_pmp_3_mask[4])
         );
  AND2X1_LVT U2792 ( .A1(n1794), .A2(io_pmp_3_addr[2]), .Y(io_pmp_3_mask[5])
         );
  AND2X1_LVT U2793 ( .A1(n1795), .A2(io_pmp_3_addr[4]), .Y(io_pmp_3_mask[7])
         );
  AND2X1_LVT U2794 ( .A1(n1796), .A2(io_pmp_3_addr[5]), .Y(io_pmp_3_mask[8])
         );
  AND2X1_LVT U2795 ( .A1(n1797), .A2(io_pmp_3_addr[6]), .Y(io_pmp_3_mask[9])
         );
  AND2X1_LVT U2796 ( .A1(n1798), .A2(io_pmp_4_addr[8]), .Y(io_pmp_4_mask[11])
         );
  AND2X1_LVT U2797 ( .A1(n1799), .A2(io_pmp_4_addr[10]), .Y(io_pmp_4_mask[13])
         );
  AND2X1_LVT U2798 ( .A1(n1800), .A2(io_pmp_4_addr[12]), .Y(io_pmp_4_mask[15])
         );
  AND2X1_LVT U2799 ( .A1(n1801), .A2(io_pmp_4_addr[13]), .Y(io_pmp_4_mask[16])
         );
  AND2X1_LVT U2800 ( .A1(n1802), .A2(io_pmp_4_addr[14]), .Y(io_pmp_4_mask[17])
         );
  AND2X1_LVT U2801 ( .A1(n1803), .A2(io_pmp_4_addr[15]), .Y(io_pmp_4_mask[18])
         );
  AND2X1_LVT U2802 ( .A1(n1804), .A2(io_pmp_4_addr[16]), .Y(io_pmp_4_mask[19])
         );
  AND2X1_LVT U2803 ( .A1(n1805), .A2(io_pmp_4_addr[17]), .Y(io_pmp_4_mask[20])
         );
  AND2X1_LVT U2804 ( .A1(n1806), .A2(io_pmp_4_addr[18]), .Y(io_pmp_4_mask[21])
         );
  AND2X1_LVT U2805 ( .A1(n1807), .A2(io_pmp_4_addr[19]), .Y(io_pmp_4_mask[22])
         );
  AND2X1_LVT U2806 ( .A1(n1808), .A2(io_pmp_4_addr[20]), .Y(io_pmp_4_mask[23])
         );
  AND2X1_LVT U2807 ( .A1(n1809), .A2(io_pmp_4_addr[21]), .Y(io_pmp_4_mask[24])
         );
  AND2X1_LVT U2808 ( .A1(n1810), .A2(io_pmp_4_addr[22]), .Y(io_pmp_4_mask[25])
         );
  AND2X1_LVT U2809 ( .A1(n1811), .A2(io_pmp_4_addr[23]), .Y(io_pmp_4_mask[26])
         );
  AND2X1_LVT U2810 ( .A1(n1812), .A2(io_pmp_4_addr[24]), .Y(io_pmp_4_mask[27])
         );
  AND2X1_LVT U2811 ( .A1(n1813), .A2(io_pmp_4_addr[25]), .Y(io_pmp_4_mask[28])
         );
  AND2X1_LVT U2812 ( .A1(n1814), .A2(io_pmp_4_addr[26]), .Y(io_pmp_4_mask[29])
         );
  AND2X1_LVT U2813 ( .A1(n1815), .A2(io_pmp_4_addr[27]), .Y(io_pmp_4_mask[30])
         );
  AND2X1_LVT U2814 ( .A1(n1816), .A2(io_pmp_4_addr[28]), .Y(io_pmp_4_mask[31])
         );
  AND2X1_LVT U2815 ( .A1(n1817), .A2(io_pmp_4_addr[0]), .Y(io_pmp_4_mask[3])
         );
  AND2X1_LVT U2816 ( .A1(n1818), .A2(io_pmp_4_addr[1]), .Y(io_pmp_4_mask[4])
         );
  AND2X1_LVT U2817 ( .A1(n1819), .A2(io_pmp_4_addr[2]), .Y(io_pmp_4_mask[5])
         );
  AND2X1_LVT U2818 ( .A1(n1820), .A2(io_pmp_4_addr[4]), .Y(io_pmp_4_mask[7])
         );
  AND2X1_LVT U2819 ( .A1(n1821), .A2(io_pmp_4_addr[5]), .Y(io_pmp_4_mask[8])
         );
  AND2X1_LVT U2820 ( .A1(n1822), .A2(io_pmp_4_addr[6]), .Y(io_pmp_4_mask[9])
         );
  AND2X1_LVT U2821 ( .A1(n1823), .A2(io_pmp_5_addr[8]), .Y(io_pmp_5_mask[11])
         );
  AND2X1_LVT U2822 ( .A1(n1824), .A2(io_pmp_5_addr[10]), .Y(io_pmp_5_mask[13])
         );
  AND2X1_LVT U2823 ( .A1(n1825), .A2(io_pmp_5_addr[12]), .Y(io_pmp_5_mask[15])
         );
  AND2X1_LVT U2824 ( .A1(n1826), .A2(io_pmp_5_addr[13]), .Y(io_pmp_5_mask[16])
         );
  AND2X1_LVT U2825 ( .A1(n1827), .A2(io_pmp_5_addr[14]), .Y(io_pmp_5_mask[17])
         );
  AND2X1_LVT U2826 ( .A1(n1828), .A2(io_pmp_5_addr[15]), .Y(io_pmp_5_mask[18])
         );
  AND2X1_LVT U2827 ( .A1(n1829), .A2(io_pmp_5_addr[16]), .Y(io_pmp_5_mask[19])
         );
  AND2X1_LVT U2828 ( .A1(n1830), .A2(io_pmp_5_addr[17]), .Y(io_pmp_5_mask[20])
         );
  AND2X1_LVT U2829 ( .A1(n1831), .A2(io_pmp_5_addr[18]), .Y(io_pmp_5_mask[21])
         );
  AND2X1_LVT U2830 ( .A1(n1832), .A2(io_pmp_5_addr[19]), .Y(io_pmp_5_mask[22])
         );
  AND2X1_LVT U2831 ( .A1(n1833), .A2(io_pmp_5_addr[20]), .Y(io_pmp_5_mask[23])
         );
  AND2X1_LVT U2832 ( .A1(n1834), .A2(io_pmp_5_addr[21]), .Y(io_pmp_5_mask[24])
         );
  AND2X1_LVT U2833 ( .A1(n1835), .A2(io_pmp_5_addr[22]), .Y(io_pmp_5_mask[25])
         );
  AND2X1_LVT U2834 ( .A1(n1836), .A2(io_pmp_5_addr[23]), .Y(io_pmp_5_mask[26])
         );
  AND2X1_LVT U2835 ( .A1(n1837), .A2(io_pmp_5_addr[24]), .Y(io_pmp_5_mask[27])
         );
  AND2X1_LVT U2836 ( .A1(n1838), .A2(io_pmp_5_addr[25]), .Y(io_pmp_5_mask[28])
         );
  AND2X1_LVT U2837 ( .A1(n1839), .A2(io_pmp_5_addr[26]), .Y(io_pmp_5_mask[29])
         );
  AND2X1_LVT U2838 ( .A1(n1840), .A2(io_pmp_5_addr[27]), .Y(io_pmp_5_mask[30])
         );
  AND2X1_LVT U2839 ( .A1(n1841), .A2(io_pmp_5_addr[28]), .Y(io_pmp_5_mask[31])
         );
  AND2X1_LVT U2840 ( .A1(n1842), .A2(io_pmp_5_addr[0]), .Y(io_pmp_5_mask[3])
         );
  AND2X1_LVT U2841 ( .A1(n1843), .A2(io_pmp_5_addr[1]), .Y(io_pmp_5_mask[4])
         );
  AND2X1_LVT U2842 ( .A1(n1844), .A2(io_pmp_5_addr[2]), .Y(io_pmp_5_mask[5])
         );
  AND2X1_LVT U2843 ( .A1(n1845), .A2(io_pmp_5_addr[4]), .Y(io_pmp_5_mask[7])
         );
  AND2X1_LVT U2844 ( .A1(n1846), .A2(io_pmp_5_addr[5]), .Y(io_pmp_5_mask[8])
         );
  AND2X1_LVT U2845 ( .A1(n1847), .A2(io_pmp_5_addr[6]), .Y(io_pmp_5_mask[9])
         );
  AND2X1_LVT U2846 ( .A1(n1848), .A2(io_pmp_6_addr[8]), .Y(io_pmp_6_mask[11])
         );
  AND2X1_LVT U2847 ( .A1(n1849), .A2(io_pmp_6_addr[10]), .Y(io_pmp_6_mask[13])
         );
  AND2X1_LVT U2848 ( .A1(n1850), .A2(io_pmp_6_addr[12]), .Y(io_pmp_6_mask[15])
         );
  AND2X1_LVT U2849 ( .A1(n1851), .A2(io_pmp_6_addr[13]), .Y(io_pmp_6_mask[16])
         );
  AND2X1_LVT U2850 ( .A1(n1852), .A2(io_pmp_6_addr[14]), .Y(io_pmp_6_mask[17])
         );
  AND2X1_LVT U2851 ( .A1(n1853), .A2(io_pmp_6_addr[15]), .Y(io_pmp_6_mask[18])
         );
  AND2X1_LVT U2852 ( .A1(n1854), .A2(io_pmp_6_addr[16]), .Y(io_pmp_6_mask[19])
         );
  AND2X1_LVT U2853 ( .A1(n1855), .A2(io_pmp_6_addr[17]), .Y(io_pmp_6_mask[20])
         );
  AND2X1_LVT U2854 ( .A1(n1856), .A2(io_pmp_6_addr[18]), .Y(io_pmp_6_mask[21])
         );
  AND2X1_LVT U2855 ( .A1(n1857), .A2(io_pmp_6_addr[19]), .Y(io_pmp_6_mask[22])
         );
  AND2X1_LVT U2856 ( .A1(n1858), .A2(io_pmp_6_addr[20]), .Y(io_pmp_6_mask[23])
         );
  AND2X1_LVT U2857 ( .A1(n1859), .A2(io_pmp_6_addr[21]), .Y(io_pmp_6_mask[24])
         );
  AND2X1_LVT U2858 ( .A1(n1860), .A2(io_pmp_6_addr[22]), .Y(io_pmp_6_mask[25])
         );
  AND2X1_LVT U2859 ( .A1(n1861), .A2(io_pmp_6_addr[23]), .Y(io_pmp_6_mask[26])
         );
  AND2X1_LVT U2860 ( .A1(n1862), .A2(io_pmp_6_addr[24]), .Y(io_pmp_6_mask[27])
         );
  AND2X1_LVT U2861 ( .A1(n1863), .A2(io_pmp_6_addr[25]), .Y(io_pmp_6_mask[28])
         );
  AND2X1_LVT U2862 ( .A1(n1864), .A2(io_pmp_6_addr[26]), .Y(io_pmp_6_mask[29])
         );
  AND2X1_LVT U2863 ( .A1(n1865), .A2(io_pmp_6_addr[27]), .Y(io_pmp_6_mask[30])
         );
  AND2X1_LVT U2864 ( .A1(n1866), .A2(io_pmp_6_addr[28]), .Y(io_pmp_6_mask[31])
         );
  AND2X1_LVT U2865 ( .A1(n1867), .A2(io_pmp_6_addr[0]), .Y(io_pmp_6_mask[3])
         );
  AND2X1_LVT U2866 ( .A1(n1868), .A2(io_pmp_6_addr[1]), .Y(io_pmp_6_mask[4])
         );
  AND2X1_LVT U2867 ( .A1(n1869), .A2(io_pmp_6_addr[2]), .Y(io_pmp_6_mask[5])
         );
  AND2X1_LVT U2868 ( .A1(n1870), .A2(io_pmp_6_addr[4]), .Y(io_pmp_6_mask[7])
         );
  AND2X1_LVT U2869 ( .A1(n1871), .A2(io_pmp_6_addr[5]), .Y(io_pmp_6_mask[8])
         );
  AND2X1_LVT U2870 ( .A1(n1872), .A2(io_pmp_6_addr[6]), .Y(io_pmp_6_mask[9])
         );
  AND2X1_LVT U2871 ( .A1(n1873), .A2(io_pmp_7_addr[8]), .Y(io_pmp_7_mask[11])
         );
  AND2X1_LVT U2872 ( .A1(n1874), .A2(io_pmp_7_addr[10]), .Y(io_pmp_7_mask[13])
         );
  AND2X1_LVT U2873 ( .A1(n1875), .A2(io_pmp_7_addr[12]), .Y(io_pmp_7_mask[15])
         );
  AND2X1_LVT U2874 ( .A1(n1876), .A2(io_pmp_7_addr[13]), .Y(io_pmp_7_mask[16])
         );
  AND2X1_LVT U2875 ( .A1(n1877), .A2(io_pmp_7_addr[14]), .Y(io_pmp_7_mask[17])
         );
  AND2X1_LVT U2876 ( .A1(n1878), .A2(io_pmp_7_addr[15]), .Y(io_pmp_7_mask[18])
         );
  AND2X1_LVT U2877 ( .A1(n1879), .A2(io_pmp_7_addr[16]), .Y(io_pmp_7_mask[19])
         );
  AND2X1_LVT U2878 ( .A1(n1880), .A2(io_pmp_7_addr[17]), .Y(io_pmp_7_mask[20])
         );
  AND2X1_LVT U2879 ( .A1(n1881), .A2(io_pmp_7_addr[18]), .Y(io_pmp_7_mask[21])
         );
  AND2X1_LVT U2880 ( .A1(n1882), .A2(io_pmp_7_addr[19]), .Y(io_pmp_7_mask[22])
         );
  AND2X1_LVT U2881 ( .A1(n1883), .A2(io_pmp_7_addr[20]), .Y(io_pmp_7_mask[23])
         );
  AND2X1_LVT U2882 ( .A1(n1884), .A2(io_pmp_7_addr[21]), .Y(io_pmp_7_mask[24])
         );
  AND2X1_LVT U2883 ( .A1(n1885), .A2(io_pmp_7_addr[22]), .Y(io_pmp_7_mask[25])
         );
  AND2X1_LVT U2884 ( .A1(n1886), .A2(io_pmp_7_addr[23]), .Y(io_pmp_7_mask[26])
         );
  AND2X1_LVT U2885 ( .A1(n1887), .A2(io_pmp_7_addr[24]), .Y(io_pmp_7_mask[27])
         );
  AND2X1_LVT U2886 ( .A1(n1888), .A2(io_pmp_7_addr[25]), .Y(io_pmp_7_mask[28])
         );
  AND2X1_LVT U2887 ( .A1(n1889), .A2(io_pmp_7_addr[26]), .Y(io_pmp_7_mask[29])
         );
  AND2X1_LVT U2888 ( .A1(n1890), .A2(io_pmp_7_addr[27]), .Y(io_pmp_7_mask[30])
         );
  AND2X1_LVT U2889 ( .A1(n1891), .A2(io_pmp_7_addr[28]), .Y(io_pmp_7_mask[31])
         );
  AND2X1_LVT U2890 ( .A1(n1892), .A2(io_pmp_7_addr[0]), .Y(io_pmp_7_mask[3])
         );
  AND2X1_LVT U2891 ( .A1(n1893), .A2(io_pmp_7_addr[1]), .Y(io_pmp_7_mask[4])
         );
  AND2X1_LVT U2892 ( .A1(n1894), .A2(io_pmp_7_addr[2]), .Y(io_pmp_7_mask[5])
         );
  AND2X1_LVT U2893 ( .A1(n1895), .A2(io_pmp_7_addr[4]), .Y(io_pmp_7_mask[7])
         );
  AND2X1_LVT U2894 ( .A1(n1896), .A2(io_pmp_7_addr[5]), .Y(io_pmp_7_mask[8])
         );
  AND2X1_LVT U2895 ( .A1(n1897), .A2(io_pmp_7_addr[6]), .Y(io_pmp_7_mask[9])
         );
  AO22X1_LVT U2896 ( .A1(n513), .A2(wdata[1]), .A3(n448), .A4(io_pc[1]), .Y(
        net34877) );
  AO22X1_LVT U2897 ( .A1(n514), .A2(wdata[1]), .A3(n449), .A4(io_pc[1]), .Y(
        net35079) );
  AO22X1_LVT U2898 ( .A1(n515), .A2(wdata[1]), .A3(n450), .A4(io_pc[1]), .Y(
        net35301) );
  AND2X1_LVT U2899 ( .A1(n504), .A2(n1484), .Y(n2169) );
  AND2X1_LVT U2900 ( .A1(n504), .A2(n1465), .Y(n2168) );
  AND2X1_LVT U2901 ( .A1(n1487), .A2(n504), .Y(n2167) );
  AND3X1_LVT U2902 ( .A1(io_rw_addr[1]), .A2(n504), .A3(n1486), .Y(n2166) );
  AO221X1_LVT U2903 ( .A1(n1899), .A2(n407), .A3(n1899), .A4(n1898), .A5(n1476), .Y(n1902) );
  OA21X1_LVT U2904 ( .A1(n1474), .A2(n1475), .A3(read_mideleg_1), .Y(n1901) );
  AND2X1_LVT U2905 ( .A1(io_rw_wdata[1]), .A2(n516), .Y(n1900) );
  NAND2X0_LVT U2906 ( .A1(n589), .A2(n1904), .Y(n1905) );
  NAND2X0_LVT U2907 ( .A1(n1474), .A2(n1905), .Y(n1906) );
  NAND2X0_LVT U2908 ( .A1(n589), .A2(n1907), .Y(n1908) );
endmodule


module BreakpointUnit_DW_cmp_J40_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [38:0] A;
  input [38:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422;

  AO221X1_LVT U201 ( .A1(1'b1), .A2(n400), .A3(B[11]), .A4(n330), .A5(n331), 
        .Y(n397) );
  AO221X1_LVT U202 ( .A1(1'b1), .A2(n406), .A3(B[19]), .A4(n320), .A5(n321), 
        .Y(n388) );
  OA221X1_LVT U203 ( .A1(1'b0), .A2(n382), .A3(A[27]), .A4(n295), .A5(n296), 
        .Y(n380) );
  INVX0_LVT U204 ( .A(A[29]), .Y(n284) );
  AO22X1_LVT U205 ( .A1(B[29]), .A2(n284), .A3(B[30]), .A4(n348), .Y(n371) );
  INVX0_LVT U206 ( .A(A[0]), .Y(n285) );
  INVX0_LVT U207 ( .A(A[2]), .Y(n286) );
  INVX0_LVT U208 ( .A(A[1]), .Y(n287) );
  AO222X1_LVT U209 ( .A1(n285), .A2(B[0]), .A3(n286), .A4(B[2]), .A5(n287), 
        .A6(B[1]), .Y(n288) );
  NAND2X0_LVT U210 ( .A1(B[2]), .A2(n286), .Y(n289) );
  NAND2X0_LVT U211 ( .A1(A[1]), .A2(n289), .Y(n290) );
  OA22X1_LVT U212 ( .A1(B[2]), .A2(n286), .A3(B[1]), .A4(n290), .Y(n291) );
  INVX0_LVT U213 ( .A(A[3]), .Y(n292) );
  NAND2X0_LVT U214 ( .A1(B[3]), .A2(n292), .Y(n293) );
  NAND2X0_LVT U215 ( .A1(n291), .A2(n288), .Y(n294) );
  NAND3X0_LVT U216 ( .A1(n294), .A2(n395), .A3(n293), .Y(n391) );
  INVX0_LVT U217 ( .A(B[27]), .Y(n295) );
  INVX0_LVT U218 ( .A(n371), .Y(n296) );
  NAND2X0_LVT U220 ( .A1(n350), .A2(B[26]), .Y(n298) );
  NAND2X0_LVT U221 ( .A1(A[25]), .A2(n298), .Y(n299) );
  OA22X1_LVT U222 ( .A1(n350), .A2(B[26]), .A3(B[25]), .A4(n299), .Y(n376) );
  NAND2X0_LVT U223 ( .A1(n355), .A2(B[18]), .Y(n300) );
  NAND2X0_LVT U224 ( .A1(A[17]), .A2(n300), .Y(n301) );
  OA22X1_LVT U225 ( .A1(n355), .A2(B[18]), .A3(B[17]), .A4(n301), .Y(n411) );
  INVX0_LVT U226 ( .A(A[25]), .Y(n302) );
  AO22X1_LVT U227 ( .A1(B[25]), .A2(n302), .A3(B[26]), .A4(n350), .Y(n378) );
  INVX0_LVT U228 ( .A(A[17]), .Y(n303) );
  AO22X1_LVT U229 ( .A1(n355), .A2(B[18]), .A3(B[17]), .A4(n303), .Y(n387) );
  NAND2X0_LVT U230 ( .A1(n361), .A2(B[6]), .Y(n304) );
  NAND2X0_LVT U231 ( .A1(A[5]), .A2(n304), .Y(n305) );
  OA22X1_LVT U232 ( .A1(n361), .A2(B[6]), .A3(B[5]), .A4(n305), .Y(n394) );
  NAND2X0_LVT U233 ( .A1(n345), .A2(B[34]), .Y(n306) );
  NAND2X0_LVT U234 ( .A1(A[33]), .A2(n306), .Y(n307) );
  OA22X1_LVT U235 ( .A1(n345), .A2(B[34]), .A3(B[33]), .A4(n307), .Y(n421) );
  INVX0_LVT U236 ( .A(A[21]), .Y(n308) );
  AO22X1_LVT U237 ( .A1(n353), .A2(B[22]), .A3(B[21]), .A4(n308), .Y(n406) );
  NAND2X0_LVT U238 ( .A1(n359), .A2(B[10]), .Y(n309) );
  NAND2X0_LVT U239 ( .A1(A[9]), .A2(n309), .Y(n310) );
  NAND2X0_LVT U240 ( .A1(n399), .A2(A[7]), .Y(n311) );
  OA22X1_LVT U241 ( .A1(B[8]), .A2(n360), .A3(B[7]), .A4(n311), .Y(n312) );
  OA222X1_LVT U242 ( .A1(n310), .A2(B[9]), .A3(n359), .A4(B[10]), .A5(n396), 
        .A6(n312), .Y(n402) );
  INVX0_LVT U243 ( .A(A[13]), .Y(n313) );
  AO22X1_LVT U244 ( .A1(n357), .A2(B[14]), .A3(B[13]), .A4(n313), .Y(n400) );
  NAND2X0_LVT U245 ( .A1(n404), .A2(A[11]), .Y(n314) );
  OA22X1_LVT U246 ( .A1(B[12]), .A2(n358), .A3(B[11]), .A4(n314), .Y(n401) );
  NAND2X0_LVT U247 ( .A1(n346), .A2(B[32]), .Y(n315) );
  NAND2X0_LVT U248 ( .A1(A[31]), .A2(n315), .Y(n316) );
  OA22X1_LVT U249 ( .A1(n346), .A2(B[32]), .A3(B[31]), .A4(n316), .Y(n422) );
  INVX0_LVT U250 ( .A(A[33]), .Y(n317) );
  AO22X1_LVT U251 ( .A1(B[33]), .A2(n317), .A3(B[34]), .A4(n345), .Y(n416) );
  NAND2X0_LVT U252 ( .A1(n395), .A2(A[3]), .Y(n318) );
  OA22X1_LVT U253 ( .A1(B[4]), .A2(n362), .A3(B[3]), .A4(n318), .Y(n393) );
  INVX0_LVT U255 ( .A(A[19]), .Y(n320) );
  INVX0_LVT U256 ( .A(n413), .Y(n321) );
  NAND2X0_LVT U257 ( .A1(n390), .A2(A[15]), .Y(n322) );
  OA22X1_LVT U258 ( .A1(B[16]), .A2(n356), .A3(B[15]), .A4(n322), .Y(n412) );
  NAND2X0_LVT U259 ( .A1(n357), .A2(B[14]), .Y(n323) );
  NAND2X0_LVT U260 ( .A1(A[13]), .A2(n323), .Y(n324) );
  OA22X1_LVT U261 ( .A1(n357), .A2(B[14]), .A3(B[13]), .A4(n324), .Y(n403) );
  INVX0_LVT U262 ( .A(A[9]), .Y(n325) );
  AO22X1_LVT U263 ( .A1(n359), .A2(B[10]), .A3(B[9]), .A4(n325), .Y(n396) );
  NAND2X0_LVT U264 ( .A1(n379), .A2(A[23]), .Y(n326) );
  OA22X1_LVT U265 ( .A1(B[24]), .A2(n351), .A3(B[23]), .A4(n326), .Y(n377) );
  NAND2X0_LVT U266 ( .A1(n348), .A2(B[30]), .Y(n327) );
  NAND2X0_LVT U267 ( .A1(A[29]), .A2(n327), .Y(n375) );
  NAND2X0_LVT U268 ( .A1(n353), .A2(B[22]), .Y(n328) );
  NAND2X0_LVT U269 ( .A1(A[21]), .A2(n328), .Y(n410) );
  INVX0_LVT U270 ( .A(A[5]), .Y(n329) );
  AO22X1_LVT U271 ( .A1(n361), .A2(B[6]), .A3(B[5]), .A4(n329), .Y(n392) );
  INVX0_LVT U272 ( .A(A[11]), .Y(n330) );
  INVX0_LVT U273 ( .A(n404), .Y(n331) );
  INVX1_LVT U275 ( .A(A[14]), .Y(n357) );
  INVX1_LVT U276 ( .A(A[4]), .Y(n362) );
  INVX1_LVT U277 ( .A(A[34]), .Y(n345) );
  INVX1_LVT U278 ( .A(A[32]), .Y(n346) );
  INVX1_LVT U279 ( .A(A[31]), .Y(n347) );
  INVX1_LVT U280 ( .A(A[12]), .Y(n358) );
  INVX1_LVT U281 ( .A(A[36]), .Y(n343) );
  INVX1_LVT U282 ( .A(A[10]), .Y(n359) );
  INVX1_LVT U283 ( .A(A[35]), .Y(n344) );
  INVX1_LVT U284 ( .A(A[8]), .Y(n360) );
  INVX1_LVT U285 ( .A(B[7]), .Y(n342) );
  INVX1_LVT U286 ( .A(B[15]), .Y(n341) );
  INVX1_LVT U287 ( .A(A[16]), .Y(n356) );
  INVX1_LVT U288 ( .A(A[23]), .Y(n352) );
  INVX1_LVT U289 ( .A(A[24]), .Y(n351) );
  INVX1_LVT U290 ( .A(A[6]), .Y(n361) );
  INVX1_LVT U291 ( .A(A[18]), .Y(n355) );
  INVX1_LVT U292 ( .A(A[22]), .Y(n353) );
  INVX1_LVT U293 ( .A(A[20]), .Y(n354) );
  INVX1_LVT U294 ( .A(A[26]), .Y(n350) );
  INVX1_LVT U295 ( .A(A[28]), .Y(n349) );
  INVX1_LVT U296 ( .A(A[30]), .Y(n348) );
  INVX0_LVT U297 ( .A(n380), .Y(n336) );
  INVX0_LVT U298 ( .A(n416), .Y(n339) );
  OAI21X1_LVT U299 ( .A1(A[15]), .A2(n341), .A3(n390), .Y(n389) );
  OAI21X1_LVT U300 ( .A1(A[7]), .A2(n342), .A3(n399), .Y(n398) );
  OA221X1_LVT U301 ( .A1(n373), .A2(n336), .A3(n372), .A4(n371), .A5(n374), 
        .Y(n370) );
  OA221X1_LVT U302 ( .A1(n402), .A2(n397), .A3(n401), .A4(n400), .A5(n403), 
        .Y(n383) );
  OA221X1_LVT U303 ( .A1(n408), .A2(n388), .A3(n407), .A4(n406), .A5(n409), 
        .Y(n367) );
  NAND2X0_LVT U304 ( .A1(n333), .A2(n334), .Y(n363) );
  AND2X1_LVT U305 ( .A1(n419), .A2(n418), .Y(n333) );
  INVX1_LVT U306 ( .A(B[37]), .Y(n335) );
  NAND2X0_LVT U307 ( .A1(n335), .A2(A[37]), .Y(n334) );
  INVX1_LVT U308 ( .A(B[38]), .Y(n337) );
  INVX1_LVT U309 ( .A(n417), .Y(n338) );
  INVX1_LVT U310 ( .A(n378), .Y(n340) );
  AO222X1_LVT U311 ( .A1(n363), .A2(n364), .A3(n337), .A4(A[38]), .A5(n365), 
        .A6(n366), .Y(GE_LT_GT_LE) );
  OAI221X1_LVT U312 ( .A1(n367), .A2(n368), .A3(n369), .A4(n368), .A5(n370), 
        .Y(n366) );
  OA22X1_LVT U313 ( .A1(n348), .A2(B[30]), .A3(n375), .A4(B[29]), .Y(n374) );
  AO22X1_LVT U314 ( .A1(n376), .A2(n377), .A3(n376), .A4(n378), .Y(n373) );
  OA22X1_LVT U315 ( .A1(n349), .A2(B[28]), .A3(n381), .A4(B[27]), .Y(n372) );
  NAND2X0_LVT U316 ( .A1(A[27]), .A2(n382), .Y(n381) );
  AO221X1_LVT U317 ( .A1(n383), .A2(n384), .A3(n383), .A4(n385), .A5(n386), 
        .Y(n369) );
  OR3X1_LVT U318 ( .A1(n387), .A2(n388), .A3(n389), .Y(n386) );
  OA221X1_LVT U319 ( .A1(n391), .A2(n392), .A3(n393), .A4(n392), .A5(n394), 
        .Y(n385) );
  NAND2X0_LVT U320 ( .A1(B[4]), .A2(n362), .Y(n395) );
  OR3X1_LVT U321 ( .A1(n396), .A2(n397), .A3(n398), .Y(n384) );
  NAND2X0_LVT U322 ( .A1(B[8]), .A2(n360), .Y(n399) );
  NAND2X0_LVT U323 ( .A1(B[12]), .A2(n358), .Y(n404) );
  NAND4X0_LVT U324 ( .A1(n380), .A2(n340), .A3(n405), .A4(n379), .Y(n368) );
  NAND2X0_LVT U325 ( .A1(B[24]), .A2(n351), .Y(n379) );
  NAND2X0_LVT U326 ( .A1(B[23]), .A2(n352), .Y(n405) );
  NAND2X0_LVT U327 ( .A1(B[28]), .A2(n349), .Y(n382) );
  OA22X1_LVT U328 ( .A1(n353), .A2(B[22]), .A3(n410), .A4(B[21]), .Y(n409) );
  AO22X1_LVT U329 ( .A1(n411), .A2(n412), .A3(n411), .A4(n387), .Y(n408) );
  NAND2X0_LVT U330 ( .A1(B[16]), .A2(n356), .Y(n390) );
  OA22X1_LVT U331 ( .A1(n354), .A2(B[20]), .A3(n414), .A4(B[19]), .Y(n407) );
  NAND2X0_LVT U332 ( .A1(A[19]), .A2(n413), .Y(n414) );
  NAND2X0_LVT U333 ( .A1(B[20]), .A2(n354), .Y(n413) );
  AND4X1_LVT U334 ( .A1(n338), .A2(n339), .A3(n364), .A4(n415), .Y(n365) );
  AOI22X1_LVT U335 ( .A1(B[32]), .A2(n346), .A3(B[31]), .A4(n347), .Y(n415) );
  OA22X1_LVT U336 ( .A1(A[37]), .A2(n335), .A3(A[38]), .A4(n337), .Y(n364) );
  AO222X1_LVT U337 ( .A1(B[36]), .A2(n420), .A3(n343), .A4(n420), .A5(B[36]), 
        .A6(n343), .Y(n419) );
  OR2X1_LVT U338 ( .A1(n344), .A2(B[35]), .Y(n420) );
  AO221X1_LVT U339 ( .A1(n421), .A2(n416), .A3(n421), .A4(n422), .A5(n417), 
        .Y(n418) );
  AO22X1_LVT U340 ( .A1(n343), .A2(B[36]), .A3(n344), .A4(B[35]), .Y(n417) );
endmodule


module BreakpointUnit_DW_cmp_J40_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [38:0] A;
  input [38:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n299, n300, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423;

  AO221X1_LVT U201 ( .A1(1'b1), .A2(n390), .A3(B[11]), .A4(n302), .A5(n303), 
        .Y(n387) );
  AO221X1_LVT U202 ( .A1(1'b1), .A2(n399), .A3(B[19]), .A4(n299), .A5(n300), 
        .Y(n375) );
  NAND2X0_LVT U203 ( .A1(n340), .A2(B[10]), .Y(n284) );
  NAND2X0_LVT U204 ( .A1(A[9]), .A2(n284), .Y(n285) );
  NAND2X0_LVT U205 ( .A1(n389), .A2(A[7]), .Y(n286) );
  OA22X1_LVT U206 ( .A1(B[8]), .A2(n342), .A3(B[7]), .A4(n286), .Y(n287) );
  OA222X1_LVT U207 ( .A1(n285), .A2(B[9]), .A3(n340), .A4(B[10]), .A5(n386), 
        .A6(n287), .Y(n392) );
  INVX0_LVT U208 ( .A(A[0]), .Y(n288) );
  INVX0_LVT U209 ( .A(A[1]), .Y(n289) );
  INVX0_LVT U210 ( .A(A[2]), .Y(n290) );
  AO222X1_LVT U211 ( .A1(n288), .A2(B[0]), .A3(n289), .A4(B[1]), .A5(n290), 
        .A6(B[2]), .Y(n291) );
  NAND2X0_LVT U212 ( .A1(B[2]), .A2(n290), .Y(n292) );
  NAND2X0_LVT U213 ( .A1(A[1]), .A2(n292), .Y(n293) );
  OA22X1_LVT U214 ( .A1(B[1]), .A2(n293), .A3(B[2]), .A4(n290), .Y(n294) );
  INVX0_LVT U215 ( .A(A[3]), .Y(n295) );
  NAND2X0_LVT U216 ( .A1(B[3]), .A2(n295), .Y(n296) );
  NAND2X0_LVT U217 ( .A1(n294), .A2(n291), .Y(n297) );
  NAND3X0_LVT U218 ( .A1(n297), .A2(n385), .A3(n296), .Y(n378) );
  INVX0_LVT U220 ( .A(A[19]), .Y(n299) );
  INVX0_LVT U221 ( .A(n410), .Y(n300) );
  INVX0_LVT U223 ( .A(A[11]), .Y(n302) );
  INVX0_LVT U224 ( .A(n396), .Y(n303) );
  INVX1_LVT U225 ( .A(B[38]), .Y(n311) );
  INVX1_LVT U226 ( .A(B[37]), .Y(n309) );
  INVX1_LVT U227 ( .A(B[15]), .Y(n316) );
  INVX1_LVT U228 ( .A(B[7]), .Y(n317) );
  INVX1_LVT U229 ( .A(A[13]), .Y(n338) );
  INVX1_LVT U230 ( .A(A[12]), .Y(n339) );
  INVX1_LVT U231 ( .A(A[14]), .Y(n337) );
  INVX1_LVT U232 ( .A(A[10]), .Y(n340) );
  INVX1_LVT U233 ( .A(A[9]), .Y(n341) );
  INVX1_LVT U234 ( .A(A[8]), .Y(n342) );
  INVX1_LVT U235 ( .A(A[6]), .Y(n343) );
  INVX1_LVT U236 ( .A(A[5]), .Y(n344) );
  INVX1_LVT U237 ( .A(A[4]), .Y(n345) );
  INVX1_LVT U238 ( .A(A[31]), .Y(n323) );
  INVX1_LVT U239 ( .A(A[32]), .Y(n322) );
  INVX1_LVT U240 ( .A(A[34]), .Y(n320) );
  INVX1_LVT U241 ( .A(A[33]), .Y(n321) );
  INVX1_LVT U242 ( .A(A[35]), .Y(n319) );
  INVX1_LVT U243 ( .A(A[36]), .Y(n318) );
  INVX1_LVT U244 ( .A(A[17]), .Y(n335) );
  INVX1_LVT U245 ( .A(A[25]), .Y(n328) );
  INVX1_LVT U246 ( .A(A[24]), .Y(n329) );
  INVX1_LVT U247 ( .A(A[23]), .Y(n330) );
  INVX1_LVT U248 ( .A(A[16]), .Y(n336) );
  INVX1_LVT U249 ( .A(A[20]), .Y(n333) );
  INVX1_LVT U250 ( .A(A[22]), .Y(n331) );
  INVX1_LVT U251 ( .A(A[21]), .Y(n332) );
  INVX1_LVT U252 ( .A(A[18]), .Y(n334) );
  INVX1_LVT U253 ( .A(A[30]), .Y(n324) );
  INVX1_LVT U254 ( .A(A[29]), .Y(n325) );
  INVX1_LVT U255 ( .A(A[28]), .Y(n326) );
  INVX1_LVT U256 ( .A(A[27]), .Y(n306) );
  INVX1_LVT U257 ( .A(A[26]), .Y(n327) );
  INVX0_LVT U258 ( .A(n367), .Y(n310) );
  INVX0_LVT U259 ( .A(n354), .Y(n314) );
  OA221X1_LVT U260 ( .A1(n356), .A2(n310), .A3(n355), .A4(n354), .A5(n357), 
        .Y(n353) );
  OA221X1_LVT U261 ( .A1(n392), .A2(n387), .A3(n391), .A4(n390), .A5(n393), 
        .Y(n370) );
  AND2X1_LVT U262 ( .A1(n304), .A2(n305), .Y(n367) );
  AND2X1_LVT U263 ( .A1(n369), .A2(n314), .Y(n304) );
  NAND2X0_LVT U264 ( .A1(n306), .A2(B[27]), .Y(n305) );
  OA221X1_LVT U265 ( .A1(n401), .A2(n375), .A3(n400), .A4(n399), .A5(n402), 
        .Y(n350) );
  NAND2X0_LVT U266 ( .A1(n307), .A2(n308), .Y(n346) );
  AND2X1_LVT U267 ( .A1(n416), .A2(n415), .Y(n307) );
  NAND2X0_LVT U268 ( .A1(n309), .A2(A[37]), .Y(n308) );
  INVX1_LVT U269 ( .A(n414), .Y(n312) );
  INVX1_LVT U270 ( .A(n413), .Y(n313) );
  INVX1_LVT U271 ( .A(n362), .Y(n315) );
  AO222X1_LVT U272 ( .A1(n346), .A2(n347), .A3(n311), .A4(A[38]), .A5(n348), 
        .A6(n349), .Y(GE_LT_GT_LE) );
  OAI221X1_LVT U273 ( .A1(n350), .A2(n351), .A3(n352), .A4(n351), .A5(n353), 
        .Y(n349) );
  OA22X1_LVT U274 ( .A1(n324), .A2(B[30]), .A3(n358), .A4(B[29]), .Y(n357) );
  NAND2X0_LVT U275 ( .A1(A[29]), .A2(n359), .Y(n358) );
  NAND2X0_LVT U276 ( .A1(B[30]), .A2(n324), .Y(n359) );
  AO22X1_LVT U277 ( .A1(n360), .A2(n361), .A3(n360), .A4(n362), .Y(n356) );
  OA22X1_LVT U278 ( .A1(n329), .A2(B[24]), .A3(n363), .A4(B[23]), .Y(n361) );
  NAND2X0_LVT U279 ( .A1(A[23]), .A2(n364), .Y(n363) );
  OA22X1_LVT U280 ( .A1(B[26]), .A2(n327), .A3(B[25]), .A4(n365), .Y(n360) );
  NAND2X0_LVT U281 ( .A1(A[25]), .A2(n366), .Y(n365) );
  NAND2X0_LVT U282 ( .A1(B[26]), .A2(n327), .Y(n366) );
  OA22X1_LVT U283 ( .A1(n326), .A2(B[28]), .A3(n368), .A4(B[27]), .Y(n355) );
  NAND2X0_LVT U284 ( .A1(A[27]), .A2(n369), .Y(n368) );
  AO221X1_LVT U285 ( .A1(n370), .A2(n371), .A3(n370), .A4(n372), .A5(n373), 
        .Y(n352) );
  OR3X1_LVT U286 ( .A1(n374), .A2(n375), .A3(n376), .Y(n373) );
  OAI21X1_LVT U287 ( .A1(A[15]), .A2(n316), .A3(n377), .Y(n376) );
  OA221X1_LVT U288 ( .A1(n378), .A2(n379), .A3(n380), .A4(n379), .A5(n381), 
        .Y(n372) );
  OA22X1_LVT U289 ( .A1(n343), .A2(B[6]), .A3(n382), .A4(B[5]), .Y(n381) );
  NAND2X0_LVT U290 ( .A1(A[5]), .A2(n383), .Y(n382) );
  NAND2X0_LVT U291 ( .A1(B[6]), .A2(n343), .Y(n383) );
  OA22X1_LVT U292 ( .A1(n384), .A2(B[3]), .A3(n345), .A4(B[4]), .Y(n380) );
  NAND2X0_LVT U293 ( .A1(A[3]), .A2(n385), .Y(n384) );
  AO22X1_LVT U294 ( .A1(B[5]), .A2(n344), .A3(B[6]), .A4(n343), .Y(n379) );
  NAND2X0_LVT U295 ( .A1(B[4]), .A2(n345), .Y(n385) );
  OR3X1_LVT U296 ( .A1(n386), .A2(n387), .A3(n388), .Y(n371) );
  OAI21X1_LVT U297 ( .A1(A[7]), .A2(n317), .A3(n389), .Y(n388) );
  OA22X1_LVT U298 ( .A1(n337), .A2(B[14]), .A3(n394), .A4(B[13]), .Y(n393) );
  NAND2X0_LVT U299 ( .A1(A[13]), .A2(n395), .Y(n394) );
  NAND2X0_LVT U300 ( .A1(B[14]), .A2(n337), .Y(n395) );
  AO22X1_LVT U301 ( .A1(B[9]), .A2(n341), .A3(B[10]), .A4(n340), .Y(n386) );
  NAND2X0_LVT U302 ( .A1(B[8]), .A2(n342), .Y(n389) );
  OA22X1_LVT U303 ( .A1(n339), .A2(B[12]), .A3(n397), .A4(B[11]), .Y(n391) );
  NAND2X0_LVT U304 ( .A1(A[11]), .A2(n396), .Y(n397) );
  NAND2X0_LVT U305 ( .A1(B[12]), .A2(n339), .Y(n396) );
  AO22X1_LVT U306 ( .A1(B[13]), .A2(n338), .A3(B[14]), .A4(n337), .Y(n390) );
  NAND4X0_LVT U307 ( .A1(n367), .A2(n315), .A3(n398), .A4(n364), .Y(n351) );
  NAND2X0_LVT U308 ( .A1(B[24]), .A2(n329), .Y(n364) );
  NAND2X0_LVT U309 ( .A1(B[23]), .A2(n330), .Y(n398) );
  AO22X1_LVT U310 ( .A1(n328), .A2(B[25]), .A3(n327), .A4(B[26]), .Y(n362) );
  NAND2X0_LVT U311 ( .A1(B[28]), .A2(n326), .Y(n369) );
  AO22X1_LVT U312 ( .A1(n325), .A2(B[29]), .A3(n324), .A4(B[30]), .Y(n354) );
  OA22X1_LVT U313 ( .A1(n331), .A2(B[22]), .A3(n403), .A4(B[21]), .Y(n402) );
  NAND2X0_LVT U314 ( .A1(A[21]), .A2(n404), .Y(n403) );
  NAND2X0_LVT U315 ( .A1(B[22]), .A2(n331), .Y(n404) );
  AO22X1_LVT U316 ( .A1(n405), .A2(n406), .A3(n405), .A4(n374), .Y(n401) );
  AO22X1_LVT U317 ( .A1(B[17]), .A2(n335), .A3(B[18]), .A4(n334), .Y(n374) );
  OA22X1_LVT U318 ( .A1(n336), .A2(B[16]), .A3(n407), .A4(B[15]), .Y(n406) );
  NAND2X0_LVT U319 ( .A1(A[15]), .A2(n377), .Y(n407) );
  NAND2X0_LVT U320 ( .A1(B[16]), .A2(n336), .Y(n377) );
  OA22X1_LVT U321 ( .A1(B[18]), .A2(n334), .A3(B[17]), .A4(n408), .Y(n405) );
  NAND2X0_LVT U322 ( .A1(A[17]), .A2(n409), .Y(n408) );
  NAND2X0_LVT U323 ( .A1(B[18]), .A2(n334), .Y(n409) );
  OA22X1_LVT U324 ( .A1(n333), .A2(B[20]), .A3(n411), .A4(B[19]), .Y(n400) );
  NAND2X0_LVT U325 ( .A1(A[19]), .A2(n410), .Y(n411) );
  NAND2X0_LVT U326 ( .A1(B[20]), .A2(n333), .Y(n410) );
  AO22X1_LVT U327 ( .A1(B[21]), .A2(n332), .A3(B[22]), .A4(n331), .Y(n399) );
  AND4X1_LVT U328 ( .A1(n312), .A2(n313), .A3(n347), .A4(n412), .Y(n348) );
  AOI22X1_LVT U329 ( .A1(B[32]), .A2(n322), .A3(B[31]), .A4(n323), .Y(n412) );
  OA22X1_LVT U330 ( .A1(A[37]), .A2(n309), .A3(A[38]), .A4(n311), .Y(n347) );
  AO222X1_LVT U331 ( .A1(B[36]), .A2(n417), .A3(n318), .A4(n417), .A5(B[36]), 
        .A6(n318), .Y(n416) );
  OR2X1_LVT U332 ( .A1(n319), .A2(B[35]), .Y(n417) );
  AO221X1_LVT U333 ( .A1(n418), .A2(n413), .A3(n418), .A4(n419), .A5(n414), 
        .Y(n415) );
  AO22X1_LVT U334 ( .A1(n318), .A2(B[36]), .A3(n319), .A4(B[35]), .Y(n414) );
  OA22X1_LVT U335 ( .A1(n420), .A2(B[31]), .A3(n322), .A4(B[32]), .Y(n419) );
  NAND2X0_LVT U336 ( .A1(A[31]), .A2(n421), .Y(n420) );
  NAND2X0_LVT U337 ( .A1(B[32]), .A2(n322), .Y(n421) );
  AO22X1_LVT U338 ( .A1(n321), .A2(B[33]), .A3(n320), .A4(B[34]), .Y(n413) );
  OA22X1_LVT U339 ( .A1(B[34]), .A2(n320), .A3(B[33]), .A4(n422), .Y(n418) );
  NAND2X0_LVT U340 ( .A1(A[33]), .A2(n423), .Y(n422) );
  NAND2X0_LVT U341 ( .A1(B[34]), .A2(n320), .Y(n423) );
endmodule


module BreakpointUnit ( io_status_prv, io_bp_0_control_action, 
        io_bp_0_control_tmatch, io_bp_0_control_m, io_bp_0_control_s, 
        io_bp_0_control_u, io_bp_0_control_x, io_bp_0_control_w, 
        io_bp_0_control_r, io_bp_0_address, io_pc, io_ea, io_xcpt_if, 
        io_xcpt_ld, io_xcpt_st, io_debug_if, io_debug_ld, io_debug_st, 
        io_status_debug_BAR );
  input [1:0] io_status_prv;
  input [1:0] io_bp_0_control_tmatch;
  input [38:0] io_bp_0_address;
  input [38:0] io_pc;
  input [38:0] io_ea;
  input io_bp_0_control_action, io_bp_0_control_m, io_bp_0_control_s,
         io_bp_0_control_u, io_bp_0_control_x, io_bp_0_control_w,
         io_bp_0_control_r, io_status_debug_BAR;
  output io_xcpt_if, io_xcpt_ld, io_xcpt_st, io_debug_if, io_debug_ld,
         io_debug_st;
  wire   n_T_9, n_T_73, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n159, n160, n161, n162, n163, n164, n165, n166;

  BreakpointUnit_DW_cmp_J40_0 gte_x_5 ( .A(io_pc), .B(io_bp_0_address), .TC(
        1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b1), .GE_LT_GT_LE(n_T_73) );
  BreakpointUnit_DW_cmp_J40_1 gte_x_2 ( .A(io_ea), .B(io_bp_0_address), .TC(
        1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b1), .GE_LT_GT_LE(n_T_9) );
  INVX0_LVT U2 ( .A(io_status_prv[1]), .Y(n1) );
  AND2X1_LVT U3 ( .A1(io_bp_0_control_u), .A2(n1), .Y(n2) );
  INVX0_LVT U4 ( .A(io_status_prv[0]), .Y(n3) );
  AO22X1_LVT U5 ( .A1(io_status_prv[1]), .A2(io_bp_0_control_m), .A3(n1), .A4(
        io_bp_0_control_s), .Y(n4) );
  OA221X1_LVT U6 ( .A1(io_status_prv[0]), .A2(n2), .A3(n3), .A4(n4), .A5(
        io_status_debug_BAR), .Y(n67) );
  INVX0_LVT U7 ( .A(io_bp_0_address[28]), .Y(n125) );
  INVX1_LVT U8 ( .A(io_bp_0_address[29]), .Y(n126) );
  INVX1_LVT U9 ( .A(io_bp_0_address[1]), .Y(n133) );
  INVX1_LVT U10 ( .A(io_bp_0_address[2]), .Y(n135) );
  INVX1_LVT U11 ( .A(io_bp_0_address[27]), .Y(n122) );
  INVX1_LVT U12 ( .A(io_bp_0_address[37]), .Y(n123) );
  INVX1_LVT U13 ( .A(io_bp_0_address[4]), .Y(n119) );
  INVX1_LVT U14 ( .A(io_bp_0_address[5]), .Y(n120) );
  INVX1_LVT U15 ( .A(io_bp_0_address[12]), .Y(n117) );
  INVX1_LVT U16 ( .A(io_bp_0_address[6]), .Y(n148) );
  INVX1_LVT U17 ( .A(io_bp_0_address[8]), .Y(n145) );
  INVX1_LVT U18 ( .A(io_bp_0_address[14]), .Y(n144) );
  INVX1_LVT U19 ( .A(io_bp_0_address[17]), .Y(n141) );
  INVX1_LVT U20 ( .A(io_bp_0_address[11]), .Y(n142) );
  INVX1_LVT U21 ( .A(io_bp_0_address[22]), .Y(n76) );
  INVX1_LVT U22 ( .A(io_bp_0_address[26]), .Y(n72) );
  INVX1_LVT U23 ( .A(io_bp_0_address[33]), .Y(n73) );
  INVX1_LVT U24 ( .A(io_bp_0_address[3]), .Y(n79) );
  INVX1_LVT U25 ( .A(io_bp_0_address[24]), .Y(n139) );
  INVX1_LVT U26 ( .A(io_bp_0_address[21]), .Y(n138) );
  INVX1_LVT U27 ( .A(io_bp_0_address[16]), .Y(n110) );
  INVX0_LVT U28 ( .A(io_bp_0_address[20]), .Y(n109) );
  INVX1_LVT U29 ( .A(io_bp_0_address[38]), .Y(n106) );
  INVX1_LVT U30 ( .A(io_bp_0_address[19]), .Y(n107) );
  INVX1_LVT U31 ( .A(io_bp_0_address[32]), .Y(n103) );
  INVX1_LVT U32 ( .A(io_bp_0_address[34]), .Y(n104) );
  INVX1_LVT U33 ( .A(io_bp_0_address[30]), .Y(n100) );
  INVX1_LVT U34 ( .A(io_bp_0_address[31]), .Y(n101) );
  INVX1_LVT U35 ( .A(io_bp_0_address[10]), .Y(n90) );
  INVX1_LVT U36 ( .A(io_bp_0_address[25]), .Y(n91) );
  INVX1_LVT U37 ( .A(io_bp_0_address[35]), .Y(n88) );
  INVX1_LVT U38 ( .A(io_bp_0_address[36]), .Y(n87) );
  INVX1_LVT U39 ( .A(io_bp_0_address[23]), .Y(n84) );
  INVX1_LVT U40 ( .A(io_bp_0_control_tmatch[0]), .Y(n70) );
  INVX1_LVT U41 ( .A(io_bp_0_control_tmatch[1]), .Y(n163) );
  INVX1_LVT U42 ( .A(io_ea[1]), .Y(n132) );
  INVX1_LVT U43 ( .A(io_ea[22]), .Y(n77) );
  INVX1_LVT U44 ( .A(io_ea[0]), .Y(n74) );
  INVX1_LVT U45 ( .A(io_ea[3]), .Y(n78) );
  INVX1_LVT U46 ( .A(io_ea[2]), .Y(n136) );
  XOR2X1_LVT U47 ( .A1(n_T_73), .A2(io_bp_0_control_tmatch[0]), .Y(n63) );
  INVX0_LVT U48 ( .A(n_T_9), .Y(n161) );
  INVX0_LVT U49 ( .A(n68), .Y(n154) );
  XOR2X1_LVT U50 ( .A1(io_pc[20]), .A2(n109), .Y(n17) );
  XOR2X1_LVT U51 ( .A1(io_pc[28]), .A2(n125), .Y(n12) );
  XOR2X1_LVT U52 ( .A1(io_pc[9]), .A2(n85), .Y(n13) );
  XOR2X1_LVT U53 ( .A1(io_pc[15]), .A2(n116), .Y(n14) );
  XOR2X1_LVT U54 ( .A1(io_pc[13]), .A2(n93), .Y(n15) );
  XOR2X1_LVT U55 ( .A1(io_pc[23]), .A2(n84), .Y(n8) );
  XOR2X1_LVT U56 ( .A1(io_pc[18]), .A2(n94), .Y(n9) );
  XOR2X1_LVT U57 ( .A1(io_pc[35]), .A2(n88), .Y(n10) );
  XOR2X1_LVT U58 ( .A1(io_pc[1]), .A2(io_bp_0_address[1]), .Y(n23) );
  XOR2X1_LVT U59 ( .A1(io_pc[0]), .A2(n131), .Y(n49) );
  XOR2X1_LVT U60 ( .A1(io_pc[3]), .A2(n79), .Y(n44) );
  XOR2X1_LVT U61 ( .A1(io_pc[7]), .A2(n147), .Y(n30) );
  XOR2X1_LVT U62 ( .A1(io_pc[31]), .A2(n101), .Y(n27) );
  XOR2X1_LVT U63 ( .A1(io_pc[27]), .A2(n122), .Y(n18) );
  XOR2X1_LVT U64 ( .A1(io_pc[29]), .A2(n126), .Y(n20) );
  XOR2X1_LVT U65 ( .A1(io_pc[38]), .A2(n106), .Y(n11) );
  NOR4X1_LVT U66 ( .A1(n160), .A2(n159), .A3(n156), .A4(n155), .Y(n164) );
  XOR2X1_LVT U67 ( .A1(io_pc[34]), .A2(n104), .Y(n51) );
  XOR2X1_LVT U68 ( .A1(io_pc[33]), .A2(n73), .Y(n52) );
  XOR2X1_LVT U69 ( .A1(io_pc[5]), .A2(n120), .Y(n53) );
  XOR2X1_LVT U70 ( .A1(io_pc[37]), .A2(n123), .Y(n54) );
  XOR2X1_LVT U71 ( .A1(io_pc[2]), .A2(n135), .Y(n50) );
  XOR2X1_LVT U72 ( .A1(io_pc[4]), .A2(n119), .Y(n45) );
  XOR2X1_LVT U73 ( .A1(io_pc[14]), .A2(n144), .Y(n46) );
  XOR2X1_LVT U74 ( .A1(io_pc[12]), .A2(n117), .Y(n47) );
  XOR2X1_LVT U75 ( .A1(io_pc[36]), .A2(n87), .Y(n36) );
  XOR2X1_LVT U76 ( .A1(io_pc[10]), .A2(n90), .Y(n37) );
  XOR2X1_LVT U77 ( .A1(io_pc[6]), .A2(n148), .Y(n38) );
  XOR2X1_LVT U78 ( .A1(io_pc[11]), .A2(n142), .Y(n39) );
  XOR2X1_LVT U79 ( .A1(io_pc[21]), .A2(n138), .Y(n32) );
  XOR2X1_LVT U80 ( .A1(io_pc[17]), .A2(n141), .Y(n33) );
  XOR2X1_LVT U81 ( .A1(io_pc[24]), .A2(n139), .Y(n34) );
  XOR2X1_LVT U82 ( .A1(io_pc[22]), .A2(n76), .Y(n35) );
  XOR2X1_LVT U83 ( .A1(io_pc[25]), .A2(n91), .Y(n28) );
  XOR2X1_LVT U84 ( .A1(io_pc[8]), .A2(n145), .Y(n29) );
  XOR2X1_LVT U85 ( .A1(io_pc[19]), .A2(n107), .Y(n31) );
  XOR2X1_LVT U86 ( .A1(io_pc[16]), .A2(n110), .Y(n24) );
  XOR2X1_LVT U87 ( .A1(io_pc[30]), .A2(n100), .Y(n25) );
  XOR2X1_LVT U88 ( .A1(io_pc[32]), .A2(n103), .Y(n26) );
  XOR2X1_LVT U89 ( .A1(io_pc[26]), .A2(n72), .Y(n19) );
  AND4X1_LVT U90 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .Y(n5) );
  AND4X1_LVT U91 ( .A1(n130), .A2(n129), .A3(n128), .A4(n127), .Y(n6) );
  NAND2X0_LVT U92 ( .A1(n154), .A2(n153), .Y(n7) );
  NAND3X0_LVT U93 ( .A1(n5), .A2(n6), .A3(n7), .Y(n155) );
  INVX1_LVT U94 ( .A(io_bp_0_address[0]), .Y(n131) );
  AND2X1_LVT U95 ( .A1(io_bp_0_address[0]), .A2(io_bp_0_control_tmatch[0]), 
        .Y(n16) );
  AND2X1_LVT U96 ( .A1(n16), .A2(io_bp_0_address[1]), .Y(n68) );
  INVX1_LVT U97 ( .A(io_bp_0_address[9]), .Y(n85) );
  INVX1_LVT U98 ( .A(io_bp_0_address[18]), .Y(n94) );
  INVX1_LVT U99 ( .A(io_bp_0_address[13]), .Y(n93) );
  INVX1_LVT U100 ( .A(io_bp_0_address[15]), .Y(n116) );
  INVX1_LVT U101 ( .A(io_bp_0_address[7]), .Y(n147) );
  INVX1_LVT U102 ( .A(io_bp_0_control_action), .Y(n69) );
  NAND4X0_LVT U103 ( .A1(n11), .A2(n10), .A3(n9), .A4(n8), .Y(n62) );
  NAND4X0_LVT U104 ( .A1(n15), .A2(n14), .A3(n13), .A4(n12), .Y(n61) );
  INVX1_LVT U105 ( .A(n16), .Y(n22) );
  NAND4X0_LVT U106 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .Y(n21) );
  AO21X1_LVT U107 ( .A1(n23), .A2(n22), .A3(n21), .Y(n60) );
  NAND4X0_LVT U108 ( .A1(n27), .A2(n26), .A3(n25), .A4(n24), .Y(n43) );
  NAND4X0_LVT U109 ( .A1(n31), .A2(n30), .A3(n29), .A4(n28), .Y(n42) );
  NAND4X0_LVT U110 ( .A1(n35), .A2(n34), .A3(n33), .A4(n32), .Y(n41) );
  NAND4X0_LVT U111 ( .A1(n39), .A2(n38), .A3(n37), .A4(n36), .Y(n40) );
  NOR4X1_LVT U112 ( .A1(n43), .A2(n42), .A3(n41), .A4(n40), .Y(n58) );
  AO21X1_LVT U113 ( .A1(io_bp_0_address[2]), .A2(n68), .A3(n44), .Y(n48) );
  AND4X1_LVT U114 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .Y(n57) );
  OA22X1_LVT U115 ( .A1(n68), .A2(n50), .A3(io_bp_0_control_tmatch[0]), .A4(
        n49), .Y(n56) );
  AND4X1_LVT U116 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .Y(n55) );
  NAND4X0_LVT U117 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .Y(n59) );
  NOR4X1_LVT U118 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .Y(n64) );
  MUX21X1_LVT U119 ( .A1(n64), .A2(n63), .S0(io_bp_0_control_tmatch[1]), .Y(
        n65) );
  AND3X1_LVT U120 ( .A1(n65), .A2(n67), .A3(io_bp_0_control_x), .Y(n66) );
  AND2X1_LVT U121 ( .A1(n66), .A2(io_bp_0_control_action), .Y(io_debug_if) );
  AND2X1_LVT U122 ( .A1(n66), .A2(n69), .Y(io_xcpt_if) );
  AOI22X1_LVT U125 ( .A1(n73), .A2(io_ea[33]), .A3(n72), .A4(io_ea[26]), .Y(
        n71) );
  OA221X1_LVT U126 ( .A1(n73), .A2(io_ea[33]), .A3(n72), .A4(io_ea[26]), .A5(
        n71), .Y(n82) );
  AO22X1_LVT U127 ( .A1(io_bp_0_address[0]), .A2(io_ea[0]), .A3(n131), .A4(n74), .Y(n75) );
  OA222X1_LVT U128 ( .A1(io_bp_0_address[22]), .A2(n77), .A3(n76), .A4(
        io_ea[22]), .A5(io_bp_0_control_tmatch[0]), .A6(n75), .Y(n81) );
  AO222X1_LVT U129 ( .A1(io_bp_0_address[3]), .A2(io_ea[3]), .A3(n79), .A4(n78), .A5(n68), .A6(io_bp_0_address[2]), .Y(n80) );
  NAND3X0_LVT U130 ( .A1(n82), .A2(n81), .A3(n80), .Y(n160) );
  AOI22X1_LVT U131 ( .A1(n84), .A2(io_ea[23]), .A3(n85), .A4(io_ea[9]), .Y(n83) );
  OA221X1_LVT U132 ( .A1(n85), .A2(io_ea[9]), .A3(n84), .A4(io_ea[23]), .A5(
        n83), .Y(n98) );
  AOI22X1_LVT U133 ( .A1(n87), .A2(io_ea[36]), .A3(n88), .A4(io_ea[35]), .Y(
        n86) );
  OA221X1_LVT U134 ( .A1(n88), .A2(io_ea[35]), .A3(n87), .A4(io_ea[36]), .A5(
        n86), .Y(n97) );
  AOI22X1_LVT U135 ( .A1(n91), .A2(io_ea[25]), .A3(n90), .A4(io_ea[10]), .Y(
        n89) );
  OA221X1_LVT U136 ( .A1(n91), .A2(io_ea[25]), .A3(n90), .A4(io_ea[10]), .A5(
        n89), .Y(n96) );
  AOI22X1_LVT U137 ( .A1(n94), .A2(io_ea[18]), .A3(n93), .A4(io_ea[13]), .Y(
        n92) );
  OA221X1_LVT U138 ( .A1(n94), .A2(io_ea[18]), .A3(n93), .A4(io_ea[13]), .A5(
        n92), .Y(n95) );
  NAND4X0_LVT U139 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .Y(n159) );
  AOI22X1_LVT U140 ( .A1(n101), .A2(io_ea[31]), .A3(n100), .A4(io_ea[30]), .Y(
        n99) );
  OA221X1_LVT U141 ( .A1(n101), .A2(io_ea[31]), .A3(n100), .A4(io_ea[30]), 
        .A5(n99), .Y(n114) );
  AOI22X1_LVT U142 ( .A1(n104), .A2(io_ea[34]), .A3(n103), .A4(io_ea[32]), .Y(
        n102) );
  OA221X1_LVT U143 ( .A1(n104), .A2(io_ea[34]), .A3(n103), .A4(io_ea[32]), 
        .A5(n102), .Y(n113) );
  AOI22X1_LVT U144 ( .A1(n107), .A2(io_ea[19]), .A3(n106), .A4(io_ea[38]), .Y(
        n105) );
  OA221X1_LVT U145 ( .A1(n107), .A2(io_ea[19]), .A3(n106), .A4(io_ea[38]), 
        .A5(n105), .Y(n112) );
  AOI22X1_LVT U146 ( .A1(n109), .A2(io_ea[20]), .A3(n110), .A4(io_ea[16]), .Y(
        n108) );
  OA221X1_LVT U147 ( .A1(n110), .A2(io_ea[16]), .A3(n109), .A4(io_ea[20]), 
        .A5(n108), .Y(n111) );
  NAND4X0_LVT U148 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .Y(n156) );
  AOI22X1_LVT U149 ( .A1(n117), .A2(io_ea[12]), .A3(n116), .A4(io_ea[15]), .Y(
        n115) );
  OA221X1_LVT U150 ( .A1(n117), .A2(io_ea[12]), .A3(n116), .A4(io_ea[15]), 
        .A5(n115), .Y(n130) );
  AOI22X1_LVT U151 ( .A1(n120), .A2(io_ea[5]), .A3(n119), .A4(io_ea[4]), .Y(
        n118) );
  OA221X1_LVT U152 ( .A1(n120), .A2(io_ea[5]), .A3(n119), .A4(io_ea[4]), .A5(
        n118), .Y(n129) );
  AOI22X1_LVT U153 ( .A1(n122), .A2(io_ea[27]), .A3(n123), .A4(io_ea[37]), .Y(
        n121) );
  OA221X1_LVT U154 ( .A1(n123), .A2(io_ea[37]), .A3(n122), .A4(io_ea[27]), 
        .A5(n121), .Y(n128) );
  AOI22X1_LVT U155 ( .A1(n126), .A2(io_ea[29]), .A3(n125), .A4(io_ea[28]), .Y(
        n124) );
  OA221X1_LVT U156 ( .A1(n126), .A2(io_ea[29]), .A3(n125), .A4(io_ea[28]), 
        .A5(n124), .Y(n127) );
  OA222X1_LVT U157 ( .A1(io_bp_0_address[1]), .A2(io_ea[1]), .A3(n133), .A4(
        n132), .A5(n70), .A6(n131), .Y(n134) );
  AO221X1_LVT U158 ( .A1(io_bp_0_address[2]), .A2(n136), .A3(n135), .A4(
        io_ea[2]), .A5(n134), .Y(n153) );
  AOI22X1_LVT U159 ( .A1(n138), .A2(io_ea[21]), .A3(n139), .A4(io_ea[24]), .Y(
        n137) );
  OA221X1_LVT U160 ( .A1(n139), .A2(io_ea[24]), .A3(n138), .A4(io_ea[21]), 
        .A5(n137), .Y(n152) );
  AOI22X1_LVT U161 ( .A1(n142), .A2(io_ea[11]), .A3(n141), .A4(io_ea[17]), .Y(
        n140) );
  OA221X1_LVT U162 ( .A1(n142), .A2(io_ea[11]), .A3(n141), .A4(io_ea[17]), 
        .A5(n140), .Y(n151) );
  AOI22X1_LVT U163 ( .A1(n144), .A2(io_ea[14]), .A3(n145), .A4(io_ea[8]), .Y(
        n143) );
  OA221X1_LVT U164 ( .A1(n145), .A2(io_ea[8]), .A3(n144), .A4(io_ea[14]), .A5(
        n143), .Y(n150) );
  AOI22X1_LVT U165 ( .A1(n148), .A2(io_ea[6]), .A3(n147), .A4(io_ea[7]), .Y(
        n146) );
  OA221X1_LVT U166 ( .A1(n148), .A2(io_ea[6]), .A3(n147), .A4(io_ea[7]), .A5(
        n146), .Y(n149) );
  AO22X1_LVT U167 ( .A1(io_bp_0_control_tmatch[0]), .A2(n161), .A3(n70), .A4(
        n_T_9), .Y(n162) );
  OA221X1_LVT U168 ( .A1(io_bp_0_control_tmatch[1]), .A2(n164), .A3(n163), 
        .A4(n162), .A5(n67), .Y(n166) );
  AND2X1_LVT U169 ( .A1(n166), .A2(io_bp_0_control_r), .Y(n165) );
  AND2X1_LVT U170 ( .A1(io_bp_0_control_action), .A2(n165), .Y(io_debug_ld) );
  AND3X1_LVT U171 ( .A1(io_bp_0_control_action), .A2(n166), .A3(
        io_bp_0_control_w), .Y(io_debug_st) );
  AND2X1_LVT U172 ( .A1(n165), .A2(n69), .Y(io_xcpt_ld) );
  AND3X1_LVT U173 ( .A1(n166), .A2(io_bp_0_control_w), .A3(n69), .Y(io_xcpt_st) );
endmodule


module ALU_DP_OP_31J40_124_1870_J40_0 ( I1, I2, I3, O1 );
  input [63:0] I1;
  input [63:0] I2;
  output [63:0] O1;
  input I3;
  wire   n442, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917;

  FADDX1_LVT U568 ( .A(I1[0]), .B(I2[0]), .CI(I3), .CO(n442), .S(O1[0]) );
  AO222X1_LVT U571 ( .A1(I1[52]), .A2(I2[52]), .A3(I1[52]), .A4(n752), .A5(
        I2[52]), .A6(n752), .Y(n741) );
  OR2X1_LVT U572 ( .A1(I1[58]), .A2(I2[58]), .Y(n703) );
  AO222X1_LVT U573 ( .A1(n703), .A2(n731), .A3(n733), .A4(n732), .A5(I1[58]), 
        .A6(I2[58]), .Y(n720) );
  AO222X1_LVT U574 ( .A1(I1[40]), .A2(I2[40]), .A3(I1[40]), .A4(n789), .A5(
        I2[40]), .A6(n789), .Y(n785) );
  AO222X1_LVT U575 ( .A1(I1[44]), .A2(I2[44]), .A3(I1[44]), .A4(n779), .A5(
        I2[44]), .A6(n779), .Y(n772) );
  AO222X1_LVT U576 ( .A1(I1[60]), .A2(I2[60]), .A3(I1[60]), .A4(n728), .A5(
        I2[60]), .A6(n728), .Y(n718) );
  AO222X1_LVT U577 ( .A1(I1[56]), .A2(I2[56]), .A3(I1[56]), .A4(n737), .A5(
        I2[56]), .A6(n737), .Y(n733) );
  OA222X1_LVT U578 ( .A1(n873), .A2(n874), .A3(n873), .A4(n875), .A5(n873), 
        .A6(n876), .Y(n827) );
  OA222X1_LVT U579 ( .A1(n913), .A2(n442), .A3(n913), .A4(n914), .A5(n913), 
        .A6(n915), .Y(n906) );
  AND2X1_LVT U580 ( .A1(n721), .A2(n722), .Y(n713) );
  FADDX1_LVT U581 ( .A(n704), .B(I1[63]), .CI(I2[63]), .S(O1[63]) );
  OA222X1_LVT U582 ( .A1(n705), .A2(n706), .A3(n705), .A4(n707), .A5(n705), 
        .A6(n708), .Y(n704) );
  AO221X1_LVT U583 ( .A1(n709), .A2(n707), .A3(n710), .A4(n711), .A5(n712), 
        .Y(n705) );
  NAND3X0_LVT U584 ( .A1(n713), .A2(n714), .A3(n715), .Y(n712) );
  NAND3X0_LVT U585 ( .A1(n716), .A2(n717), .A3(n718), .Y(n715) );
  NAND4X0_LVT U586 ( .A1(n719), .A2(n720), .A3(n716), .A4(n717), .Y(n714) );
  NAND3X0_LVT U587 ( .A1(I1[61]), .A2(I2[61]), .A3(n717), .Y(n722) );
  NAND2X0_LVT U588 ( .A1(I1[62]), .A2(I2[62]), .Y(n721) );
  AND2X1_LVT U589 ( .A1(n723), .A2(n710), .Y(n707) );
  AND4X1_LVT U590 ( .A1(n719), .A2(n724), .A3(n716), .A4(n717), .Y(n710) );
  OR2X1_LVT U591 ( .A1(I1[62]), .A2(I2[62]), .Y(n717) );
  FADDX1_LVT U592 ( .A(I1[62]), .B(I2[62]), .CI(n725), .S(O1[62]) );
  AO22X1_LVT U593 ( .A1(I1[61]), .A2(I2[61]), .A3(n726), .A4(n716), .Y(n725)
         );
  OR2X1_LVT U594 ( .A1(I1[61]), .A2(I2[61]), .Y(n716) );
  FADDX1_LVT U595 ( .A(I1[61]), .B(I2[61]), .CI(n726), .S(O1[61]) );
  AO21X1_LVT U596 ( .A1(n719), .A2(n727), .A3(n718), .Y(n726) );
  OA22X1_LVT U597 ( .A1(I1[60]), .A2(I2[60]), .A3(I1[59]), .A4(I2[59]), .Y(
        n719) );
  FADDX1_LVT U598 ( .A(I1[60]), .B(I2[60]), .CI(n729), .S(O1[60]) );
  AO221X1_LVT U599 ( .A1(n727), .A2(I1[59]), .A3(n727), .A4(I2[59]), .A5(n728), 
        .Y(n729) );
  AND2X1_LVT U600 ( .A1(I1[59]), .A2(I2[59]), .Y(n728) );
  FADDX1_LVT U601 ( .A(I1[59]), .B(I2[59]), .CI(n727), .S(O1[59]) );
  AO21X1_LVT U602 ( .A1(n724), .A2(n730), .A3(n720), .Y(n727) );
  AND2X1_LVT U603 ( .A1(n732), .A2(n734), .Y(n724) );
  OA22X1_LVT U604 ( .A1(I1[58]), .A2(I2[58]), .A3(I1[57]), .A4(I2[57]), .Y(
        n732) );
  FADDX1_LVT U605 ( .A(I1[58]), .B(I2[58]), .CI(n735), .S(O1[58]) );
  OA22X1_LVT U606 ( .A1(n731), .A2(n736), .A3(I1[57]), .A4(I2[57]), .Y(n735)
         );
  AND2X1_LVT U607 ( .A1(I1[57]), .A2(I2[57]), .Y(n731) );
  FADDX1_LVT U608 ( .A(I1[57]), .B(I2[57]), .CI(n736), .S(O1[57]) );
  AO21X1_LVT U609 ( .A1(n734), .A2(n730), .A3(n733), .Y(n736) );
  OA22X1_LVT U610 ( .A1(I1[56]), .A2(I2[56]), .A3(I1[55]), .A4(I2[55]), .Y(
        n734) );
  FADDX1_LVT U611 ( .A(I1[56]), .B(I2[56]), .CI(n738), .S(O1[56]) );
  OA22X1_LVT U612 ( .A1(n737), .A2(n730), .A3(I1[55]), .A4(I2[55]), .Y(n738)
         );
  AND2X1_LVT U613 ( .A1(I1[55]), .A2(I2[55]), .Y(n737) );
  FADDX1_LVT U614 ( .A(I1[55]), .B(I2[55]), .CI(n730), .S(O1[55]) );
  AO21X1_LVT U615 ( .A1(n723), .A2(n739), .A3(n711), .Y(n730) );
  AO221X1_LVT U616 ( .A1(n740), .A2(n741), .A3(n742), .A4(n743), .A5(n744), 
        .Y(n711) );
  AO22X1_LVT U617 ( .A1(I1[54]), .A2(I2[54]), .A3(n745), .A4(n746), .Y(n744)
         );
  OR2X1_LVT U618 ( .A1(I2[54]), .A2(I1[54]), .Y(n746) );
  AND2X1_LVT U619 ( .A1(n743), .A2(n747), .Y(n723) );
  AND2X1_LVT U620 ( .A1(n740), .A2(n748), .Y(n743) );
  OA22X1_LVT U621 ( .A1(I1[54]), .A2(I2[54]), .A3(I1[53]), .A4(I2[53]), .Y(
        n740) );
  FADDX1_LVT U622 ( .A(I1[54]), .B(I2[54]), .CI(n749), .S(O1[54]) );
  OA22X1_LVT U623 ( .A1(n745), .A2(n750), .A3(I1[53]), .A4(I2[53]), .Y(n749)
         );
  AND2X1_LVT U624 ( .A1(I1[53]), .A2(I2[53]), .Y(n745) );
  FADDX1_LVT U625 ( .A(I1[53]), .B(I2[53]), .CI(n750), .S(O1[53]) );
  AO21X1_LVT U626 ( .A1(n748), .A2(n751), .A3(n741), .Y(n750) );
  OA22X1_LVT U627 ( .A1(I1[52]), .A2(I2[52]), .A3(I1[51]), .A4(I2[51]), .Y(
        n748) );
  FADDX1_LVT U628 ( .A(I1[52]), .B(I2[52]), .CI(n753), .S(O1[52]) );
  OA22X1_LVT U629 ( .A1(n752), .A2(n751), .A3(I1[51]), .A4(I2[51]), .Y(n753)
         );
  AND2X1_LVT U630 ( .A1(I1[51]), .A2(I2[51]), .Y(n752) );
  FADDX1_LVT U631 ( .A(I1[51]), .B(I2[51]), .CI(n751), .S(O1[51]) );
  AO21X1_LVT U632 ( .A1(n747), .A2(n739), .A3(n742), .Y(n751) );
  AO222X1_LVT U633 ( .A1(I1[50]), .A2(I2[50]), .A3(n754), .A4(n755), .A5(n756), 
        .A6(n757), .Y(n742) );
  OR2X1_LVT U634 ( .A1(I2[50]), .A2(I1[50]), .Y(n755) );
  AND2X1_LVT U635 ( .A1(n756), .A2(n758), .Y(n747) );
  OA22X1_LVT U636 ( .A1(I1[50]), .A2(I2[50]), .A3(I1[49]), .A4(I2[49]), .Y(
        n756) );
  FADDX1_LVT U637 ( .A(I1[50]), .B(I2[50]), .CI(n759), .S(O1[50]) );
  OA22X1_LVT U638 ( .A1(n754), .A2(n760), .A3(I1[49]), .A4(I2[49]), .Y(n759)
         );
  AND2X1_LVT U639 ( .A1(I1[49]), .A2(I2[49]), .Y(n754) );
  FADDX1_LVT U640 ( .A(I1[49]), .B(I2[49]), .CI(n760), .S(O1[49]) );
  AO21X1_LVT U641 ( .A1(n758), .A2(n739), .A3(n757), .Y(n760) );
  AO22X1_LVT U642 ( .A1(I1[48]), .A2(I2[48]), .A3(n761), .A4(n762), .Y(n757)
         );
  OR2X1_LVT U643 ( .A1(I1[48]), .A2(I2[48]), .Y(n762) );
  OA22X1_LVT U644 ( .A1(I1[48]), .A2(I2[48]), .A3(I1[47]), .A4(I2[47]), .Y(
        n758) );
  FADDX1_LVT U645 ( .A(I1[48]), .B(I2[48]), .CI(n763), .S(O1[48]) );
  OA22X1_LVT U646 ( .A1(n761), .A2(n739), .A3(I1[47]), .A4(I2[47]), .Y(n763)
         );
  AND2X1_LVT U647 ( .A1(I1[47]), .A2(I2[47]), .Y(n761) );
  FADDX1_LVT U648 ( .A(I1[47]), .B(I2[47]), .CI(n739), .S(O1[47]) );
  AO21X1_LVT U649 ( .A1(n706), .A2(n708), .A3(n709), .Y(n739) );
  AO221X1_LVT U650 ( .A1(n764), .A2(n765), .A3(n766), .A4(n767), .A5(n768), 
        .Y(n709) );
  AO222X1_LVT U651 ( .A1(I1[46]), .A2(I2[46]), .A3(n769), .A4(n770), .A5(n771), 
        .A6(n772), .Y(n768) );
  OR2X1_LVT U652 ( .A1(I2[46]), .A2(I1[46]), .Y(n770) );
  AND2X1_LVT U653 ( .A1(n766), .A2(n773), .Y(n706) );
  AND2X1_LVT U654 ( .A1(n774), .A2(n765), .Y(n766) );
  AND2X1_LVT U655 ( .A1(n771), .A2(n775), .Y(n765) );
  OA22X1_LVT U656 ( .A1(I1[46]), .A2(I2[46]), .A3(I1[45]), .A4(I2[45]), .Y(
        n771) );
  FADDX1_LVT U657 ( .A(I1[46]), .B(I2[46]), .CI(n776), .S(O1[46]) );
  OA22X1_LVT U658 ( .A1(n769), .A2(n777), .A3(I1[45]), .A4(I2[45]), .Y(n776)
         );
  AND2X1_LVT U659 ( .A1(I1[45]), .A2(I2[45]), .Y(n769) );
  FADDX1_LVT U660 ( .A(I1[45]), .B(I2[45]), .CI(n777), .S(O1[45]) );
  AO21X1_LVT U661 ( .A1(n775), .A2(n778), .A3(n772), .Y(n777) );
  OA22X1_LVT U662 ( .A1(I1[44]), .A2(I2[44]), .A3(I1[43]), .A4(I2[43]), .Y(
        n775) );
  FADDX1_LVT U663 ( .A(I1[44]), .B(I2[44]), .CI(n780), .S(O1[44]) );
  OA22X1_LVT U664 ( .A1(n779), .A2(n778), .A3(I1[43]), .A4(I2[43]), .Y(n780)
         );
  AND2X1_LVT U665 ( .A1(I1[43]), .A2(I2[43]), .Y(n779) );
  FADDX1_LVT U666 ( .A(I1[43]), .B(I2[43]), .CI(n778), .S(O1[43]) );
  AO21X1_LVT U667 ( .A1(n774), .A2(n781), .A3(n764), .Y(n778) );
  AO222X1_LVT U668 ( .A1(I1[42]), .A2(I2[42]), .A3(n782), .A4(n783), .A5(n784), 
        .A6(n785), .Y(n764) );
  OR2X1_LVT U669 ( .A1(I2[42]), .A2(I1[42]), .Y(n783) );
  AND2X1_LVT U670 ( .A1(n784), .A2(n786), .Y(n774) );
  OA22X1_LVT U671 ( .A1(I1[42]), .A2(I2[42]), .A3(I1[41]), .A4(I2[41]), .Y(
        n784) );
  FADDX1_LVT U672 ( .A(I1[42]), .B(I2[42]), .CI(n787), .S(O1[42]) );
  OA22X1_LVT U673 ( .A1(n782), .A2(n788), .A3(I1[41]), .A4(I2[41]), .Y(n787)
         );
  AND2X1_LVT U674 ( .A1(I1[41]), .A2(I2[41]), .Y(n782) );
  FADDX1_LVT U675 ( .A(I1[41]), .B(I2[41]), .CI(n788), .S(O1[41]) );
  AO21X1_LVT U676 ( .A1(n786), .A2(n781), .A3(n785), .Y(n788) );
  OA22X1_LVT U677 ( .A1(I1[40]), .A2(I2[40]), .A3(I1[39]), .A4(I2[39]), .Y(
        n786) );
  FADDX1_LVT U678 ( .A(I1[40]), .B(I2[40]), .CI(n790), .S(O1[40]) );
  OA22X1_LVT U679 ( .A1(n789), .A2(n781), .A3(I1[39]), .A4(I2[39]), .Y(n790)
         );
  AND2X1_LVT U680 ( .A1(I1[39]), .A2(I2[39]), .Y(n789) );
  FADDX1_LVT U681 ( .A(I1[39]), .B(I2[39]), .CI(n781), .S(O1[39]) );
  AO21X1_LVT U682 ( .A1(n773), .A2(n708), .A3(n767), .Y(n781) );
  AO221X1_LVT U683 ( .A1(n791), .A2(n792), .A3(n793), .A4(n794), .A5(n795), 
        .Y(n767) );
  AO22X1_LVT U684 ( .A1(I1[38]), .A2(I2[38]), .A3(n796), .A4(n797), .Y(n795)
         );
  OR2X1_LVT U685 ( .A1(I2[38]), .A2(I1[38]), .Y(n797) );
  AND2X1_LVT U686 ( .A1(n794), .A2(n798), .Y(n773) );
  AND2X1_LVT U687 ( .A1(n791), .A2(n799), .Y(n794) );
  OA22X1_LVT U688 ( .A1(I1[38]), .A2(I2[38]), .A3(I1[37]), .A4(I2[37]), .Y(
        n791) );
  FADDX1_LVT U689 ( .A(I1[38]), .B(I2[38]), .CI(n800), .S(O1[38]) );
  OA22X1_LVT U690 ( .A1(n796), .A2(n801), .A3(I1[37]), .A4(I2[37]), .Y(n800)
         );
  AND2X1_LVT U691 ( .A1(I1[37]), .A2(I2[37]), .Y(n796) );
  FADDX1_LVT U692 ( .A(I1[37]), .B(I2[37]), .CI(n801), .S(O1[37]) );
  AO21X1_LVT U693 ( .A1(n799), .A2(n802), .A3(n792), .Y(n801) );
  AO22X1_LVT U694 ( .A1(I1[36]), .A2(I2[36]), .A3(n803), .A4(n804), .Y(n792)
         );
  OR2X1_LVT U695 ( .A1(I1[36]), .A2(I2[36]), .Y(n804) );
  OA22X1_LVT U696 ( .A1(I1[36]), .A2(I2[36]), .A3(I1[35]), .A4(I2[35]), .Y(
        n799) );
  FADDX1_LVT U697 ( .A(I1[36]), .B(I2[36]), .CI(n805), .S(O1[36]) );
  OA22X1_LVT U698 ( .A1(n803), .A2(n802), .A3(I1[35]), .A4(I2[35]), .Y(n805)
         );
  AND2X1_LVT U699 ( .A1(I1[35]), .A2(I2[35]), .Y(n803) );
  FADDX1_LVT U700 ( .A(I1[35]), .B(I2[35]), .CI(n802), .S(O1[35]) );
  AO21X1_LVT U701 ( .A1(n798), .A2(n708), .A3(n793), .Y(n802) );
  AO222X1_LVT U702 ( .A1(I1[34]), .A2(I2[34]), .A3(n806), .A4(n807), .A5(n808), 
        .A6(n809), .Y(n793) );
  OR2X1_LVT U703 ( .A1(I2[34]), .A2(I1[34]), .Y(n807) );
  AND2X1_LVT U704 ( .A1(n808), .A2(n810), .Y(n798) );
  OA22X1_LVT U705 ( .A1(I1[34]), .A2(I2[34]), .A3(I1[33]), .A4(I2[33]), .Y(
        n808) );
  FADDX1_LVT U706 ( .A(I1[34]), .B(I2[34]), .CI(n811), .S(O1[34]) );
  OA22X1_LVT U707 ( .A1(n806), .A2(n812), .A3(I1[33]), .A4(I2[33]), .Y(n811)
         );
  AND2X1_LVT U708 ( .A1(I1[33]), .A2(I2[33]), .Y(n806) );
  FADDX1_LVT U709 ( .A(I1[33]), .B(I2[33]), .CI(n812), .S(O1[33]) );
  AO21X1_LVT U710 ( .A1(n810), .A2(n708), .A3(n809), .Y(n812) );
  AO22X1_LVT U711 ( .A1(I1[32]), .A2(I2[32]), .A3(n813), .A4(n814), .Y(n809)
         );
  OR2X1_LVT U712 ( .A1(I1[32]), .A2(I2[32]), .Y(n814) );
  OA22X1_LVT U713 ( .A1(I1[32]), .A2(I2[32]), .A3(I1[31]), .A4(I2[31]), .Y(
        n810) );
  FADDX1_LVT U714 ( .A(I1[32]), .B(I2[32]), .CI(n815), .S(O1[32]) );
  AO221X1_LVT U715 ( .A1(n708), .A2(I1[31]), .A3(n708), .A4(I2[31]), .A5(n813), 
        .Y(n815) );
  AND2X1_LVT U716 ( .A1(I1[31]), .A2(I2[31]), .Y(n813) );
  FADDX1_LVT U717 ( .A(I1[31]), .B(I2[31]), .CI(n708), .S(O1[31]) );
  AO221X1_LVT U718 ( .A1(n816), .A2(n817), .A3(n816), .A4(n818), .A5(n819), 
        .Y(n708) );
  AO221X1_LVT U719 ( .A1(n820), .A2(n821), .A3(n822), .A4(n823), .A5(n824), 
        .Y(n819) );
  AO22X1_LVT U720 ( .A1(I1[30]), .A2(I2[30]), .A3(n825), .A4(n826), .Y(n824)
         );
  OR2X1_LVT U721 ( .A1(I2[30]), .A2(I1[30]), .Y(n826) );
  AND2X1_LVT U722 ( .A1(n827), .A2(n828), .Y(n818) );
  AND2X1_LVT U723 ( .A1(n829), .A2(n823), .Y(n816) );
  AND2X1_LVT U724 ( .A1(n820), .A2(n830), .Y(n823) );
  OA22X1_LVT U725 ( .A1(I1[30]), .A2(I2[30]), .A3(I1[29]), .A4(I2[29]), .Y(
        n820) );
  FADDX1_LVT U726 ( .A(I1[30]), .B(I2[30]), .CI(n831), .S(O1[30]) );
  AO221X1_LVT U727 ( .A1(n832), .A2(I1[29]), .A3(n832), .A4(I2[29]), .A5(n825), 
        .Y(n831) );
  AND2X1_LVT U728 ( .A1(I1[29]), .A2(I2[29]), .Y(n825) );
  FADDX1_LVT U729 ( .A(I1[29]), .B(I2[29]), .CI(n832), .S(O1[29]) );
  AO21X1_LVT U730 ( .A1(n830), .A2(n833), .A3(n821), .Y(n832) );
  AO22X1_LVT U731 ( .A1(I1[28]), .A2(I2[28]), .A3(n834), .A4(n835), .Y(n821)
         );
  OR2X1_LVT U732 ( .A1(I1[28]), .A2(I2[28]), .Y(n835) );
  OA22X1_LVT U733 ( .A1(I1[28]), .A2(I2[28]), .A3(I1[27]), .A4(I2[27]), .Y(
        n830) );
  FADDX1_LVT U734 ( .A(I1[28]), .B(I2[28]), .CI(n836), .S(O1[28]) );
  AO221X1_LVT U735 ( .A1(n833), .A2(I1[27]), .A3(n833), .A4(I2[27]), .A5(n834), 
        .Y(n836) );
  AND2X1_LVT U736 ( .A1(I1[27]), .A2(I2[27]), .Y(n834) );
  FADDX1_LVT U737 ( .A(I1[27]), .B(I2[27]), .CI(n833), .S(O1[27]) );
  AO21X1_LVT U738 ( .A1(n829), .A2(n837), .A3(n822), .Y(n833) );
  AO222X1_LVT U739 ( .A1(I1[26]), .A2(I2[26]), .A3(n838), .A4(n839), .A5(n840), 
        .A6(n841), .Y(n822) );
  OR2X1_LVT U740 ( .A1(I2[26]), .A2(I1[26]), .Y(n839) );
  AND2X1_LVT U741 ( .A1(n840), .A2(n842), .Y(n829) );
  OA22X1_LVT U742 ( .A1(I1[26]), .A2(I2[26]), .A3(I1[25]), .A4(I2[25]), .Y(
        n840) );
  FADDX1_LVT U743 ( .A(I1[26]), .B(I2[26]), .CI(n843), .S(O1[26]) );
  AO221X1_LVT U744 ( .A1(n844), .A2(I1[25]), .A3(n844), .A4(I2[25]), .A5(n838), 
        .Y(n843) );
  AND2X1_LVT U745 ( .A1(I1[25]), .A2(I2[25]), .Y(n838) );
  FADDX1_LVT U746 ( .A(I1[25]), .B(I2[25]), .CI(n844), .S(O1[25]) );
  AO21X1_LVT U747 ( .A1(n842), .A2(n837), .A3(n841), .Y(n844) );
  AO22X1_LVT U748 ( .A1(I1[24]), .A2(I2[24]), .A3(n845), .A4(n846), .Y(n841)
         );
  OR2X1_LVT U749 ( .A1(I1[24]), .A2(I2[24]), .Y(n846) );
  OA22X1_LVT U750 ( .A1(I1[24]), .A2(I2[24]), .A3(I1[23]), .A4(I2[23]), .Y(
        n842) );
  FADDX1_LVT U751 ( .A(I1[24]), .B(I2[24]), .CI(n847), .S(O1[24]) );
  AO221X1_LVT U752 ( .A1(n837), .A2(I1[23]), .A3(n837), .A4(I2[23]), .A5(n845), 
        .Y(n847) );
  AND2X1_LVT U753 ( .A1(I1[23]), .A2(I2[23]), .Y(n845) );
  FADDX1_LVT U754 ( .A(I1[23]), .B(I2[23]), .CI(n837), .S(O1[23]) );
  AO21X1_LVT U755 ( .A1(n828), .A2(n827), .A3(n817), .Y(n837) );
  AO221X1_LVT U756 ( .A1(n848), .A2(n849), .A3(n850), .A4(n851), .A5(n852), 
        .Y(n817) );
  AO22X1_LVT U757 ( .A1(I1[22]), .A2(I2[22]), .A3(n853), .A4(n854), .Y(n852)
         );
  OR2X1_LVT U758 ( .A1(I2[22]), .A2(I1[22]), .Y(n854) );
  AND2X1_LVT U759 ( .A1(n855), .A2(n851), .Y(n828) );
  AND2X1_LVT U760 ( .A1(n848), .A2(n856), .Y(n851) );
  OA22X1_LVT U761 ( .A1(I1[22]), .A2(I2[22]), .A3(I1[21]), .A4(I2[21]), .Y(
        n848) );
  FADDX1_LVT U762 ( .A(I1[22]), .B(I2[22]), .CI(n857), .S(O1[22]) );
  AO221X1_LVT U763 ( .A1(n858), .A2(I1[21]), .A3(n858), .A4(I2[21]), .A5(n853), 
        .Y(n857) );
  AND2X1_LVT U764 ( .A1(I1[21]), .A2(I2[21]), .Y(n853) );
  FADDX1_LVT U765 ( .A(I1[21]), .B(I2[21]), .CI(n858), .S(O1[21]) );
  AO21X1_LVT U766 ( .A1(n856), .A2(n859), .A3(n849), .Y(n858) );
  AO22X1_LVT U767 ( .A1(I1[20]), .A2(I2[20]), .A3(n860), .A4(n861), .Y(n849)
         );
  OR2X1_LVT U768 ( .A1(I1[20]), .A2(I2[20]), .Y(n861) );
  OA22X1_LVT U769 ( .A1(I1[20]), .A2(I2[20]), .A3(I1[19]), .A4(I2[19]), .Y(
        n856) );
  FADDX1_LVT U770 ( .A(I1[20]), .B(I2[20]), .CI(n862), .S(O1[20]) );
  AO221X1_LVT U771 ( .A1(n859), .A2(I1[19]), .A3(n859), .A4(I2[19]), .A5(n860), 
        .Y(n862) );
  AND2X1_LVT U772 ( .A1(I1[19]), .A2(I2[19]), .Y(n860) );
  FADDX1_LVT U773 ( .A(I1[19]), .B(I2[19]), .CI(n859), .S(O1[19]) );
  AO21X1_LVT U774 ( .A1(n827), .A2(n855), .A3(n850), .Y(n859) );
  AO222X1_LVT U775 ( .A1(I1[18]), .A2(I2[18]), .A3(n863), .A4(n864), .A5(n865), 
        .A6(n866), .Y(n850) );
  OR2X1_LVT U776 ( .A1(I2[18]), .A2(I1[18]), .Y(n864) );
  AND2X1_LVT U777 ( .A1(n865), .A2(n867), .Y(n855) );
  OA22X1_LVT U778 ( .A1(I1[18]), .A2(I2[18]), .A3(I1[17]), .A4(I2[17]), .Y(
        n865) );
  FADDX1_LVT U779 ( .A(I1[18]), .B(I2[18]), .CI(n868), .S(O1[18]) );
  AO221X1_LVT U780 ( .A1(n869), .A2(I1[17]), .A3(n869), .A4(I2[17]), .A5(n863), 
        .Y(n868) );
  AND2X1_LVT U781 ( .A1(I1[17]), .A2(I2[17]), .Y(n863) );
  FADDX1_LVT U782 ( .A(I1[17]), .B(I2[17]), .CI(n869), .S(O1[17]) );
  AO21X1_LVT U783 ( .A1(n867), .A2(n827), .A3(n866), .Y(n869) );
  AO22X1_LVT U784 ( .A1(I1[16]), .A2(I2[16]), .A3(n870), .A4(n871), .Y(n866)
         );
  OR2X1_LVT U785 ( .A1(I1[16]), .A2(I2[16]), .Y(n871) );
  OA22X1_LVT U786 ( .A1(I1[16]), .A2(I2[16]), .A3(I1[15]), .A4(I2[15]), .Y(
        n867) );
  FADDX1_LVT U787 ( .A(I1[16]), .B(I2[16]), .CI(n872), .S(O1[16]) );
  OA22X1_LVT U788 ( .A1(n827), .A2(n870), .A3(I1[15]), .A4(I2[15]), .Y(n872)
         );
  AND2X1_LVT U789 ( .A1(I1[15]), .A2(I2[15]), .Y(n870) );
  FADDX1_LVT U790 ( .A(n827), .B(I1[15]), .CI(I2[15]), .S(O1[15]) );
  AO221X1_LVT U791 ( .A1(n877), .A2(n878), .A3(n879), .A4(n874), .A5(n880), 
        .Y(n873) );
  AO22X1_LVT U792 ( .A1(I1[14]), .A2(I2[14]), .A3(n881), .A4(n882), .Y(n880)
         );
  OR2X1_LVT U793 ( .A1(I2[14]), .A2(I1[14]), .Y(n882) );
  AND2X1_LVT U794 ( .A1(n877), .A2(n883), .Y(n874) );
  OA22X1_LVT U795 ( .A1(I1[14]), .A2(I2[14]), .A3(I1[13]), .A4(I2[13]), .Y(
        n877) );
  FADDX1_LVT U796 ( .A(I1[14]), .B(I2[14]), .CI(n884), .S(O1[14]) );
  OA22X1_LVT U797 ( .A1(n881), .A2(n885), .A3(I1[13]), .A4(I2[13]), .Y(n884)
         );
  AND2X1_LVT U798 ( .A1(I1[13]), .A2(I2[13]), .Y(n881) );
  FADDX1_LVT U799 ( .A(I1[13]), .B(I2[13]), .CI(n885), .S(O1[13]) );
  AO21X1_LVT U800 ( .A1(n883), .A2(n886), .A3(n878), .Y(n885) );
  AO22X1_LVT U801 ( .A1(I1[12]), .A2(I2[12]), .A3(n887), .A4(n888), .Y(n878)
         );
  OR2X1_LVT U802 ( .A1(I1[12]), .A2(I2[12]), .Y(n888) );
  OA22X1_LVT U803 ( .A1(I1[12]), .A2(I2[12]), .A3(I1[11]), .A4(I2[11]), .Y(
        n883) );
  FADDX1_LVT U804 ( .A(I1[12]), .B(I2[12]), .CI(n889), .S(O1[12]) );
  OA22X1_LVT U805 ( .A1(n887), .A2(n886), .A3(I1[11]), .A4(I2[11]), .Y(n889)
         );
  AND2X1_LVT U806 ( .A1(I1[11]), .A2(I2[11]), .Y(n887) );
  FADDX1_LVT U807 ( .A(I1[11]), .B(I2[11]), .CI(n886), .S(O1[11]) );
  AO21X1_LVT U808 ( .A1(n875), .A2(n876), .A3(n879), .Y(n886) );
  AO222X1_LVT U809 ( .A1(I1[10]), .A2(I2[10]), .A3(n890), .A4(n891), .A5(n892), 
        .A6(n893), .Y(n879) );
  OR2X1_LVT U810 ( .A1(I2[10]), .A2(I1[10]), .Y(n891) );
  AND2X1_LVT U811 ( .A1(n892), .A2(n894), .Y(n875) );
  OA22X1_LVT U812 ( .A1(I1[10]), .A2(I2[10]), .A3(I1[9]), .A4(I2[9]), .Y(n892)
         );
  FADDX1_LVT U813 ( .A(I1[10]), .B(I2[10]), .CI(n895), .S(O1[10]) );
  OA22X1_LVT U814 ( .A1(n890), .A2(n896), .A3(I1[9]), .A4(I2[9]), .Y(n895) );
  AND2X1_LVT U815 ( .A1(I1[9]), .A2(I2[9]), .Y(n890) );
  FADDX1_LVT U816 ( .A(I1[9]), .B(I2[9]), .CI(n896), .S(O1[9]) );
  AO21X1_LVT U817 ( .A1(n894), .A2(n876), .A3(n893), .Y(n896) );
  AO22X1_LVT U818 ( .A1(I1[8]), .A2(I2[8]), .A3(n897), .A4(n898), .Y(n893) );
  OR2X1_LVT U819 ( .A1(I1[8]), .A2(I2[8]), .Y(n898) );
  OA22X1_LVT U820 ( .A1(I1[8]), .A2(I2[8]), .A3(I1[7]), .A4(I2[7]), .Y(n894)
         );
  FADDX1_LVT U821 ( .A(I1[8]), .B(I2[8]), .CI(n899), .S(O1[8]) );
  AO221X1_LVT U822 ( .A1(n876), .A2(I1[7]), .A3(n876), .A4(I2[7]), .A5(n897), 
        .Y(n899) );
  AND2X1_LVT U823 ( .A1(I1[7]), .A2(I2[7]), .Y(n897) );
  FADDX1_LVT U824 ( .A(I1[7]), .B(I2[7]), .CI(n876), .S(O1[7]) );
  AO221X1_LVT U825 ( .A1(n900), .A2(n901), .A3(n900), .A4(n902), .A5(n903), 
        .Y(n876) );
  AO22X1_LVT U826 ( .A1(I1[6]), .A2(I2[6]), .A3(n904), .A4(n905), .Y(n903) );
  OR2X1_LVT U827 ( .A1(I1[6]), .A2(I2[6]), .Y(n905) );
  AND2X1_LVT U828 ( .A1(n906), .A2(n907), .Y(n901) );
  OA22X1_LVT U829 ( .A1(I1[6]), .A2(I2[6]), .A3(I1[5]), .A4(I2[5]), .Y(n900)
         );
  FADDX1_LVT U830 ( .A(I1[6]), .B(I2[6]), .CI(n908), .S(O1[6]) );
  AO221X1_LVT U831 ( .A1(n909), .A2(I1[5]), .A3(n909), .A4(I2[5]), .A5(n904), 
        .Y(n908) );
  AND2X1_LVT U832 ( .A1(I1[5]), .A2(I2[5]), .Y(n904) );
  FADDX1_LVT U833 ( .A(I1[5]), .B(I2[5]), .CI(n909), .S(O1[5]) );
  AO21X1_LVT U834 ( .A1(n907), .A2(n906), .A3(n902), .Y(n909) );
  AO22X1_LVT U835 ( .A1(I1[4]), .A2(I2[4]), .A3(n910), .A4(n911), .Y(n902) );
  OR2X1_LVT U836 ( .A1(I1[4]), .A2(I2[4]), .Y(n911) );
  OA22X1_LVT U837 ( .A1(I1[4]), .A2(I2[4]), .A3(I1[3]), .A4(I2[3]), .Y(n907)
         );
  FADDX1_LVT U838 ( .A(I1[4]), .B(I2[4]), .CI(n912), .S(O1[4]) );
  OA22X1_LVT U839 ( .A1(n906), .A2(n910), .A3(I1[3]), .A4(I2[3]), .Y(n912) );
  AND2X1_LVT U840 ( .A1(I1[3]), .A2(I2[3]), .Y(n910) );
  FADDX1_LVT U841 ( .A(n906), .B(I1[3]), .CI(I2[3]), .S(O1[3]) );
  AO22X1_LVT U842 ( .A1(I1[2]), .A2(I2[2]), .A3(n916), .A4(n914), .Y(n913) );
  OR2X1_LVT U843 ( .A1(I1[2]), .A2(I2[2]), .Y(n914) );
  FADDX1_LVT U844 ( .A(I1[2]), .B(I2[2]), .CI(n917), .S(O1[2]) );
  AO21X1_LVT U845 ( .A1(n442), .A2(n915), .A3(n916), .Y(n917) );
  AND2X1_LVT U846 ( .A1(I2[1]), .A2(I1[1]), .Y(n916) );
  OR2X1_LVT U847 ( .A1(I2[1]), .A2(I1[1]), .Y(n915) );
  FADDX1_LVT U848 ( .A(n442), .B(I2[1]), .CI(I1[1]), .S(O1[1]) );
endmodule


module ALU_DW_rightsh_J40_0 ( A, DATA_TC, SH, B );
  input [64:0] A;
  input [5:0] SH;
  output [64:0] B;
  input DATA_TC;
  wire   n492, n493, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841;

  IBUFFX2_LVT U418 ( .A(n502), .Y(n504) );
  IBUFFX2_LVT U419 ( .A(n506), .Y(n493) );
  IBUFFX2_LVT U420 ( .A(n506), .Y(n508) );
  IBUFFX2_LVT U421 ( .A(n506), .Y(n507) );
  IBUFFX2_LVT U422 ( .A(n502), .Y(n505) );
  IBUFFX2_LVT U423 ( .A(n502), .Y(n503) );
  IBUFFX2_LVT U424 ( .A(n512), .Y(n514) );
  IBUFFX2_LVT U425 ( .A(n512), .Y(n515) );
  IBUFFX2_LVT U426 ( .A(n512), .Y(n513) );
  IBUFFX2_LVT U427 ( .A(n499), .Y(n500) );
  IBUFFX2_LVT U428 ( .A(n499), .Y(n501) );
  IBUFFX4_LVT U429 ( .A(n499), .Y(n495) );
  IBUFFX2_LVT U430 ( .A(n509), .Y(n510) );
  IBUFFX2_LVT U431 ( .A(n509), .Y(n511) );
  IBUFFX4_LVT U432 ( .A(n509), .Y(n492) );
  IBUFFX2_LVT U433 ( .A(n517), .Y(n520) );
  IBUFFX2_LVT U434 ( .A(n517), .Y(n518) );
  NBUFFX4_LVT U435 ( .A(SH[5]), .Y(n499) );
  NBUFFX2_LVT U436 ( .A(SH[4]), .Y(n517) );
  NBUFFX2_LVT U437 ( .A(SH[3]), .Y(n512) );
  INVX1_LVT U438 ( .A(n517), .Y(n519) );
  INVX1_LVT U439 ( .A(n512), .Y(n516) );
  NBUFFX2_LVT U440 ( .A(SH[2]), .Y(n509) );
  NBUFFX2_LVT U441 ( .A(SH[1]), .Y(n506) );
  NBUFFX2_LVT U442 ( .A(SH[0]), .Y(n502) );
  INVX1_LVT U443 ( .A(n517), .Y(n521) );
  NBUFFX2_LVT U444 ( .A(A[64]), .Y(n496) );
  NBUFFX2_LVT U445 ( .A(A[64]), .Y(n497) );
  NBUFFX2_LVT U446 ( .A(A[64]), .Y(n498) );
  AO22X1_LVT U447 ( .A1(n499), .A2(n522), .A3(n495), .A4(n523), .Y(B[9]) );
  AO22X1_LVT U448 ( .A1(n517), .A2(n524), .A3(n518), .A4(n525), .Y(n523) );
  AO22X1_LVT U449 ( .A1(n512), .A2(n526), .A3(n513), .A4(n527), .Y(n525) );
  AO22X1_LVT U450 ( .A1(n499), .A2(n528), .A3(n495), .A4(n529), .Y(B[8]) );
  AO22X1_LVT U451 ( .A1(n517), .A2(n530), .A3(n518), .A4(n531), .Y(n529) );
  AO22X1_LVT U452 ( .A1(n512), .A2(n532), .A3(n514), .A4(n533), .Y(n531) );
  AO22X1_LVT U453 ( .A1(n499), .A2(n534), .A3(n495), .A4(n535), .Y(B[7]) );
  AO22X1_LVT U454 ( .A1(n517), .A2(n536), .A3(n518), .A4(n537), .Y(n535) );
  AO22X1_LVT U455 ( .A1(n512), .A2(n538), .A3(n516), .A4(n539), .Y(n537) );
  AO22X1_LVT U456 ( .A1(n509), .A2(n540), .A3(n492), .A4(n541), .Y(n539) );
  AO22X1_LVT U457 ( .A1(n499), .A2(n542), .A3(n495), .A4(n543), .Y(B[6]) );
  AO22X1_LVT U458 ( .A1(n517), .A2(n544), .A3(n518), .A4(n545), .Y(n543) );
  AO22X1_LVT U459 ( .A1(n512), .A2(n546), .A3(n513), .A4(n547), .Y(n545) );
  AO22X1_LVT U460 ( .A1(n509), .A2(n548), .A3(n492), .A4(n549), .Y(n547) );
  AO22X1_LVT U461 ( .A1(n499), .A2(A[64]), .A3(n495), .A4(n550), .Y(B[63]) );
  AO22X1_LVT U462 ( .A1(n499), .A2(A[64]), .A3(n495), .A4(n551), .Y(B[62]) );
  AO22X1_LVT U463 ( .A1(n499), .A2(A[64]), .A3(n495), .A4(n552), .Y(B[61]) );
  AO22X1_LVT U464 ( .A1(n499), .A2(n498), .A3(n495), .A4(n553), .Y(B[60]) );
  AO22X1_LVT U465 ( .A1(n499), .A2(n554), .A3(n495), .A4(n555), .Y(B[5]) );
  AO22X1_LVT U466 ( .A1(n517), .A2(n556), .A3(n518), .A4(n557), .Y(n555) );
  AO22X1_LVT U467 ( .A1(n512), .A2(n558), .A3(n514), .A4(n559), .Y(n557) );
  AO22X1_LVT U468 ( .A1(n509), .A2(n560), .A3(n511), .A4(n561), .Y(n559) );
  AO22X1_LVT U469 ( .A1(n499), .A2(n498), .A3(n495), .A4(n562), .Y(B[59]) );
  AO22X1_LVT U470 ( .A1(n499), .A2(n498), .A3(n495), .A4(n563), .Y(B[58]) );
  AO22X1_LVT U471 ( .A1(n499), .A2(n498), .A3(n495), .A4(n564), .Y(B[57]) );
  AO22X1_LVT U472 ( .A1(n499), .A2(n498), .A3(n495), .A4(n565), .Y(B[56]) );
  AO22X1_LVT U473 ( .A1(n499), .A2(n498), .A3(n495), .A4(n566), .Y(B[55]) );
  AO22X1_LVT U474 ( .A1(n499), .A2(n498), .A3(n495), .A4(n567), .Y(B[54]) );
  AO22X1_LVT U475 ( .A1(n499), .A2(n498), .A3(n495), .A4(n568), .Y(B[53]) );
  AO22X1_LVT U476 ( .A1(n499), .A2(n498), .A3(n495), .A4(n569), .Y(B[52]) );
  AO22X1_LVT U477 ( .A1(n499), .A2(n498), .A3(n495), .A4(n570), .Y(B[51]) );
  AO22X1_LVT U478 ( .A1(n499), .A2(n498), .A3(n495), .A4(n571), .Y(B[50]) );
  AO22X1_LVT U479 ( .A1(n499), .A2(n572), .A3(n495), .A4(n573), .Y(B[4]) );
  AO22X1_LVT U480 ( .A1(n517), .A2(n574), .A3(n518), .A4(n575), .Y(n573) );
  AO22X1_LVT U481 ( .A1(n512), .A2(n576), .A3(n513), .A4(n577), .Y(n575) );
  AO22X1_LVT U482 ( .A1(n509), .A2(n578), .A3(n492), .A4(n579), .Y(n577) );
  AO22X1_LVT U483 ( .A1(n499), .A2(n498), .A3(n495), .A4(n580), .Y(B[49]) );
  AO22X1_LVT U484 ( .A1(n499), .A2(n498), .A3(n495), .A4(n581), .Y(B[48]) );
  AO22X1_LVT U485 ( .A1(n499), .A2(n498), .A3(n495), .A4(n582), .Y(B[47]) );
  AO22X1_LVT U486 ( .A1(n499), .A2(n498), .A3(n495), .A4(n583), .Y(B[46]) );
  AO22X1_LVT U487 ( .A1(n499), .A2(n498), .A3(n500), .A4(n584), .Y(B[45]) );
  AO22X1_LVT U488 ( .A1(n499), .A2(A[64]), .A3(n500), .A4(n585), .Y(B[44]) );
  AO22X1_LVT U489 ( .A1(n499), .A2(A[64]), .A3(n500), .A4(n586), .Y(B[43]) );
  AO22X1_LVT U490 ( .A1(n499), .A2(n498), .A3(n500), .A4(n587), .Y(B[42]) );
  AO22X1_LVT U491 ( .A1(n499), .A2(A[64]), .A3(n500), .A4(n522), .Y(B[41]) );
  AO22X1_LVT U492 ( .A1(n517), .A2(n588), .A3(n518), .A4(n589), .Y(n522) );
  AO22X1_LVT U493 ( .A1(n499), .A2(A[64]), .A3(n500), .A4(n528), .Y(B[40]) );
  AO22X1_LVT U494 ( .A1(n517), .A2(n590), .A3(n518), .A4(n591), .Y(n528) );
  AO22X1_LVT U495 ( .A1(n499), .A2(n592), .A3(n500), .A4(n593), .Y(B[3]) );
  AO22X1_LVT U496 ( .A1(n517), .A2(n594), .A3(n518), .A4(n595), .Y(n593) );
  AO22X1_LVT U497 ( .A1(n512), .A2(n596), .A3(n514), .A4(n597), .Y(n595) );
  AO22X1_LVT U498 ( .A1(n509), .A2(n541), .A3(n492), .A4(n598), .Y(n597) );
  AO22X1_LVT U499 ( .A1(n506), .A2(n599), .A3(n507), .A4(n600), .Y(n598) );
  AO22X1_LVT U500 ( .A1(n506), .A2(n601), .A3(n507), .A4(n602), .Y(n541) );
  AO22X1_LVT U501 ( .A1(n499), .A2(A[64]), .A3(n500), .A4(n534), .Y(B[39]) );
  AO22X1_LVT U502 ( .A1(n517), .A2(n603), .A3(n518), .A4(n604), .Y(n534) );
  AO22X1_LVT U503 ( .A1(n499), .A2(n498), .A3(n500), .A4(n542), .Y(B[38]) );
  AO22X1_LVT U504 ( .A1(n517), .A2(n605), .A3(n518), .A4(n606), .Y(n542) );
  AO22X1_LVT U505 ( .A1(n499), .A2(A[64]), .A3(n500), .A4(n554), .Y(B[37]) );
  AO22X1_LVT U506 ( .A1(n517), .A2(n607), .A3(n518), .A4(n608), .Y(n554) );
  AO22X1_LVT U507 ( .A1(n499), .A2(n497), .A3(n500), .A4(n572), .Y(B[36]) );
  AO22X1_LVT U508 ( .A1(n517), .A2(n609), .A3(n519), .A4(n610), .Y(n572) );
  AO22X1_LVT U509 ( .A1(n499), .A2(n497), .A3(n500), .A4(n592), .Y(B[35]) );
  AO22X1_LVT U510 ( .A1(n517), .A2(n611), .A3(n519), .A4(n612), .Y(n592) );
  AO22X1_LVT U511 ( .A1(n499), .A2(n497), .A3(n495), .A4(n613), .Y(B[34]) );
  AO22X1_LVT U512 ( .A1(n499), .A2(n497), .A3(n495), .A4(n614), .Y(B[33]) );
  AO22X1_LVT U513 ( .A1(n499), .A2(n497), .A3(n501), .A4(n615), .Y(B[32]) );
  AO22X1_LVT U514 ( .A1(n499), .A2(n550), .A3(n500), .A4(n616), .Y(B[31]) );
  AO22X1_LVT U515 ( .A1(n517), .A2(n617), .A3(n519), .A4(n618), .Y(n616) );
  AO22X1_LVT U516 ( .A1(n517), .A2(n497), .A3(n519), .A4(n619), .Y(n550) );
  AO22X1_LVT U517 ( .A1(n499), .A2(n551), .A3(n495), .A4(n620), .Y(B[30]) );
  AO22X1_LVT U518 ( .A1(n517), .A2(n621), .A3(n519), .A4(n622), .Y(n620) );
  AO22X1_LVT U519 ( .A1(n517), .A2(n497), .A3(n519), .A4(n623), .Y(n551) );
  AO22X1_LVT U520 ( .A1(n499), .A2(n613), .A3(n495), .A4(n624), .Y(B[2]) );
  AO22X1_LVT U521 ( .A1(n517), .A2(n625), .A3(n519), .A4(n626), .Y(n624) );
  AO22X1_LVT U522 ( .A1(n512), .A2(n627), .A3(n516), .A4(n628), .Y(n626) );
  AO22X1_LVT U523 ( .A1(n509), .A2(n549), .A3(n511), .A4(n629), .Y(n628) );
  AO22X1_LVT U524 ( .A1(n506), .A2(n630), .A3(n508), .A4(n631), .Y(n629) );
  AO22X1_LVT U525 ( .A1(n506), .A2(n632), .A3(n508), .A4(n633), .Y(n549) );
  AO22X1_LVT U526 ( .A1(n517), .A2(n634), .A3(n519), .A4(n635), .Y(n613) );
  AO22X1_LVT U527 ( .A1(n499), .A2(n552), .A3(n495), .A4(n636), .Y(B[29]) );
  AO22X1_LVT U528 ( .A1(n517), .A2(n637), .A3(n519), .A4(n638), .Y(n636) );
  AO22X1_LVT U529 ( .A1(n517), .A2(n497), .A3(n519), .A4(n639), .Y(n552) );
  AO22X1_LVT U530 ( .A1(n499), .A2(n553), .A3(n495), .A4(n640), .Y(B[28]) );
  AO22X1_LVT U531 ( .A1(n517), .A2(n641), .A3(n519), .A4(n642), .Y(n640) );
  AO22X1_LVT U532 ( .A1(n517), .A2(n497), .A3(n519), .A4(n643), .Y(n553) );
  AO22X1_LVT U533 ( .A1(n499), .A2(n562), .A3(n495), .A4(n644), .Y(B[27]) );
  AO22X1_LVT U534 ( .A1(n517), .A2(n645), .A3(n520), .A4(n646), .Y(n644) );
  AO22X1_LVT U535 ( .A1(n517), .A2(n497), .A3(n520), .A4(n647), .Y(n562) );
  AO22X1_LVT U536 ( .A1(n499), .A2(n563), .A3(n495), .A4(n648), .Y(B[26]) );
  AO22X1_LVT U537 ( .A1(n517), .A2(n649), .A3(n520), .A4(n650), .Y(n648) );
  AO22X1_LVT U538 ( .A1(n517), .A2(n497), .A3(n520), .A4(n651), .Y(n563) );
  AO22X1_LVT U539 ( .A1(n499), .A2(n564), .A3(n495), .A4(n652), .Y(B[25]) );
  AO22X1_LVT U540 ( .A1(n517), .A2(n589), .A3(n520), .A4(n524), .Y(n652) );
  AO22X1_LVT U541 ( .A1(n512), .A2(n653), .A3(n516), .A4(n654), .Y(n524) );
  AO22X1_LVT U542 ( .A1(n512), .A2(n655), .A3(n513), .A4(n656), .Y(n589) );
  AO22X1_LVT U543 ( .A1(n517), .A2(n497), .A3(n520), .A4(n588), .Y(n564) );
  AO22X1_LVT U544 ( .A1(n512), .A2(n498), .A3(n516), .A4(n657), .Y(n588) );
  AO22X1_LVT U545 ( .A1(n499), .A2(n565), .A3(n495), .A4(n658), .Y(B[24]) );
  AO22X1_LVT U546 ( .A1(n517), .A2(n591), .A3(n520), .A4(n530), .Y(n658) );
  AO22X1_LVT U547 ( .A1(n512), .A2(n659), .A3(n514), .A4(n660), .Y(n530) );
  AO22X1_LVT U548 ( .A1(n512), .A2(n661), .A3(n513), .A4(n662), .Y(n591) );
  AO22X1_LVT U549 ( .A1(n517), .A2(n498), .A3(n520), .A4(n590), .Y(n565) );
  AO22X1_LVT U550 ( .A1(n512), .A2(n498), .A3(n513), .A4(n663), .Y(n590) );
  AO22X1_LVT U551 ( .A1(n499), .A2(n566), .A3(n501), .A4(n664), .Y(B[23]) );
  AO22X1_LVT U552 ( .A1(n517), .A2(n604), .A3(n520), .A4(n536), .Y(n664) );
  AO22X1_LVT U553 ( .A1(n512), .A2(n665), .A3(n513), .A4(n666), .Y(n536) );
  AO22X1_LVT U554 ( .A1(n512), .A2(n667), .A3(n513), .A4(n668), .Y(n604) );
  AO22X1_LVT U555 ( .A1(n517), .A2(n498), .A3(n520), .A4(n603), .Y(n566) );
  AO22X1_LVT U556 ( .A1(n512), .A2(n669), .A3(n513), .A4(n670), .Y(n603) );
  AO22X1_LVT U557 ( .A1(n499), .A2(n567), .A3(n501), .A4(n671), .Y(B[22]) );
  AO22X1_LVT U558 ( .A1(n517), .A2(n606), .A3(n520), .A4(n544), .Y(n671) );
  AO22X1_LVT U559 ( .A1(n512), .A2(n672), .A3(n513), .A4(n673), .Y(n544) );
  AO22X1_LVT U560 ( .A1(n512), .A2(n674), .A3(n513), .A4(n675), .Y(n606) );
  AO22X1_LVT U561 ( .A1(n517), .A2(n498), .A3(n520), .A4(n605), .Y(n567) );
  AO22X1_LVT U562 ( .A1(n512), .A2(n676), .A3(n513), .A4(n677), .Y(n605) );
  AO22X1_LVT U563 ( .A1(n499), .A2(n568), .A3(n501), .A4(n678), .Y(B[21]) );
  AO22X1_LVT U564 ( .A1(n517), .A2(n608), .A3(n520), .A4(n556), .Y(n678) );
  AO22X1_LVT U565 ( .A1(n512), .A2(n679), .A3(n513), .A4(n680), .Y(n556) );
  AO22X1_LVT U566 ( .A1(n512), .A2(n681), .A3(n513), .A4(n682), .Y(n608) );
  AO22X1_LVT U567 ( .A1(n517), .A2(n498), .A3(n518), .A4(n607), .Y(n568) );
  AO22X1_LVT U568 ( .A1(n512), .A2(n683), .A3(n513), .A4(n684), .Y(n607) );
  AO22X1_LVT U569 ( .A1(n499), .A2(n569), .A3(n501), .A4(n685), .Y(B[20]) );
  AO22X1_LVT U570 ( .A1(n517), .A2(n610), .A3(n518), .A4(n574), .Y(n685) );
  AO22X1_LVT U571 ( .A1(n512), .A2(n686), .A3(n513), .A4(n687), .Y(n574) );
  AO22X1_LVT U572 ( .A1(n512), .A2(n688), .A3(n514), .A4(n689), .Y(n610) );
  AO22X1_LVT U573 ( .A1(n517), .A2(n498), .A3(n518), .A4(n609), .Y(n569) );
  AO22X1_LVT U574 ( .A1(n512), .A2(n690), .A3(n514), .A4(n691), .Y(n609) );
  AO22X1_LVT U575 ( .A1(n499), .A2(n614), .A3(n501), .A4(n692), .Y(B[1]) );
  AO22X1_LVT U576 ( .A1(n517), .A2(n693), .A3(n520), .A4(n694), .Y(n692) );
  AO22X1_LVT U577 ( .A1(n512), .A2(n527), .A3(n514), .A4(n695), .Y(n694) );
  AO22X1_LVT U578 ( .A1(n509), .A2(n561), .A3(n492), .A4(n696), .Y(n695) );
  AO22X1_LVT U579 ( .A1(n506), .A2(n600), .A3(n507), .A4(n697), .Y(n696) );
  AO22X1_LVT U580 ( .A1(n502), .A2(A[2]), .A3(n504), .A4(A[1]), .Y(n697) );
  AO22X1_LVT U581 ( .A1(n502), .A2(A[4]), .A3(n504), .A4(A[3]), .Y(n600) );
  AO22X1_LVT U582 ( .A1(n506), .A2(n602), .A3(n508), .A4(n599), .Y(n561) );
  AO22X1_LVT U583 ( .A1(n502), .A2(A[6]), .A3(n504), .A4(A[5]), .Y(n599) );
  AO22X1_LVT U584 ( .A1(n502), .A2(A[8]), .A3(n504), .A4(A[7]), .Y(n602) );
  AO22X1_LVT U585 ( .A1(n509), .A2(n698), .A3(n492), .A4(n560), .Y(n527) );
  AO22X1_LVT U586 ( .A1(n506), .A2(n699), .A3(n507), .A4(n601), .Y(n560) );
  AO22X1_LVT U587 ( .A1(n502), .A2(A[10]), .A3(n504), .A4(A[9]), .Y(n601) );
  AO22X1_LVT U588 ( .A1(n517), .A2(n700), .A3(n520), .A4(n701), .Y(n614) );
  AO22X1_LVT U589 ( .A1(n499), .A2(n570), .A3(n501), .A4(n702), .Y(B[19]) );
  AO22X1_LVT U590 ( .A1(n517), .A2(n612), .A3(n520), .A4(n594), .Y(n702) );
  AO22X1_LVT U591 ( .A1(n512), .A2(n703), .A3(n514), .A4(n704), .Y(n594) );
  AO22X1_LVT U592 ( .A1(n512), .A2(n705), .A3(n514), .A4(n706), .Y(n612) );
  AO22X1_LVT U593 ( .A1(n517), .A2(n498), .A3(n518), .A4(n611), .Y(n570) );
  AO22X1_LVT U594 ( .A1(n512), .A2(n707), .A3(n514), .A4(n708), .Y(n611) );
  AO22X1_LVT U595 ( .A1(n499), .A2(n571), .A3(n501), .A4(n709), .Y(B[18]) );
  AO22X1_LVT U596 ( .A1(n517), .A2(n635), .A3(n520), .A4(n625), .Y(n709) );
  AO22X1_LVT U597 ( .A1(n512), .A2(n710), .A3(n514), .A4(n711), .Y(n625) );
  AO22X1_LVT U598 ( .A1(n512), .A2(n712), .A3(n514), .A4(n713), .Y(n635) );
  AO22X1_LVT U599 ( .A1(n517), .A2(n498), .A3(n518), .A4(n634), .Y(n571) );
  AO22X1_LVT U600 ( .A1(n512), .A2(n714), .A3(n514), .A4(n715), .Y(n634) );
  AO22X1_LVT U601 ( .A1(n499), .A2(n580), .A3(n501), .A4(n716), .Y(B[17]) );
  AO22X1_LVT U602 ( .A1(n517), .A2(n701), .A3(n518), .A4(n693), .Y(n716) );
  AO22X1_LVT U603 ( .A1(n512), .A2(n654), .A3(n514), .A4(n526), .Y(n693) );
  AO22X1_LVT U604 ( .A1(n509), .A2(n717), .A3(n511), .A4(n718), .Y(n526) );
  AO22X1_LVT U605 ( .A1(n509), .A2(n719), .A3(n492), .A4(n720), .Y(n654) );
  AO22X1_LVT U606 ( .A1(n512), .A2(n656), .A3(n514), .A4(n653), .Y(n701) );
  AO22X1_LVT U607 ( .A1(n509), .A2(n721), .A3(n492), .A4(n722), .Y(n653) );
  AO22X1_LVT U608 ( .A1(n509), .A2(n723), .A3(n492), .A4(n724), .Y(n656) );
  AO22X1_LVT U609 ( .A1(n517), .A2(n498), .A3(n518), .A4(n700), .Y(n580) );
  AO22X1_LVT U610 ( .A1(n512), .A2(n657), .A3(n514), .A4(n655), .Y(n700) );
  AO22X1_LVT U611 ( .A1(n509), .A2(n725), .A3(n510), .A4(n726), .Y(n655) );
  AO22X1_LVT U612 ( .A1(n509), .A2(n727), .A3(n510), .A4(n728), .Y(n657) );
  AO22X1_LVT U613 ( .A1(n499), .A2(n581), .A3(n501), .A4(n729), .Y(B[16]) );
  AO22X1_LVT U614 ( .A1(n517), .A2(n730), .A3(n520), .A4(n731), .Y(n729) );
  AO22X1_LVT U615 ( .A1(n517), .A2(n498), .A3(n520), .A4(n732), .Y(n581) );
  AO22X1_LVT U616 ( .A1(n499), .A2(n582), .A3(n501), .A4(n733), .Y(B[15]) );
  AO22X1_LVT U617 ( .A1(n517), .A2(n618), .A3(n518), .A4(n734), .Y(n733) );
  AO22X1_LVT U618 ( .A1(n512), .A2(n666), .A3(n515), .A4(n538), .Y(n734) );
  AO22X1_LVT U619 ( .A1(n509), .A2(n735), .A3(n510), .A4(n736), .Y(n538) );
  AO22X1_LVT U620 ( .A1(n509), .A2(n737), .A3(n510), .A4(n738), .Y(n666) );
  AO22X1_LVT U621 ( .A1(n512), .A2(n668), .A3(n515), .A4(n665), .Y(n618) );
  AO22X1_LVT U622 ( .A1(n509), .A2(n739), .A3(n510), .A4(n740), .Y(n665) );
  AO22X1_LVT U623 ( .A1(n509), .A2(n741), .A3(n510), .A4(n742), .Y(n668) );
  AO22X1_LVT U624 ( .A1(n517), .A2(n619), .A3(n518), .A4(n617), .Y(n582) );
  AO22X1_LVT U625 ( .A1(n512), .A2(n670), .A3(n515), .A4(n667), .Y(n617) );
  AO22X1_LVT U626 ( .A1(n509), .A2(n743), .A3(n510), .A4(n744), .Y(n667) );
  AO22X1_LVT U627 ( .A1(n509), .A2(n745), .A3(n510), .A4(n746), .Y(n670) );
  AO22X1_LVT U628 ( .A1(n512), .A2(n497), .A3(n515), .A4(n669), .Y(n619) );
  AO22X1_LVT U629 ( .A1(n509), .A2(n496), .A3(n510), .A4(n747), .Y(n669) );
  AO22X1_LVT U630 ( .A1(n499), .A2(n583), .A3(n501), .A4(n748), .Y(B[14]) );
  AO22X1_LVT U631 ( .A1(n517), .A2(n622), .A3(n518), .A4(n749), .Y(n748) );
  AO22X1_LVT U632 ( .A1(n512), .A2(n673), .A3(n515), .A4(n546), .Y(n749) );
  AO22X1_LVT U633 ( .A1(n509), .A2(n750), .A3(n510), .A4(n751), .Y(n546) );
  AO22X1_LVT U634 ( .A1(n509), .A2(n752), .A3(n510), .A4(n753), .Y(n673) );
  AO22X1_LVT U635 ( .A1(n512), .A2(n675), .A3(n515), .A4(n672), .Y(n622) );
  AO22X1_LVT U636 ( .A1(n509), .A2(n754), .A3(n510), .A4(n755), .Y(n672) );
  AO22X1_LVT U637 ( .A1(n509), .A2(n756), .A3(n511), .A4(n757), .Y(n675) );
  AO22X1_LVT U638 ( .A1(n517), .A2(n623), .A3(n520), .A4(n621), .Y(n583) );
  AO22X1_LVT U639 ( .A1(n512), .A2(n677), .A3(n515), .A4(n674), .Y(n621) );
  AO22X1_LVT U640 ( .A1(n509), .A2(n758), .A3(n511), .A4(n759), .Y(n674) );
  AO22X1_LVT U641 ( .A1(n509), .A2(n760), .A3(n511), .A4(n761), .Y(n677) );
  AO22X1_LVT U642 ( .A1(n512), .A2(n496), .A3(n515), .A4(n676), .Y(n623) );
  AO22X1_LVT U643 ( .A1(n509), .A2(n496), .A3(n511), .A4(n762), .Y(n676) );
  AO22X1_LVT U644 ( .A1(n499), .A2(n584), .A3(n501), .A4(n763), .Y(B[13]) );
  AO22X1_LVT U645 ( .A1(n517), .A2(n638), .A3(n520), .A4(n764), .Y(n763) );
  AO22X1_LVT U646 ( .A1(n512), .A2(n680), .A3(n515), .A4(n558), .Y(n764) );
  AO22X1_LVT U647 ( .A1(n509), .A2(n718), .A3(n511), .A4(n698), .Y(n558) );
  AO22X1_LVT U648 ( .A1(n506), .A2(n765), .A3(n508), .A4(n766), .Y(n698) );
  AO22X1_LVT U649 ( .A1(n506), .A2(n767), .A3(n507), .A4(n768), .Y(n718) );
  AO22X1_LVT U650 ( .A1(n509), .A2(n720), .A3(n511), .A4(n717), .Y(n680) );
  AO22X1_LVT U651 ( .A1(n506), .A2(n769), .A3(n508), .A4(n770), .Y(n717) );
  AO22X1_LVT U652 ( .A1(n506), .A2(n771), .A3(n507), .A4(n772), .Y(n720) );
  AO22X1_LVT U653 ( .A1(n512), .A2(n682), .A3(n515), .A4(n679), .Y(n638) );
  AO22X1_LVT U654 ( .A1(n509), .A2(n722), .A3(n511), .A4(n719), .Y(n679) );
  AO22X1_LVT U655 ( .A1(n506), .A2(n773), .A3(n507), .A4(n774), .Y(n719) );
  AO22X1_LVT U656 ( .A1(n506), .A2(n775), .A3(n507), .A4(n776), .Y(n722) );
  AO22X1_LVT U657 ( .A1(n509), .A2(n724), .A3(n511), .A4(n721), .Y(n682) );
  AO22X1_LVT U658 ( .A1(n506), .A2(n777), .A3(n507), .A4(n778), .Y(n721) );
  AO22X1_LVT U659 ( .A1(n506), .A2(n779), .A3(n507), .A4(n780), .Y(n724) );
  AO22X1_LVT U660 ( .A1(n517), .A2(n639), .A3(n520), .A4(n637), .Y(n584) );
  AO22X1_LVT U661 ( .A1(n512), .A2(n684), .A3(n515), .A4(n681), .Y(n637) );
  AO22X1_LVT U662 ( .A1(n509), .A2(n726), .A3(n511), .A4(n723), .Y(n681) );
  AO22X1_LVT U663 ( .A1(n506), .A2(n781), .A3(n507), .A4(n782), .Y(n723) );
  AO22X1_LVT U664 ( .A1(n506), .A2(n783), .A3(n507), .A4(n784), .Y(n726) );
  AO22X1_LVT U665 ( .A1(n509), .A2(n728), .A3(n511), .A4(n725), .Y(n684) );
  AO22X1_LVT U666 ( .A1(n506), .A2(n785), .A3(n507), .A4(n786), .Y(n725) );
  AO22X1_LVT U667 ( .A1(n506), .A2(n787), .A3(n507), .A4(n788), .Y(n728) );
  AO22X1_LVT U668 ( .A1(n512), .A2(n496), .A3(n515), .A4(n683), .Y(n639) );
  AO22X1_LVT U669 ( .A1(n509), .A2(n496), .A3(n511), .A4(n727), .Y(n683) );
  AO22X1_LVT U670 ( .A1(n506), .A2(n789), .A3(n507), .A4(n790), .Y(n727) );
  AO22X1_LVT U671 ( .A1(n499), .A2(n585), .A3(n495), .A4(n791), .Y(B[12]) );
  AO22X1_LVT U672 ( .A1(n517), .A2(n642), .A3(n520), .A4(n792), .Y(n791) );
  AO22X1_LVT U673 ( .A1(n512), .A2(n687), .A3(n516), .A4(n576), .Y(n792) );
  AO22X1_LVT U674 ( .A1(n509), .A2(n793), .A3(n511), .A4(n794), .Y(n576) );
  AO22X1_LVT U675 ( .A1(n509), .A2(n795), .A3(n492), .A4(n796), .Y(n687) );
  AO22X1_LVT U676 ( .A1(n512), .A2(n689), .A3(n516), .A4(n686), .Y(n642) );
  AO22X1_LVT U677 ( .A1(n509), .A2(n797), .A3(n492), .A4(n798), .Y(n686) );
  AO22X1_LVT U678 ( .A1(n509), .A2(n799), .A3(n492), .A4(n800), .Y(n689) );
  AO22X1_LVT U679 ( .A1(n517), .A2(n643), .A3(n520), .A4(n641), .Y(n585) );
  AO22X1_LVT U680 ( .A1(n512), .A2(n691), .A3(n516), .A4(n688), .Y(n641) );
  AO22X1_LVT U681 ( .A1(n509), .A2(n801), .A3(n492), .A4(n802), .Y(n688) );
  AO22X1_LVT U682 ( .A1(n509), .A2(n803), .A3(n492), .A4(n804), .Y(n691) );
  AO22X1_LVT U683 ( .A1(n512), .A2(n496), .A3(n516), .A4(n690), .Y(n643) );
  AO22X1_LVT U684 ( .A1(n509), .A2(n496), .A3(n492), .A4(n805), .Y(n690) );
  AO22X1_LVT U685 ( .A1(n499), .A2(n586), .A3(n501), .A4(n806), .Y(B[11]) );
  AO22X1_LVT U686 ( .A1(n517), .A2(n646), .A3(n518), .A4(n807), .Y(n806) );
  AO22X1_LVT U687 ( .A1(n512), .A2(n704), .A3(n516), .A4(n596), .Y(n807) );
  AO22X1_LVT U688 ( .A1(n509), .A2(n736), .A3(n492), .A4(n540), .Y(n596) );
  AO22X1_LVT U689 ( .A1(n506), .A2(n766), .A3(n507), .A4(n699), .Y(n540) );
  AO22X1_LVT U690 ( .A1(n502), .A2(A[12]), .A3(n504), .A4(A[11]), .Y(n699) );
  AO22X1_LVT U691 ( .A1(n502), .A2(A[14]), .A3(n504), .A4(A[13]), .Y(n766) );
  AO22X1_LVT U692 ( .A1(n506), .A2(n768), .A3(n507), .A4(n765), .Y(n736) );
  AO22X1_LVT U693 ( .A1(n502), .A2(A[16]), .A3(n504), .A4(A[15]), .Y(n765) );
  AO22X1_LVT U694 ( .A1(n502), .A2(A[18]), .A3(n504), .A4(A[17]), .Y(n768) );
  AO22X1_LVT U695 ( .A1(n509), .A2(n738), .A3(n492), .A4(n735), .Y(n704) );
  AO22X1_LVT U696 ( .A1(n506), .A2(n770), .A3(n507), .A4(n767), .Y(n735) );
  AO22X1_LVT U697 ( .A1(n502), .A2(A[20]), .A3(n504), .A4(A[19]), .Y(n767) );
  AO22X1_LVT U698 ( .A1(n502), .A2(A[22]), .A3(n504), .A4(A[21]), .Y(n770) );
  AO22X1_LVT U699 ( .A1(n506), .A2(n772), .A3(n507), .A4(n769), .Y(n738) );
  AO22X1_LVT U700 ( .A1(n502), .A2(A[24]), .A3(n504), .A4(A[23]), .Y(n769) );
  AO22X1_LVT U701 ( .A1(n502), .A2(A[26]), .A3(n503), .A4(A[25]), .Y(n772) );
  AO22X1_LVT U702 ( .A1(n512), .A2(n706), .A3(n516), .A4(n703), .Y(n646) );
  AO22X1_LVT U703 ( .A1(n509), .A2(n740), .A3(n492), .A4(n737), .Y(n703) );
  AO22X1_LVT U704 ( .A1(n506), .A2(n774), .A3(n507), .A4(n771), .Y(n737) );
  AO22X1_LVT U705 ( .A1(n502), .A2(A[28]), .A3(n503), .A4(A[27]), .Y(n771) );
  AO22X1_LVT U706 ( .A1(n502), .A2(A[30]), .A3(n503), .A4(A[29]), .Y(n774) );
  AO22X1_LVT U707 ( .A1(n506), .A2(n776), .A3(n493), .A4(n773), .Y(n740) );
  AO22X1_LVT U708 ( .A1(n502), .A2(A[32]), .A3(n503), .A4(A[31]), .Y(n773) );
  AO22X1_LVT U709 ( .A1(n502), .A2(A[34]), .A3(n503), .A4(A[33]), .Y(n776) );
  AO22X1_LVT U710 ( .A1(n509), .A2(n742), .A3(n492), .A4(n739), .Y(n706) );
  AO22X1_LVT U711 ( .A1(n506), .A2(n778), .A3(n493), .A4(n775), .Y(n739) );
  AO22X1_LVT U712 ( .A1(n502), .A2(A[36]), .A3(n503), .A4(A[35]), .Y(n775) );
  AO22X1_LVT U713 ( .A1(n502), .A2(A[38]), .A3(n503), .A4(A[37]), .Y(n778) );
  AO22X1_LVT U714 ( .A1(n506), .A2(n780), .A3(n507), .A4(n777), .Y(n742) );
  AO22X1_LVT U715 ( .A1(n502), .A2(A[40]), .A3(n503), .A4(A[39]), .Y(n777) );
  AO22X1_LVT U716 ( .A1(n502), .A2(A[42]), .A3(n503), .A4(A[41]), .Y(n780) );
  AO22X1_LVT U717 ( .A1(n517), .A2(n647), .A3(n518), .A4(n645), .Y(n586) );
  AO22X1_LVT U718 ( .A1(n512), .A2(n708), .A3(n516), .A4(n705), .Y(n645) );
  AO22X1_LVT U719 ( .A1(n509), .A2(n744), .A3(n492), .A4(n741), .Y(n705) );
  AO22X1_LVT U720 ( .A1(n506), .A2(n782), .A3(n508), .A4(n779), .Y(n741) );
  AO22X1_LVT U721 ( .A1(n502), .A2(A[44]), .A3(n503), .A4(A[43]), .Y(n779) );
  AO22X1_LVT U722 ( .A1(n502), .A2(A[46]), .A3(n503), .A4(A[45]), .Y(n782) );
  AO22X1_LVT U723 ( .A1(n506), .A2(n784), .A3(n508), .A4(n781), .Y(n744) );
  AO22X1_LVT U724 ( .A1(n502), .A2(A[48]), .A3(n503), .A4(A[47]), .Y(n781) );
  AO22X1_LVT U725 ( .A1(n502), .A2(A[50]), .A3(n505), .A4(A[49]), .Y(n784) );
  AO22X1_LVT U726 ( .A1(n509), .A2(n746), .A3(n492), .A4(n743), .Y(n708) );
  AO22X1_LVT U727 ( .A1(n506), .A2(n786), .A3(n493), .A4(n783), .Y(n743) );
  AO22X1_LVT U728 ( .A1(n502), .A2(A[52]), .A3(n503), .A4(A[51]), .Y(n783) );
  AO22X1_LVT U729 ( .A1(n502), .A2(A[54]), .A3(n503), .A4(A[53]), .Y(n786) );
  AO22X1_LVT U730 ( .A1(n506), .A2(n788), .A3(n508), .A4(n785), .Y(n746) );
  AO22X1_LVT U731 ( .A1(n502), .A2(A[56]), .A3(n505), .A4(A[55]), .Y(n785) );
  AO22X1_LVT U732 ( .A1(n502), .A2(A[58]), .A3(n503), .A4(A[57]), .Y(n788) );
  AO22X1_LVT U733 ( .A1(n512), .A2(n496), .A3(n516), .A4(n707), .Y(n647) );
  AO22X1_LVT U734 ( .A1(n509), .A2(n747), .A3(n492), .A4(n745), .Y(n707) );
  AO22X1_LVT U735 ( .A1(n506), .A2(n790), .A3(n493), .A4(n787), .Y(n745) );
  AO22X1_LVT U736 ( .A1(n502), .A2(A[60]), .A3(n503), .A4(A[59]), .Y(n787) );
  AO22X1_LVT U737 ( .A1(n502), .A2(A[62]), .A3(n505), .A4(A[61]), .Y(n790) );
  AO22X1_LVT U738 ( .A1(n506), .A2(n496), .A3(n507), .A4(n789), .Y(n747) );
  AO22X1_LVT U739 ( .A1(n502), .A2(n496), .A3(n505), .A4(A[63]), .Y(n789) );
  AO22X1_LVT U740 ( .A1(n499), .A2(n587), .A3(n501), .A4(n808), .Y(B[10]) );
  AO22X1_LVT U741 ( .A1(n517), .A2(n650), .A3(n521), .A4(n809), .Y(n808) );
  AO22X1_LVT U742 ( .A1(n512), .A2(n711), .A3(n516), .A4(n627), .Y(n809) );
  AO22X1_LVT U743 ( .A1(n509), .A2(n751), .A3(n492), .A4(n548), .Y(n627) );
  AO22X1_LVT U744 ( .A1(n506), .A2(n810), .A3(n507), .A4(n811), .Y(n548) );
  AO22X1_LVT U745 ( .A1(n506), .A2(n812), .A3(n508), .A4(n813), .Y(n751) );
  AO22X1_LVT U746 ( .A1(n509), .A2(n753), .A3(n492), .A4(n750), .Y(n711) );
  AO22X1_LVT U747 ( .A1(n506), .A2(n814), .A3(n508), .A4(n815), .Y(n750) );
  AO22X1_LVT U748 ( .A1(n506), .A2(n816), .A3(n508), .A4(n817), .Y(n753) );
  AO22X1_LVT U749 ( .A1(n512), .A2(n713), .A3(n516), .A4(n710), .Y(n650) );
  AO22X1_LVT U750 ( .A1(n509), .A2(n755), .A3(n492), .A4(n752), .Y(n710) );
  AO22X1_LVT U751 ( .A1(n506), .A2(n818), .A3(n508), .A4(n819), .Y(n752) );
  AO22X1_LVT U752 ( .A1(n506), .A2(n820), .A3(n508), .A4(n821), .Y(n755) );
  AO22X1_LVT U753 ( .A1(n509), .A2(n757), .A3(n492), .A4(n754), .Y(n713) );
  AO22X1_LVT U754 ( .A1(n506), .A2(n822), .A3(n508), .A4(n823), .Y(n754) );
  AO22X1_LVT U755 ( .A1(n506), .A2(n824), .A3(n508), .A4(n825), .Y(n757) );
  AO22X1_LVT U756 ( .A1(n517), .A2(n651), .A3(n521), .A4(n649), .Y(n587) );
  AO22X1_LVT U757 ( .A1(n512), .A2(n715), .A3(n516), .A4(n712), .Y(n649) );
  AO22X1_LVT U758 ( .A1(n509), .A2(n759), .A3(n492), .A4(n756), .Y(n712) );
  AO22X1_LVT U759 ( .A1(n506), .A2(n826), .A3(n508), .A4(n827), .Y(n756) );
  AO22X1_LVT U760 ( .A1(n506), .A2(n828), .A3(n508), .A4(n829), .Y(n759) );
  AO22X1_LVT U761 ( .A1(n509), .A2(n761), .A3(n492), .A4(n758), .Y(n715) );
  AO22X1_LVT U762 ( .A1(n506), .A2(n830), .A3(n508), .A4(n831), .Y(n758) );
  AO22X1_LVT U763 ( .A1(n506), .A2(n832), .A3(n508), .A4(n833), .Y(n761) );
  AO22X1_LVT U764 ( .A1(n512), .A2(n496), .A3(n516), .A4(n714), .Y(n651) );
  AO22X1_LVT U765 ( .A1(n509), .A2(n762), .A3(n492), .A4(n760), .Y(n714) );
  AO22X1_LVT U766 ( .A1(n506), .A2(n834), .A3(n508), .A4(n835), .Y(n760) );
  AO22X1_LVT U767 ( .A1(n506), .A2(n496), .A3(n508), .A4(n836), .Y(n762) );
  AO22X1_LVT U768 ( .A1(n499), .A2(n615), .A3(n500), .A4(n837), .Y(B[0]) );
  AO22X1_LVT U769 ( .A1(n517), .A2(n731), .A3(n521), .A4(n838), .Y(n837) );
  AO22X1_LVT U770 ( .A1(n512), .A2(n533), .A3(n513), .A4(n839), .Y(n838) );
  AO22X1_LVT U771 ( .A1(n509), .A2(n579), .A3(n492), .A4(n840), .Y(n839) );
  AO22X1_LVT U772 ( .A1(n506), .A2(n631), .A3(n493), .A4(n841), .Y(n840) );
  AO22X1_LVT U773 ( .A1(n502), .A2(A[1]), .A3(n504), .A4(A[0]), .Y(n841) );
  AO22X1_LVT U774 ( .A1(n502), .A2(A[3]), .A3(n504), .A4(A[2]), .Y(n631) );
  AO22X1_LVT U775 ( .A1(n506), .A2(n633), .A3(n493), .A4(n630), .Y(n579) );
  AO22X1_LVT U776 ( .A1(n502), .A2(A[5]), .A3(n504), .A4(A[4]), .Y(n630) );
  AO22X1_LVT U777 ( .A1(n502), .A2(A[7]), .A3(n504), .A4(A[6]), .Y(n633) );
  AO22X1_LVT U778 ( .A1(n509), .A2(n794), .A3(n492), .A4(n578), .Y(n533) );
  AO22X1_LVT U779 ( .A1(n506), .A2(n811), .A3(n493), .A4(n632), .Y(n578) );
  AO22X1_LVT U780 ( .A1(n502), .A2(A[9]), .A3(n504), .A4(A[8]), .Y(n632) );
  AO22X1_LVT U781 ( .A1(n502), .A2(A[11]), .A3(n504), .A4(A[10]), .Y(n811) );
  AO22X1_LVT U782 ( .A1(n506), .A2(n813), .A3(n493), .A4(n810), .Y(n794) );
  AO22X1_LVT U783 ( .A1(n502), .A2(A[13]), .A3(n504), .A4(A[12]), .Y(n810) );
  AO22X1_LVT U784 ( .A1(n502), .A2(A[15]), .A3(n504), .A4(A[14]), .Y(n813) );
  AO22X1_LVT U785 ( .A1(n512), .A2(n660), .A3(n516), .A4(n532), .Y(n731) );
  AO22X1_LVT U786 ( .A1(n509), .A2(n796), .A3(n492), .A4(n793), .Y(n532) );
  AO22X1_LVT U787 ( .A1(n506), .A2(n815), .A3(n493), .A4(n812), .Y(n793) );
  AO22X1_LVT U788 ( .A1(n502), .A2(A[17]), .A3(n504), .A4(A[16]), .Y(n812) );
  AO22X1_LVT U789 ( .A1(n502), .A2(A[19]), .A3(n504), .A4(A[18]), .Y(n815) );
  AO22X1_LVT U790 ( .A1(n506), .A2(n817), .A3(n493), .A4(n814), .Y(n796) );
  AO22X1_LVT U791 ( .A1(n502), .A2(A[21]), .A3(n504), .A4(A[20]), .Y(n814) );
  AO22X1_LVT U792 ( .A1(n502), .A2(A[23]), .A3(n504), .A4(A[22]), .Y(n817) );
  AO22X1_LVT U793 ( .A1(n509), .A2(n798), .A3(n492), .A4(n795), .Y(n660) );
  AO22X1_LVT U794 ( .A1(n506), .A2(n819), .A3(n493), .A4(n816), .Y(n795) );
  AO22X1_LVT U795 ( .A1(n502), .A2(A[25]), .A3(n504), .A4(A[24]), .Y(n816) );
  AO22X1_LVT U796 ( .A1(n502), .A2(A[27]), .A3(n504), .A4(A[26]), .Y(n819) );
  AO22X1_LVT U797 ( .A1(n506), .A2(n821), .A3(n493), .A4(n818), .Y(n798) );
  AO22X1_LVT U798 ( .A1(n502), .A2(A[29]), .A3(n504), .A4(A[28]), .Y(n818) );
  AO22X1_LVT U799 ( .A1(n502), .A2(A[31]), .A3(n504), .A4(A[30]), .Y(n821) );
  AO22X1_LVT U800 ( .A1(n517), .A2(n732), .A3(n521), .A4(n730), .Y(n615) );
  AO22X1_LVT U801 ( .A1(n512), .A2(n662), .A3(n514), .A4(n659), .Y(n730) );
  AO22X1_LVT U802 ( .A1(n509), .A2(n800), .A3(n492), .A4(n797), .Y(n659) );
  AO22X1_LVT U803 ( .A1(n506), .A2(n823), .A3(n493), .A4(n820), .Y(n797) );
  AO22X1_LVT U804 ( .A1(n502), .A2(A[33]), .A3(n505), .A4(A[32]), .Y(n820) );
  AO22X1_LVT U805 ( .A1(n502), .A2(A[35]), .A3(n505), .A4(A[34]), .Y(n823) );
  AO22X1_LVT U806 ( .A1(n506), .A2(n825), .A3(n493), .A4(n822), .Y(n800) );
  AO22X1_LVT U807 ( .A1(n502), .A2(A[37]), .A3(n505), .A4(A[36]), .Y(n822) );
  AO22X1_LVT U808 ( .A1(n502), .A2(A[39]), .A3(n505), .A4(A[38]), .Y(n825) );
  AO22X1_LVT U809 ( .A1(n509), .A2(n802), .A3(n510), .A4(n799), .Y(n662) );
  AO22X1_LVT U810 ( .A1(n506), .A2(n827), .A3(n493), .A4(n824), .Y(n799) );
  AO22X1_LVT U811 ( .A1(n502), .A2(A[41]), .A3(n505), .A4(A[40]), .Y(n824) );
  AO22X1_LVT U812 ( .A1(n502), .A2(A[43]), .A3(n505), .A4(A[42]), .Y(n827) );
  AO22X1_LVT U813 ( .A1(n506), .A2(n829), .A3(n493), .A4(n826), .Y(n802) );
  AO22X1_LVT U814 ( .A1(n502), .A2(A[45]), .A3(n505), .A4(A[44]), .Y(n826) );
  AO22X1_LVT U815 ( .A1(n502), .A2(A[47]), .A3(n505), .A4(A[46]), .Y(n829) );
  AO22X1_LVT U816 ( .A1(n512), .A2(n663), .A3(n515), .A4(n661), .Y(n732) );
  AO22X1_LVT U817 ( .A1(n509), .A2(n804), .A3(n511), .A4(n801), .Y(n661) );
  AO22X1_LVT U818 ( .A1(n506), .A2(n831), .A3(n493), .A4(n828), .Y(n801) );
  AO22X1_LVT U819 ( .A1(n502), .A2(A[49]), .A3(n505), .A4(A[48]), .Y(n828) );
  AO22X1_LVT U820 ( .A1(n502), .A2(A[51]), .A3(n505), .A4(A[50]), .Y(n831) );
  AO22X1_LVT U821 ( .A1(n506), .A2(n833), .A3(n493), .A4(n830), .Y(n804) );
  AO22X1_LVT U822 ( .A1(n502), .A2(A[53]), .A3(n505), .A4(A[52]), .Y(n830) );
  AO22X1_LVT U823 ( .A1(n502), .A2(A[55]), .A3(n505), .A4(A[54]), .Y(n833) );
  AO22X1_LVT U824 ( .A1(n509), .A2(n805), .A3(n510), .A4(n803), .Y(n663) );
  AO22X1_LVT U825 ( .A1(n506), .A2(n835), .A3(n493), .A4(n832), .Y(n803) );
  AO22X1_LVT U826 ( .A1(n502), .A2(A[57]), .A3(n503), .A4(A[56]), .Y(n832) );
  AO22X1_LVT U827 ( .A1(n502), .A2(A[59]), .A3(n503), .A4(A[58]), .Y(n835) );
  AO22X1_LVT U828 ( .A1(n506), .A2(n836), .A3(n493), .A4(n834), .Y(n805) );
  AO22X1_LVT U829 ( .A1(n502), .A2(A[61]), .A3(n503), .A4(A[60]), .Y(n834) );
  AO22X1_LVT U830 ( .A1(n502), .A2(A[63]), .A3(n505), .A4(A[62]), .Y(n836) );
endmodule


module ALU ( io_dw, io_fn, io_in2, io_in1, io_out, io_adder_out, io_cmp_out );
  input [3:0] io_fn;
  input [63:0] io_in2;
  input [63:0] io_in1;
  output [63:0] io_out;
  output [63:0] io_adder_out;
  input io_dw;
  output io_cmp_out;
  wire   n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, shamt_5_, n_T_100_64_, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, SYNOPSYS_UNCONNECTED_1;
  wire   [63:0] in2_inv;
  wire   [63:0] shin;
  wire   [63:0] n_T_101;

  ALU_DP_OP_31J40_124_1870_J40_0 DP_OP_31J40_124_1870 ( .I1(io_in1), .I2(
        in2_inv), .I3(io_fn[3]), .O1({n607, n608, n609, n610, n611, n612, n613, 
        n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
        n626, n627, n628, n629, n630, io_adder_out[39:0]}) );
  ALU_DW_rightsh_J40_0 ashr_7 ( .A({n_T_100_64_, shin}), .DATA_TC(1'b1), .SH({
        shamt_5_, io_in2[4:0]}), .B({SYNOPSYS_UNCONNECTED_1, n_T_101}) );
  AO221X1_LVT U3 ( .A1(1'b1), .A2(n42), .A3(io_adder_out[13]), .A4(n434), .A5(
        n43), .Y(io_out[13]) );
  INVX0_LVT U4 ( .A(io_in1[25]), .Y(n1) );
  INVX0_LVT U5 ( .A(in2_inv[25]), .Y(n2) );
  AO22X1_LVT U6 ( .A1(io_in1[25]), .A2(in2_inv[25]), .A3(n1), .A4(n2), .Y(n392) );
  NAND3X0_LVT U7 ( .A1(io_in1[34]), .A2(io_in2[34]), .A3(n603), .Y(n3) );
  OA21X1_LVT U8 ( .A1(n605), .A2(n452), .A3(n3), .Y(n4) );
  AOI22X1_LVT U9 ( .A1(n124), .A2(n_T_101[34]), .A3(n598), .A4(n_T_101[29]), 
        .Y(n5) );
  NAND2X0_LVT U10 ( .A1(io_adder_out[34]), .A2(n602), .Y(n6) );
  NAND4X0_LVT U11 ( .A1(n115), .A2(n4), .A3(n5), .A4(n6), .Y(io_out[34]) );
  INVX0_LVT U12 ( .A(n_T_101[28]), .Y(n7) );
  OA22X1_LVT U13 ( .A1(n605), .A2(n453), .A3(n123), .A4(n7), .Y(n8) );
  AOI22X1_LVT U14 ( .A1(n602), .A2(io_adder_out[35]), .A3(n124), .A4(
        n_T_101[35]), .Y(n9) );
  NAND3X0_LVT U15 ( .A1(io_in1[35]), .A2(io_in2[35]), .A3(n603), .Y(n10) );
  NAND4X0_LVT U16 ( .A1(n8), .A2(n115), .A3(n9), .A4(n10), .Y(io_out[35]) );
  INVX0_LVT U17 ( .A(io_in1[14]), .Y(n11) );
  INVX0_LVT U18 ( .A(in2_inv[14]), .Y(n12) );
  AO22X1_LVT U19 ( .A1(io_in1[14]), .A2(in2_inv[14]), .A3(n11), .A4(n12), .Y(
        n326) );
  NAND3X0_LVT U20 ( .A1(io_in1[36]), .A2(n603), .A3(io_in2[36]), .Y(n13) );
  OA21X1_LVT U21 ( .A1(n605), .A2(n454), .A3(n13), .Y(n14) );
  AOI22X1_LVT U22 ( .A1(n_T_101[27]), .A2(n598), .A3(n_T_101[36]), .A4(n124), 
        .Y(n15) );
  NAND2X0_LVT U23 ( .A1(n602), .A2(io_adder_out[36]), .Y(n16) );
  NAND4X0_LVT U24 ( .A1(n14), .A2(n115), .A3(n15), .A4(n16), .Y(io_out[36]) );
  INVX0_LVT U25 ( .A(io_in1[12]), .Y(n17) );
  INVX0_LVT U26 ( .A(in2_inv[12]), .Y(n18) );
  AO22X1_LVT U27 ( .A1(io_in1[12]), .A2(in2_inv[12]), .A3(n17), .A4(n18), .Y(
        n319) );
  INVX0_LVT U28 ( .A(io_in1[7]), .Y(n19) );
  INVX0_LVT U29 ( .A(in2_inv[7]), .Y(n20) );
  AO22X1_LVT U30 ( .A1(io_in1[7]), .A2(in2_inv[7]), .A3(n19), .A4(n20), .Y(
        n288) );
  INVX0_LVT U31 ( .A(io_in1[39]), .Y(n21) );
  INVX0_LVT U32 ( .A(in2_inv[39]), .Y(n22) );
  AO22X1_LVT U33 ( .A1(io_in1[39]), .A2(in2_inv[39]), .A3(n21), .A4(n22), .Y(
        n457) );
  NAND3X0_LVT U34 ( .A1(io_in1[37]), .A2(n603), .A3(io_in2[37]), .Y(n23) );
  OA21X1_LVT U35 ( .A1(n605), .A2(n455), .A3(n23), .Y(n24) );
  AOI22X1_LVT U36 ( .A1(n_T_101[37]), .A2(n124), .A3(n_T_101[26]), .A4(n598), 
        .Y(n25) );
  NAND2X0_LVT U37 ( .A1(n602), .A2(io_adder_out[37]), .Y(n26) );
  NAND4X0_LVT U38 ( .A1(n24), .A2(n115), .A3(n25), .A4(n26), .Y(io_out[37]) );
  INVX0_LVT U39 ( .A(io_in1[6]), .Y(n27) );
  INVX0_LVT U40 ( .A(in2_inv[6]), .Y(n28) );
  AO22X1_LVT U41 ( .A1(io_in1[6]), .A2(in2_inv[6]), .A3(n27), .A4(n28), .Y(
        n282) );
  INVX0_LVT U42 ( .A(io_in1[13]), .Y(n29) );
  INVX0_LVT U43 ( .A(in2_inv[13]), .Y(n30) );
  AO22X1_LVT U44 ( .A1(io_in1[13]), .A2(in2_inv[13]), .A3(n29), .A4(n30), .Y(
        n324) );
  INVX0_LVT U45 ( .A(io_in1[63]), .Y(n31) );
  INVX0_LVT U46 ( .A(in2_inv[63]), .Y(n32) );
  AO22X1_LVT U47 ( .A1(io_in1[63]), .A2(in2_inv[63]), .A3(n31), .A4(n32), .Y(
        n604) );
  INVX0_LVT U48 ( .A(io_in1[10]), .Y(n33) );
  INVX0_LVT U49 ( .A(in2_inv[10]), .Y(n34) );
  AO22X1_LVT U50 ( .A1(io_in1[10]), .A2(in2_inv[10]), .A3(n33), .A4(n34), .Y(
        n307) );
  INVX0_LVT U51 ( .A(io_in1[16]), .Y(n35) );
  INVX0_LVT U52 ( .A(in2_inv[16]), .Y(n36) );
  AO22X1_LVT U53 ( .A1(io_in1[16]), .A2(in2_inv[16]), .A3(n35), .A4(n36), .Y(
        n338) );
  NAND3X0_LVT U54 ( .A1(io_in1[38]), .A2(n603), .A3(io_in2[38]), .Y(n37) );
  OA21X1_LVT U55 ( .A1(n605), .A2(n456), .A3(n37), .Y(n38) );
  AOI22X1_LVT U56 ( .A1(n_T_101[25]), .A2(n598), .A3(n_T_101[38]), .A4(n124), 
        .Y(n39) );
  NAND2X0_LVT U57 ( .A1(n602), .A2(io_adder_out[38]), .Y(n40) );
  NAND4X0_LVT U58 ( .A1(n38), .A2(n115), .A3(n39), .A4(n40), .Y(io_out[38]) );
  NAND3X0_LVT U59 ( .A1(io_in1[13]), .A2(io_in2[13]), .A3(n122), .Y(n41) );
  OAI21X1_LVT U60 ( .A1(n423), .A2(n324), .A3(n41), .Y(n42) );
  AO22X1_LVT U61 ( .A1(n441), .A2(n_T_101[50]), .A3(n121), .A4(n_T_101[13]), 
        .Y(n43) );
  INVX0_LVT U63 ( .A(io_in1[15]), .Y(n45) );
  INVX0_LVT U64 ( .A(in2_inv[15]), .Y(n46) );
  AO22X1_LVT U65 ( .A1(io_in1[15]), .A2(in2_inv[15]), .A3(n45), .A4(n46), .Y(
        n331) );
  INVX0_LVT U66 ( .A(io_in1[30]), .Y(n47) );
  INVX0_LVT U67 ( .A(in2_inv[30]), .Y(n48) );
  AO22X1_LVT U68 ( .A1(io_in1[30]), .A2(in2_inv[30]), .A3(n47), .A4(n48), .Y(
        n422) );
  INVX0_LVT U69 ( .A(n_T_101[24]), .Y(n49) );
  OA22X1_LVT U70 ( .A1(n605), .A2(n457), .A3(n123), .A4(n49), .Y(n50) );
  AOI22X1_LVT U71 ( .A1(n602), .A2(io_adder_out[39]), .A3(n124), .A4(
        n_T_101[39]), .Y(n51) );
  NAND3X0_LVT U72 ( .A1(io_in1[39]), .A2(io_in2[39]), .A3(n603), .Y(n52) );
  NAND4X0_LVT U73 ( .A1(n50), .A2(n115), .A3(n51), .A4(n52), .Y(io_out[39]) );
  INVX0_LVT U74 ( .A(io_in1[18]), .Y(n53) );
  INVX0_LVT U75 ( .A(in2_inv[18]), .Y(n54) );
  AO22X1_LVT U76 ( .A1(io_in1[18]), .A2(in2_inv[18]), .A3(n53), .A4(n54), .Y(
        n350) );
  INVX0_LVT U77 ( .A(io_in1[26]), .Y(n55) );
  INVX0_LVT U78 ( .A(in2_inv[26]), .Y(n56) );
  AO22X1_LVT U79 ( .A1(io_in1[26]), .A2(in2_inv[26]), .A3(n55), .A4(n56), .Y(
        n398) );
  INVX0_LVT U80 ( .A(io_in1[35]), .Y(n57) );
  INVX0_LVT U81 ( .A(in2_inv[35]), .Y(n58) );
  AO22X1_LVT U82 ( .A1(io_in1[35]), .A2(in2_inv[35]), .A3(n57), .A4(n58), .Y(
        n453) );
  INVX0_LVT U83 ( .A(n_T_101[0]), .Y(n59) );
  OA22X1_LVT U84 ( .A1(n605), .A2(n604), .A3(n123), .A4(n59), .Y(n60) );
  AOI22X1_LVT U85 ( .A1(n607), .A2(n602), .A3(n124), .A4(n_T_101[63]), .Y(n61)
         );
  NAND3X0_LVT U86 ( .A1(io_in1[63]), .A2(io_in2[63]), .A3(n603), .Y(n62) );
  NAND4X0_LVT U87 ( .A1(n60), .A2(n115), .A3(n61), .A4(n62), .Y(io_out[63]) );
  INVX0_LVT U88 ( .A(io_in1[17]), .Y(n63) );
  INVX0_LVT U89 ( .A(in2_inv[17]), .Y(n64) );
  AO22X1_LVT U90 ( .A1(io_in1[17]), .A2(in2_inv[17]), .A3(n63), .A4(n64), .Y(
        n344) );
  INVX0_LVT U91 ( .A(io_in1[29]), .Y(n65) );
  INVX0_LVT U92 ( .A(in2_inv[29]), .Y(n66) );
  AO22X1_LVT U93 ( .A1(io_in1[29]), .A2(in2_inv[29]), .A3(n65), .A4(n66), .Y(
        n416) );
  INVX0_LVT U94 ( .A(io_in1[32]), .Y(n67) );
  INVX0_LVT U95 ( .A(in2_inv[32]), .Y(n68) );
  AO22X1_LVT U96 ( .A1(io_in1[32]), .A2(in2_inv[32]), .A3(n67), .A4(n68), .Y(
        n437) );
  INVX0_LVT U97 ( .A(io_in1[34]), .Y(n69) );
  INVX0_LVT U98 ( .A(in2_inv[34]), .Y(n70) );
  AO22X1_LVT U99 ( .A1(io_in1[34]), .A2(in2_inv[34]), .A3(n69), .A4(n70), .Y(
        n452) );
  INVX0_LVT U100 ( .A(io_in1[36]), .Y(n71) );
  INVX0_LVT U101 ( .A(in2_inv[36]), .Y(n72) );
  AO22X1_LVT U102 ( .A1(io_in1[36]), .A2(in2_inv[36]), .A3(n71), .A4(n72), .Y(
        n454) );
  INVX0_LVT U103 ( .A(io_in1[37]), .Y(n73) );
  INVX0_LVT U104 ( .A(in2_inv[37]), .Y(n74) );
  AO22X1_LVT U105 ( .A1(io_in1[37]), .A2(in2_inv[37]), .A3(n73), .A4(n74), .Y(
        n455) );
  INVX0_LVT U106 ( .A(io_in1[52]), .Y(n75) );
  INVX0_LVT U107 ( .A(in2_inv[52]), .Y(n76) );
  AO22X1_LVT U108 ( .A1(io_in1[52]), .A2(in2_inv[52]), .A3(n75), .A4(n76), .Y(
        n532) );
  INVX0_LVT U109 ( .A(io_in1[61]), .Y(n77) );
  INVX0_LVT U110 ( .A(in2_inv[61]), .Y(n78) );
  AO22X1_LVT U111 ( .A1(io_in1[61]), .A2(in2_inv[61]), .A3(n77), .A4(n78), .Y(
        n588) );
  INVX0_LVT U112 ( .A(io_in1[19]), .Y(n79) );
  INVX0_LVT U113 ( .A(in2_inv[19]), .Y(n80) );
  AO22X1_LVT U114 ( .A1(io_in1[19]), .A2(in2_inv[19]), .A3(n79), .A4(n80), .Y(
        n356) );
  INVX0_LVT U115 ( .A(io_in1[27]), .Y(n81) );
  INVX0_LVT U116 ( .A(in2_inv[27]), .Y(n82) );
  AO22X1_LVT U117 ( .A1(io_in1[27]), .A2(in2_inv[27]), .A3(n81), .A4(n82), .Y(
        n404) );
  INVX0_LVT U118 ( .A(io_in1[38]), .Y(n83) );
  INVX0_LVT U119 ( .A(in2_inv[38]), .Y(n84) );
  AO22X1_LVT U120 ( .A1(io_in1[38]), .A2(in2_inv[38]), .A3(n83), .A4(n84), .Y(
        n456) );
  INVX0_LVT U121 ( .A(io_in1[47]), .Y(n85) );
  INVX0_LVT U122 ( .A(in2_inv[47]), .Y(n86) );
  AO22X1_LVT U123 ( .A1(io_in1[47]), .A2(in2_inv[47]), .A3(n85), .A4(n86), .Y(
        n501) );
  INVX0_LVT U124 ( .A(io_in1[48]), .Y(n87) );
  INVX0_LVT U125 ( .A(in2_inv[48]), .Y(n88) );
  AO22X1_LVT U126 ( .A1(io_in1[48]), .A2(in2_inv[48]), .A3(n87), .A4(n88), .Y(
        n508) );
  INVX0_LVT U127 ( .A(io_in1[53]), .Y(n89) );
  INVX0_LVT U128 ( .A(in2_inv[53]), .Y(n90) );
  AO22X1_LVT U129 ( .A1(io_in1[53]), .A2(in2_inv[53]), .A3(n89), .A4(n90), .Y(
        n538) );
  INVX0_LVT U130 ( .A(io_in1[33]), .Y(n91) );
  INVX0_LVT U131 ( .A(in2_inv[33]), .Y(n92) );
  AO22X1_LVT U132 ( .A1(io_in1[33]), .A2(in2_inv[33]), .A3(n91), .A4(n92), .Y(
        n446) );
  INVX0_LVT U133 ( .A(io_in1[40]), .Y(n93) );
  INVX0_LVT U134 ( .A(in2_inv[40]), .Y(n94) );
  AO22X1_LVT U135 ( .A1(io_in1[40]), .A2(in2_inv[40]), .A3(n93), .A4(n94), .Y(
        n459) );
  INVX0_LVT U136 ( .A(io_in1[41]), .Y(n95) );
  INVX0_LVT U137 ( .A(in2_inv[41]), .Y(n96) );
  AO22X1_LVT U138 ( .A1(io_in1[41]), .A2(in2_inv[41]), .A3(n95), .A4(n96), .Y(
        n465) );
  INVX0_LVT U139 ( .A(io_in1[42]), .Y(n97) );
  INVX0_LVT U140 ( .A(in2_inv[42]), .Y(n98) );
  AO22X1_LVT U141 ( .A1(io_in1[42]), .A2(in2_inv[42]), .A3(n97), .A4(n98), .Y(
        n471) );
  INVX0_LVT U142 ( .A(io_in1[43]), .Y(n99) );
  INVX0_LVT U143 ( .A(in2_inv[43]), .Y(n100) );
  AO22X1_LVT U144 ( .A1(io_in1[43]), .A2(in2_inv[43]), .A3(n99), .A4(n100), 
        .Y(n477) );
  INVX0_LVT U145 ( .A(io_in1[44]), .Y(n101) );
  INVX0_LVT U146 ( .A(in2_inv[44]), .Y(n102) );
  AO22X1_LVT U147 ( .A1(io_in1[44]), .A2(in2_inv[44]), .A3(n101), .A4(n102), 
        .Y(n483) );
  INVX0_LVT U148 ( .A(io_in1[45]), .Y(n103) );
  INVX0_LVT U149 ( .A(in2_inv[45]), .Y(n104) );
  AO22X1_LVT U150 ( .A1(io_in1[45]), .A2(in2_inv[45]), .A3(n103), .A4(n104), 
        .Y(n489) );
  INVX0_LVT U151 ( .A(io_in1[49]), .Y(n105) );
  INVX0_LVT U152 ( .A(in2_inv[49]), .Y(n106) );
  AO22X1_LVT U153 ( .A1(io_in1[49]), .A2(in2_inv[49]), .A3(n105), .A4(n106), 
        .Y(n514) );
  INVX0_LVT U154 ( .A(io_in1[50]), .Y(n107) );
  INVX0_LVT U155 ( .A(in2_inv[50]), .Y(n108) );
  AO22X1_LVT U156 ( .A1(io_in1[50]), .A2(in2_inv[50]), .A3(n107), .A4(n108), 
        .Y(n520) );
  INVX0_LVT U157 ( .A(io_in1[51]), .Y(n109) );
  INVX0_LVT U158 ( .A(in2_inv[51]), .Y(n110) );
  AO22X1_LVT U159 ( .A1(io_in1[51]), .A2(in2_inv[51]), .A3(n109), .A4(n110), 
        .Y(n526) );
  INVX0_LVT U160 ( .A(io_in1[56]), .Y(n111) );
  INVX0_LVT U161 ( .A(in2_inv[56]), .Y(n112) );
  AO22X1_LVT U162 ( .A1(io_in1[56]), .A2(in2_inv[56]), .A3(n111), .A4(n112), 
        .Y(n556) );
  INVX0_LVT U163 ( .A(io_in1[57]), .Y(n113) );
  INVX0_LVT U164 ( .A(in2_inv[57]), .Y(n114) );
  AO22X1_LVT U165 ( .A1(io_in1[57]), .A2(in2_inv[57]), .A3(n113), .A4(n114), 
        .Y(n562) );
  OR2X4_LVT U166 ( .A1(n121), .A2(n200), .Y(n234) );
  AND2X2_LVT U167 ( .A1(n125), .A2(shin[63]), .Y(n_T_100_64_) );
  INVX1_LVT U168 ( .A(io_in2[9]), .Y(n299) );
  OR2X1_LVT U169 ( .A1(n116), .A2(n200), .Y(n199) );
  INVX1_LVT U170 ( .A(io_in1[3]), .Y(n133) );
  INVX1_LVT U171 ( .A(io_in1[20]), .Y(n153) );
  INVX1_LVT U172 ( .A(io_in1[4]), .Y(n134) );
  INVX1_LVT U173 ( .A(io_in1[21]), .Y(n154) );
  INVX1_LVT U174 ( .A(io_in1[5]), .Y(n130) );
  INVX1_LVT U175 ( .A(io_in1[9]), .Y(n135) );
  INVX1_LVT U176 ( .A(io_in1[23]), .Y(n152) );
  INVX1_LVT U177 ( .A(io_in1[22]), .Y(n151) );
  INVX1_LVT U178 ( .A(io_in1[24]), .Y(n150) );
  INVX1_LVT U179 ( .A(io_in1[0]), .Y(n132) );
  INVX1_LVT U180 ( .A(n598), .Y(n123) );
  INVX0_LVT U181 ( .A(n243), .Y(n238) );
  INVX1_LVT U182 ( .A(io_fn[0]), .Y(n237) );
  INVX1_LVT U183 ( .A(io_fn[2]), .Y(n236) );
  INVX1_LVT U184 ( .A(io_fn[3]), .Y(n126) );
  INVX0_LVT U185 ( .A(n235), .Y(n250) );
  NBUFFX2_LVT U186 ( .A(n606), .Y(n115) );
  INVX0_LVT U187 ( .A(n_T_101[30]), .Y(n448) );
  INVX0_LVT U188 ( .A(n_T_101[32]), .Y(n439) );
  INVX0_LVT U189 ( .A(n_T_101[16]), .Y(n503) );
  INVX0_LVT U190 ( .A(n428), .Y(n131) );
  XOR2X1_LVT U191 ( .A1(in2_inv[31]), .A2(io_in1[31]), .Y(n428) );
  XOR2X1_LVT U192 ( .A1(io_in2[16]), .A2(io_fn[3]), .Y(in2_inv[16]) );
  XOR2X1_LVT U193 ( .A1(io_in2[14]), .A2(n125), .Y(in2_inv[14]) );
  XOR2X1_LVT U194 ( .A1(io_in2[17]), .A2(n125), .Y(in2_inv[17]) );
  XOR2X1_LVT U195 ( .A1(io_in2[15]), .A2(n125), .Y(in2_inv[15]) );
  XOR2X1_LVT U196 ( .A1(io_in2[29]), .A2(n125), .Y(in2_inv[29]) );
  XOR2X1_LVT U197 ( .A1(io_in2[30]), .A2(io_fn[3]), .Y(in2_inv[30]) );
  XOR2X1_LVT U198 ( .A1(io_in2[18]), .A2(n125), .Y(in2_inv[18]) );
  XOR2X1_LVT U199 ( .A1(io_in2[25]), .A2(n125), .Y(in2_inv[25]) );
  XOR2X1_LVT U200 ( .A1(io_in2[19]), .A2(n125), .Y(in2_inv[19]) );
  XOR2X1_LVT U201 ( .A1(io_in2[20]), .A2(n125), .Y(in2_inv[20]) );
  XOR2X1_LVT U202 ( .A1(io_in2[23]), .A2(n125), .Y(in2_inv[23]) );
  XOR2X1_LVT U203 ( .A1(io_in2[24]), .A2(n125), .Y(in2_inv[24]) );
  XOR2X1_LVT U204 ( .A1(io_in2[26]), .A2(n125), .Y(in2_inv[26]) );
  XOR2X1_LVT U205 ( .A1(io_in2[1]), .A2(n125), .Y(in2_inv[1]) );
  XOR2X1_LVT U206 ( .A1(io_in2[2]), .A2(n125), .Y(in2_inv[2]) );
  XOR2X1_LVT U207 ( .A1(io_in2[11]), .A2(n125), .Y(in2_inv[11]) );
  XOR2X1_LVT U208 ( .A1(io_in2[28]), .A2(n125), .Y(in2_inv[28]) );
  XOR2X1_LVT U209 ( .A1(io_in2[27]), .A2(n125), .Y(in2_inv[27]) );
  XOR2X1_LVT U210 ( .A1(io_in2[12]), .A2(n125), .Y(in2_inv[12]) );
  XOR2X1_LVT U211 ( .A1(io_in2[21]), .A2(n125), .Y(in2_inv[21]) );
  XOR2X1_LVT U212 ( .A1(io_in2[22]), .A2(n125), .Y(in2_inv[22]) );
  XOR2X1_LVT U213 ( .A1(io_in2[13]), .A2(n125), .Y(in2_inv[13]) );
  XOR2X1_LVT U214 ( .A1(io_in2[51]), .A2(n125), .Y(in2_inv[51]) );
  XOR2X1_LVT U215 ( .A1(io_in2[63]), .A2(n125), .Y(in2_inv[63]) );
  XOR2X1_LVT U216 ( .A1(io_in2[10]), .A2(n125), .Y(in2_inv[10]) );
  XOR2X1_LVT U217 ( .A1(io_in2[6]), .A2(n125), .Y(in2_inv[6]) );
  XOR2X1_LVT U218 ( .A1(io_in2[44]), .A2(n125), .Y(in2_inv[44]) );
  XOR2X1_LVT U219 ( .A1(io_in2[43]), .A2(n125), .Y(in2_inv[43]) );
  XOR2X1_LVT U220 ( .A1(io_in2[45]), .A2(n125), .Y(in2_inv[45]) );
  XOR2X1_LVT U221 ( .A1(io_in2[46]), .A2(n125), .Y(in2_inv[46]) );
  XOR2X1_LVT U222 ( .A1(io_in2[53]), .A2(n125), .Y(in2_inv[53]) );
  XOR2X1_LVT U223 ( .A1(io_in2[52]), .A2(n125), .Y(in2_inv[52]) );
  XOR2X1_LVT U224 ( .A1(io_in2[54]), .A2(n125), .Y(in2_inv[54]) );
  XOR2X1_LVT U225 ( .A1(io_in2[8]), .A2(n125), .Y(in2_inv[8]) );
  XOR2X1_LVT U226 ( .A1(io_in2[38]), .A2(n125), .Y(in2_inv[38]) );
  XOR2X1_LVT U227 ( .A1(io_in2[39]), .A2(n125), .Y(in2_inv[39]) );
  XOR2X1_LVT U228 ( .A1(io_in2[58]), .A2(n125), .Y(in2_inv[58]) );
  XOR2X1_LVT U229 ( .A1(io_in2[57]), .A2(n125), .Y(in2_inv[57]) );
  XOR2X1_LVT U230 ( .A1(io_in2[0]), .A2(n125), .Y(in2_inv[0]) );
  XOR2X1_LVT U231 ( .A1(io_in2[55]), .A2(n125), .Y(in2_inv[55]) );
  XOR2X1_LVT U232 ( .A1(io_in2[48]), .A2(n125), .Y(in2_inv[48]) );
  XOR2X1_LVT U233 ( .A1(io_in2[56]), .A2(n125), .Y(in2_inv[56]) );
  XOR2X1_LVT U234 ( .A1(io_in2[61]), .A2(n125), .Y(in2_inv[61]) );
  XOR2X1_LVT U235 ( .A1(io_in2[47]), .A2(n125), .Y(in2_inv[47]) );
  XOR2X1_LVT U236 ( .A1(io_in2[62]), .A2(n125), .Y(in2_inv[62]) );
  XOR2X1_LVT U237 ( .A1(io_in2[49]), .A2(n125), .Y(in2_inv[49]) );
  XOR2X1_LVT U238 ( .A1(io_in2[59]), .A2(n125), .Y(in2_inv[59]) );
  XOR2X1_LVT U239 ( .A1(io_in2[50]), .A2(n125), .Y(in2_inv[50]) );
  XOR2X1_LVT U240 ( .A1(io_in2[60]), .A2(n125), .Y(in2_inv[60]) );
  XOR2X1_LVT U241 ( .A1(io_in2[4]), .A2(n125), .Y(in2_inv[4]) );
  XOR2X1_LVT U242 ( .A1(io_in2[35]), .A2(n125), .Y(in2_inv[35]) );
  XOR2X1_LVT U243 ( .A1(io_in2[32]), .A2(n125), .Y(in2_inv[32]) );
  XOR2X1_LVT U244 ( .A1(io_in2[41]), .A2(n125), .Y(in2_inv[41]) );
  XOR2X1_LVT U245 ( .A1(io_in2[31]), .A2(n125), .Y(in2_inv[31]) );
  XOR2X1_LVT U246 ( .A1(io_in2[33]), .A2(n125), .Y(in2_inv[33]) );
  XOR2X1_LVT U247 ( .A1(io_in2[42]), .A2(n125), .Y(in2_inv[42]) );
  XOR2X1_LVT U248 ( .A1(io_in2[34]), .A2(n125), .Y(in2_inv[34]) );
  XOR2X1_LVT U249 ( .A1(io_in2[40]), .A2(n125), .Y(in2_inv[40]) );
  XOR2X1_LVT U250 ( .A1(io_in2[37]), .A2(n125), .Y(in2_inv[37]) );
  XOR2X1_LVT U251 ( .A1(io_in2[36]), .A2(n125), .Y(in2_inv[36]) );
  NOR2X1_LVT U252 ( .A1(io_fn[0]), .A2(io_fn[2]), .Y(n244) );
  XOR2X1_LVT U253 ( .A1(io_in2[5]), .A2(io_fn[3]), .Y(in2_inv[5]) );
  INVX1_LVT U254 ( .A(n435), .Y(n423) );
  AND2X1_LVT U255 ( .A1(n441), .A2(io_dw), .Y(n598) );
  AND2X1_LVT U256 ( .A1(n122), .A2(io_dw), .Y(n603) );
  INVX1_LVT U257 ( .A(n593), .Y(n605) );
  INVX1_LVT U258 ( .A(n118), .Y(n122) );
  INVX1_LVT U259 ( .A(n116), .Y(n121) );
  NAND3X0_LVT U260 ( .A1(n165), .A2(io_fn[0]), .A3(n243), .Y(n116) );
  AND2X1_LVT U261 ( .A1(io_dw), .A2(n434), .Y(n602) );
  AND3X1_LVT U262 ( .A1(n244), .A2(n243), .A3(n242), .Y(n434) );
  INVX1_LVT U263 ( .A(n126), .Y(n125) );
  AND2X1_LVT U264 ( .A1(io_dw), .A2(io_in2[5]), .Y(shamt_5_) );
  NAND2X0_LVT U265 ( .A1(n125), .A2(n241), .Y(n242) );
  XOR2X1_LVT U266 ( .A1(n164), .A2(io_fn[0]), .Y(io_cmp_out) );
  XOR2X1_LVT U267 ( .A1(in2_inv[21]), .A2(n154), .Y(n368) );
  XOR2X1_LVT U268 ( .A1(in2_inv[20]), .A2(n153), .Y(n362) );
  XOR2X1_LVT U269 ( .A1(in2_inv[23]), .A2(n152), .Y(n380) );
  XOR2X1_LVT U270 ( .A1(in2_inv[22]), .A2(n151), .Y(n374) );
  XOR2X1_LVT U271 ( .A1(in2_inv[24]), .A2(n150), .Y(n386) );
  XNOR2X1_LVT U272 ( .A1(in2_inv[8]), .A2(io_in1[8]), .Y(n294) );
  XNOR2X1_LVT U273 ( .A1(in2_inv[28]), .A2(io_in1[28]), .Y(n410) );
  XNOR2X1_LVT U274 ( .A1(in2_inv[11]), .A2(io_in1[11]), .Y(n313) );
  XOR2X1_LVT U275 ( .A1(io_in2[9]), .A2(n135), .Y(n136) );
  XOR2X1_LVT U276 ( .A1(in2_inv[4]), .A2(n134), .Y(n270) );
  XOR2X1_LVT U277 ( .A1(in2_inv[3]), .A2(n133), .Y(n264) );
  XOR2X1_LVT U278 ( .A1(in2_inv[0]), .A2(n132), .Y(n240) );
  XOR2X1_LVT U279 ( .A1(in2_inv[5]), .A2(n130), .Y(n276) );
  XOR2X1_LVT U280 ( .A1(in2_inv[1]), .A2(io_in1[1]), .Y(n251) );
  XOR2X1_LVT U281 ( .A1(in2_inv[2]), .A2(io_in1[2]), .Y(n257) );
  XOR2X1_LVT U282 ( .A1(in2_inv[59]), .A2(io_in1[59]), .Y(n573) );
  XOR2X1_LVT U283 ( .A1(in2_inv[60]), .A2(io_in1[60]), .Y(n580) );
  XOR2X1_LVT U284 ( .A1(in2_inv[62]), .A2(io_in1[62]), .Y(n594) );
  XNOR2X1_LVT U285 ( .A1(in2_inv[58]), .A2(io_in1[58]), .Y(n568) );
  XNOR2X1_LVT U286 ( .A1(in2_inv[55]), .A2(io_in1[55]), .Y(n550) );
  XNOR2X1_LVT U287 ( .A1(in2_inv[54]), .A2(io_in1[54]), .Y(n544) );
  XNOR2X1_LVT U288 ( .A1(in2_inv[46]), .A2(io_in1[46]), .Y(n495) );
  INVX1_LVT U289 ( .A(n117), .Y(n124) );
  XOR2X1_LVT U290 ( .A1(io_in2[3]), .A2(io_fn[3]), .Y(in2_inv[3]) );
  XOR2X1_LVT U291 ( .A1(io_in2[7]), .A2(io_fn[3]), .Y(in2_inv[7]) );
  XOR2X1_LVT U292 ( .A1(io_in2[9]), .A2(io_fn[3]), .Y(in2_inv[9]) );
  NBUFFX2_LVT U293 ( .A(n199), .Y(n119) );
  NBUFFX2_LVT U294 ( .A(n232), .Y(n120) );
  NAND2X0_LVT U295 ( .A1(io_dw), .A2(n121), .Y(n117) );
  NAND2X0_LVT U296 ( .A1(n238), .A2(io_fn[2]), .Y(n118) );
  MUX21X1_LVT U297 ( .A1(n607), .A2(io_fn[1]), .S0(io_in2[63]), .Y(n128) );
  INVX1_LVT U298 ( .A(io_fn[1]), .Y(n241) );
  MUX21X1_LVT U299 ( .A1(n241), .A2(n607), .S0(io_in2[63]), .Y(n127) );
  MUX21X1_LVT U300 ( .A1(n128), .A2(n127), .S0(io_in1[63]), .Y(n129) );
  NAND2X0_LVT U301 ( .A1(n129), .A2(n125), .Y(n235) );
  NAND4X0_LVT U302 ( .A1(n131), .A2(n604), .A3(n288), .A4(n276), .Y(n141) );
  AND4X1_LVT U303 ( .A1(n240), .A2(n264), .A3(n270), .A4(n282), .Y(n139) );
  NAND2X0_LVT U304 ( .A1(n136), .A2(n126), .Y(n137) );
  NOR4X1_LVT U305 ( .A1(n137), .A2(n594), .A3(n580), .A4(n573), .Y(n138) );
  NAND4X0_LVT U306 ( .A1(n139), .A2(n138), .A3(n356), .A4(n422), .Y(n140) );
  NOR4X1_LVT U307 ( .A1(n257), .A2(n251), .A3(n141), .A4(n140), .Y(n162) );
  NAND4X0_LVT U308 ( .A1(n562), .A2(n556), .A3(n538), .A4(n550), .Y(n145) );
  NAND4X0_LVT U309 ( .A1(n532), .A2(n526), .A3(n520), .A4(n514), .Y(n144) );
  NAND4X0_LVT U310 ( .A1(n508), .A2(n501), .A3(n489), .A4(n483), .Y(n143) );
  NAND4X0_LVT U311 ( .A1(n477), .A2(n471), .A3(n465), .A4(n459), .Y(n142) );
  NOR4X1_LVT U312 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .Y(n161) );
  NAND4X0_LVT U313 ( .A1(n588), .A2(n568), .A3(n544), .A4(n495), .Y(n149) );
  NAND4X0_LVT U314 ( .A1(n457), .A2(n456), .A3(n455), .A4(n454), .Y(n148) );
  NAND4X0_LVT U315 ( .A1(n453), .A2(n452), .A3(n446), .A4(n437), .Y(n147) );
  NAND4X0_LVT U316 ( .A1(n326), .A2(n331), .A3(n319), .A4(n324), .Y(n146) );
  NOR4X1_LVT U317 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .Y(n160) );
  NAND4X0_LVT U318 ( .A1(n307), .A2(n313), .A3(n410), .A4(n294), .Y(n158) );
  NAND4X0_LVT U319 ( .A1(n416), .A2(n398), .A3(n404), .A4(n386), .Y(n157) );
  NAND4X0_LVT U320 ( .A1(n392), .A2(n374), .A3(n380), .A4(n362), .Y(n156) );
  NAND4X0_LVT U321 ( .A1(n368), .A2(n350), .A3(n338), .A4(n344), .Y(n155) );
  NOR4X1_LVT U322 ( .A1(n158), .A2(n157), .A3(n156), .A4(n155), .Y(n159) );
  NAND4X0_LVT U323 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .Y(n163) );
  NAND2X0_LVT U324 ( .A1(n235), .A2(n163), .Y(n164) );
  MUX21X1_LVT U325 ( .A1(io_fn[1]), .A2(n126), .S0(io_fn[2]), .Y(n165) );
  NAND2X0_LVT U326 ( .A1(io_fn[1]), .A2(n126), .Y(n243) );
  AOI22X1_LVT U327 ( .A1(io_in1[0]), .A2(n116), .A3(io_in1[63]), .A4(n124), 
        .Y(n167) );
  INVX1_LVT U328 ( .A(io_dw), .Y(n440) );
  AND2X1_LVT U329 ( .A1(n440), .A2(n125), .Y(n166) );
  NAND2X0_LVT U330 ( .A1(io_in1[31]), .A2(n166), .Y(n200) );
  NAND2X0_LVT U331 ( .A1(n167), .A2(n199), .Y(shin[63]) );
  AOI22X1_LVT U332 ( .A1(io_in1[1]), .A2(n116), .A3(io_in1[62]), .A4(n124), 
        .Y(n168) );
  NAND2X0_LVT U333 ( .A1(n199), .A2(n168), .Y(shin[62]) );
  AOI22X1_LVT U334 ( .A1(io_in1[2]), .A2(n116), .A3(io_in1[61]), .A4(n124), 
        .Y(n169) );
  NAND2X0_LVT U335 ( .A1(n119), .A2(n169), .Y(shin[61]) );
  AOI22X1_LVT U336 ( .A1(io_in1[3]), .A2(n116), .A3(io_in1[60]), .A4(n124), 
        .Y(n170) );
  NAND2X0_LVT U337 ( .A1(n119), .A2(n170), .Y(shin[60]) );
  AOI22X1_LVT U338 ( .A1(io_in1[4]), .A2(n116), .A3(io_in1[59]), .A4(n124), 
        .Y(n171) );
  NAND2X0_LVT U339 ( .A1(n119), .A2(n171), .Y(shin[59]) );
  AOI22X1_LVT U340 ( .A1(io_in1[5]), .A2(n116), .A3(io_in1[58]), .A4(n124), 
        .Y(n172) );
  NAND2X0_LVT U341 ( .A1(n119), .A2(n172), .Y(shin[58]) );
  AOI22X1_LVT U342 ( .A1(io_in1[6]), .A2(n116), .A3(io_in1[57]), .A4(n124), 
        .Y(n173) );
  NAND2X0_LVT U343 ( .A1(n199), .A2(n173), .Y(shin[57]) );
  AOI22X1_LVT U344 ( .A1(io_in1[7]), .A2(n116), .A3(io_in1[56]), .A4(n124), 
        .Y(n174) );
  NAND2X0_LVT U345 ( .A1(n119), .A2(n174), .Y(shin[56]) );
  AOI22X1_LVT U346 ( .A1(io_in1[8]), .A2(n116), .A3(io_in1[55]), .A4(n124), 
        .Y(n175) );
  NAND2X0_LVT U347 ( .A1(n199), .A2(n175), .Y(shin[55]) );
  AOI22X1_LVT U348 ( .A1(io_in1[9]), .A2(n116), .A3(io_in1[54]), .A4(n124), 
        .Y(n176) );
  NAND2X0_LVT U349 ( .A1(n199), .A2(n176), .Y(shin[54]) );
  AOI22X1_LVT U350 ( .A1(io_in1[10]), .A2(n116), .A3(io_in1[53]), .A4(n124), 
        .Y(n177) );
  NAND2X0_LVT U351 ( .A1(n199), .A2(n177), .Y(shin[53]) );
  AOI22X1_LVT U352 ( .A1(io_in1[11]), .A2(n116), .A3(io_in1[52]), .A4(n124), 
        .Y(n178) );
  NAND2X0_LVT U353 ( .A1(n199), .A2(n178), .Y(shin[52]) );
  AOI22X1_LVT U354 ( .A1(io_in1[12]), .A2(n116), .A3(io_in1[51]), .A4(n124), 
        .Y(n179) );
  NAND2X0_LVT U355 ( .A1(n199), .A2(n179), .Y(shin[51]) );
  AOI22X1_LVT U356 ( .A1(io_in1[13]), .A2(n116), .A3(io_in1[50]), .A4(n124), 
        .Y(n180) );
  NAND2X0_LVT U357 ( .A1(n199), .A2(n180), .Y(shin[50]) );
  AOI22X1_LVT U358 ( .A1(io_in1[14]), .A2(n116), .A3(io_in1[49]), .A4(n124), 
        .Y(n181) );
  NAND2X0_LVT U359 ( .A1(n199), .A2(n181), .Y(shin[49]) );
  AOI22X1_LVT U360 ( .A1(io_in1[15]), .A2(n116), .A3(io_in1[48]), .A4(n124), 
        .Y(n182) );
  NAND2X0_LVT U361 ( .A1(n199), .A2(n182), .Y(shin[48]) );
  AOI22X1_LVT U362 ( .A1(io_in1[16]), .A2(n116), .A3(io_in1[47]), .A4(n124), 
        .Y(n183) );
  NAND2X0_LVT U363 ( .A1(n199), .A2(n183), .Y(shin[47]) );
  AOI22X1_LVT U364 ( .A1(io_in1[17]), .A2(n116), .A3(io_in1[46]), .A4(n124), 
        .Y(n184) );
  NAND2X0_LVT U365 ( .A1(n199), .A2(n184), .Y(shin[46]) );
  AOI22X1_LVT U366 ( .A1(io_in1[18]), .A2(n116), .A3(io_in1[45]), .A4(n124), 
        .Y(n185) );
  NAND2X0_LVT U367 ( .A1(n199), .A2(n185), .Y(shin[45]) );
  AOI22X1_LVT U368 ( .A1(io_in1[19]), .A2(n116), .A3(io_in1[44]), .A4(n124), 
        .Y(n186) );
  NAND2X0_LVT U369 ( .A1(n199), .A2(n186), .Y(shin[44]) );
  AOI22X1_LVT U370 ( .A1(io_in1[20]), .A2(n116), .A3(io_in1[43]), .A4(n124), 
        .Y(n187) );
  NAND2X0_LVT U371 ( .A1(n119), .A2(n187), .Y(shin[43]) );
  AOI22X1_LVT U372 ( .A1(io_in1[21]), .A2(n116), .A3(io_in1[42]), .A4(n124), 
        .Y(n188) );
  NAND2X0_LVT U373 ( .A1(n119), .A2(n188), .Y(shin[42]) );
  AOI22X1_LVT U374 ( .A1(io_in1[22]), .A2(n116), .A3(io_in1[41]), .A4(n124), 
        .Y(n189) );
  NAND2X0_LVT U375 ( .A1(n119), .A2(n189), .Y(shin[41]) );
  AOI22X1_LVT U376 ( .A1(io_in1[23]), .A2(n116), .A3(io_in1[40]), .A4(n124), 
        .Y(n190) );
  NAND2X0_LVT U377 ( .A1(n119), .A2(n190), .Y(shin[40]) );
  AOI22X1_LVT U378 ( .A1(io_in1[24]), .A2(n116), .A3(io_in1[39]), .A4(n124), 
        .Y(n191) );
  NAND2X0_LVT U379 ( .A1(n119), .A2(n191), .Y(shin[39]) );
  AOI22X1_LVT U380 ( .A1(io_in1[38]), .A2(n124), .A3(io_in1[25]), .A4(n116), 
        .Y(n192) );
  NAND2X0_LVT U381 ( .A1(n119), .A2(n192), .Y(shin[38]) );
  AOI22X1_LVT U382 ( .A1(io_in1[37]), .A2(n124), .A3(io_in1[26]), .A4(n116), 
        .Y(n193) );
  NAND2X0_LVT U383 ( .A1(n119), .A2(n193), .Y(shin[37]) );
  AOI22X1_LVT U384 ( .A1(io_in1[36]), .A2(n124), .A3(io_in1[27]), .A4(n116), 
        .Y(n194) );
  NAND2X0_LVT U385 ( .A1(n119), .A2(n194), .Y(shin[36]) );
  AOI22X1_LVT U386 ( .A1(io_in1[35]), .A2(n124), .A3(io_in1[28]), .A4(n116), 
        .Y(n195) );
  NAND2X0_LVT U387 ( .A1(n119), .A2(n195), .Y(shin[35]) );
  AOI22X1_LVT U388 ( .A1(io_in1[34]), .A2(n124), .A3(io_in1[29]), .A4(n116), 
        .Y(n196) );
  NAND2X0_LVT U389 ( .A1(n119), .A2(n196), .Y(shin[34]) );
  AOI22X1_LVT U390 ( .A1(io_in1[33]), .A2(n124), .A3(io_in1[30]), .A4(n116), 
        .Y(n197) );
  NAND2X0_LVT U391 ( .A1(n119), .A2(n197), .Y(shin[33]) );
  AOI22X1_LVT U392 ( .A1(io_in1[32]), .A2(n124), .A3(io_in1[31]), .A4(n116), 
        .Y(n198) );
  NAND2X0_LVT U393 ( .A1(n119), .A2(n198), .Y(shin[32]) );
  NOR2X0_LVT U394 ( .A1(n440), .A2(n121), .Y(n232) );
  AOI22X1_LVT U395 ( .A1(io_in1[32]), .A2(n120), .A3(n121), .A4(io_in1[31]), 
        .Y(n201) );
  NAND2X0_LVT U396 ( .A1(n234), .A2(n201), .Y(shin[31]) );
  AOI22X1_LVT U397 ( .A1(io_in1[30]), .A2(n121), .A3(io_in1[33]), .A4(n120), 
        .Y(n202) );
  NAND2X0_LVT U398 ( .A1(n234), .A2(n202), .Y(shin[30]) );
  AOI22X1_LVT U399 ( .A1(io_in1[34]), .A2(n120), .A3(n121), .A4(io_in1[29]), 
        .Y(n203) );
  NAND2X0_LVT U400 ( .A1(n234), .A2(n203), .Y(shin[29]) );
  AOI22X1_LVT U401 ( .A1(io_in1[35]), .A2(n120), .A3(n121), .A4(io_in1[28]), 
        .Y(n204) );
  NAND2X0_LVT U402 ( .A1(n234), .A2(n204), .Y(shin[28]) );
  AOI22X1_LVT U403 ( .A1(io_in1[36]), .A2(n120), .A3(n121), .A4(io_in1[27]), 
        .Y(n205) );
  NAND2X0_LVT U404 ( .A1(n234), .A2(n205), .Y(shin[27]) );
  AOI22X1_LVT U405 ( .A1(io_in1[37]), .A2(n120), .A3(n121), .A4(io_in1[26]), 
        .Y(n206) );
  NAND2X0_LVT U406 ( .A1(n234), .A2(n206), .Y(shin[26]) );
  AOI22X1_LVT U407 ( .A1(io_in1[38]), .A2(n120), .A3(n121), .A4(io_in1[25]), 
        .Y(n207) );
  NAND2X0_LVT U408 ( .A1(n234), .A2(n207), .Y(shin[25]) );
  AOI22X1_LVT U409 ( .A1(io_in1[24]), .A2(n121), .A3(io_in1[39]), .A4(n120), 
        .Y(n208) );
  NAND2X0_LVT U410 ( .A1(n234), .A2(n208), .Y(shin[24]) );
  AOI22X1_LVT U411 ( .A1(io_in1[23]), .A2(n121), .A3(io_in1[40]), .A4(n232), 
        .Y(n209) );
  NAND2X0_LVT U412 ( .A1(n234), .A2(n209), .Y(shin[23]) );
  AOI22X1_LVT U413 ( .A1(io_in1[22]), .A2(n121), .A3(io_in1[41]), .A4(n232), 
        .Y(n210) );
  NAND2X0_LVT U414 ( .A1(n234), .A2(n210), .Y(shin[22]) );
  AOI22X1_LVT U415 ( .A1(io_in1[21]), .A2(n121), .A3(io_in1[42]), .A4(n232), 
        .Y(n211) );
  NAND2X0_LVT U416 ( .A1(n234), .A2(n211), .Y(shin[21]) );
  AOI22X1_LVT U417 ( .A1(io_in1[20]), .A2(n121), .A3(io_in1[43]), .A4(n120), 
        .Y(n212) );
  NAND2X0_LVT U418 ( .A1(n234), .A2(n212), .Y(shin[20]) );
  AOI22X1_LVT U419 ( .A1(io_in1[19]), .A2(n121), .A3(io_in1[44]), .A4(n232), 
        .Y(n213) );
  NAND2X0_LVT U420 ( .A1(n234), .A2(n213), .Y(shin[19]) );
  AOI22X1_LVT U421 ( .A1(io_in1[18]), .A2(n121), .A3(io_in1[45]), .A4(n120), 
        .Y(n214) );
  NAND2X0_LVT U422 ( .A1(n234), .A2(n214), .Y(shin[18]) );
  AOI22X1_LVT U423 ( .A1(io_in1[17]), .A2(n121), .A3(io_in1[46]), .A4(n232), 
        .Y(n215) );
  NAND2X0_LVT U424 ( .A1(n234), .A2(n215), .Y(shin[17]) );
  AOI22X1_LVT U425 ( .A1(io_in1[16]), .A2(n121), .A3(io_in1[47]), .A4(n232), 
        .Y(n216) );
  NAND2X0_LVT U426 ( .A1(n234), .A2(n216), .Y(shin[16]) );
  AOI22X1_LVT U427 ( .A1(io_in1[15]), .A2(n121), .A3(io_in1[48]), .A4(n120), 
        .Y(n217) );
  NAND2X0_LVT U428 ( .A1(n234), .A2(n217), .Y(shin[15]) );
  AOI22X1_LVT U429 ( .A1(io_in1[14]), .A2(n121), .A3(io_in1[49]), .A4(n232), 
        .Y(n218) );
  NAND2X0_LVT U430 ( .A1(n234), .A2(n218), .Y(shin[14]) );
  AOI22X1_LVT U431 ( .A1(io_in1[13]), .A2(n121), .A3(io_in1[50]), .A4(n120), 
        .Y(n219) );
  NAND2X0_LVT U432 ( .A1(n234), .A2(n219), .Y(shin[13]) );
  AOI22X1_LVT U433 ( .A1(io_in1[12]), .A2(n121), .A3(io_in1[51]), .A4(n232), 
        .Y(n220) );
  NAND2X0_LVT U434 ( .A1(n234), .A2(n220), .Y(shin[12]) );
  AOI22X1_LVT U435 ( .A1(io_in1[11]), .A2(n121), .A3(io_in1[52]), .A4(n232), 
        .Y(n221) );
  NAND2X0_LVT U436 ( .A1(n234), .A2(n221), .Y(shin[11]) );
  AOI22X1_LVT U437 ( .A1(io_in1[10]), .A2(n121), .A3(io_in1[53]), .A4(n232), 
        .Y(n222) );
  NAND2X0_LVT U438 ( .A1(n234), .A2(n222), .Y(shin[10]) );
  AOI22X1_LVT U439 ( .A1(io_in1[9]), .A2(n121), .A3(io_in1[54]), .A4(n232), 
        .Y(n223) );
  NAND2X0_LVT U440 ( .A1(n234), .A2(n223), .Y(shin[9]) );
  AOI22X1_LVT U441 ( .A1(io_in1[8]), .A2(n121), .A3(io_in1[55]), .A4(n232), 
        .Y(n224) );
  NAND2X0_LVT U442 ( .A1(n234), .A2(n224), .Y(shin[8]) );
  AOI22X1_LVT U443 ( .A1(io_in1[7]), .A2(n121), .A3(io_in1[56]), .A4(n120), 
        .Y(n225) );
  NAND2X0_LVT U444 ( .A1(n234), .A2(n225), .Y(shin[7]) );
  AOI22X1_LVT U445 ( .A1(io_in1[6]), .A2(n121), .A3(io_in1[57]), .A4(n232), 
        .Y(n226) );
  NAND2X0_LVT U446 ( .A1(n234), .A2(n226), .Y(shin[6]) );
  AOI22X1_LVT U447 ( .A1(io_in1[5]), .A2(n121), .A3(io_in1[58]), .A4(n120), 
        .Y(n227) );
  NAND2X0_LVT U448 ( .A1(n234), .A2(n227), .Y(shin[5]) );
  AOI22X1_LVT U449 ( .A1(io_in1[4]), .A2(n121), .A3(io_in1[59]), .A4(n232), 
        .Y(n228) );
  NAND2X0_LVT U450 ( .A1(n234), .A2(n228), .Y(shin[4]) );
  AOI22X1_LVT U451 ( .A1(io_in1[3]), .A2(n121), .A3(io_in1[60]), .A4(n120), 
        .Y(n229) );
  NAND2X0_LVT U452 ( .A1(n234), .A2(n229), .Y(shin[3]) );
  AOI22X1_LVT U453 ( .A1(io_in1[2]), .A2(n121), .A3(io_in1[61]), .A4(n232), 
        .Y(n230) );
  NAND2X0_LVT U454 ( .A1(n234), .A2(n230), .Y(shin[2]) );
  AOI22X1_LVT U455 ( .A1(io_in1[1]), .A2(n121), .A3(io_in1[62]), .A4(n120), 
        .Y(n231) );
  NAND2X0_LVT U456 ( .A1(n234), .A2(n231), .Y(shin[1]) );
  AOI22X1_LVT U457 ( .A1(n121), .A2(io_in1[0]), .A3(io_in1[63]), .A4(n120), 
        .Y(n233) );
  NAND2X0_LVT U458 ( .A1(n234), .A2(n233), .Y(shin[0]) );
  AND4X1_LVT U459 ( .A1(n241), .A2(n236), .A3(n126), .A4(io_fn[0]), .Y(n441)
         );
  NAND2X0_LVT U460 ( .A1(n_T_101[63]), .A2(n441), .Y(n248) );
  AND3X1_LVT U461 ( .A1(n126), .A2(io_fn[2]), .A3(n237), .Y(n435) );
  NAND3X0_LVT U462 ( .A1(io_in2[0]), .A2(n122), .A3(io_in1[0]), .Y(n239) );
  OA21X1_LVT U463 ( .A1(n423), .A2(n240), .A3(n239), .Y(n247) );
  NAND2X0_LVT U464 ( .A1(n_T_101[0]), .A2(n121), .Y(n246) );
  NAND2X0_LVT U465 ( .A1(io_adder_out[0]), .A2(n434), .Y(n245) );
  NAND4X0_LVT U466 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .Y(n249) );
  AO21X1_LVT U467 ( .A1(io_fn[2]), .A2(n250), .A3(n249), .Y(io_out[0]) );
  NAND2X0_LVT U468 ( .A1(n_T_101[62]), .A2(n441), .Y(n255) );
  NAND2X0_LVT U469 ( .A1(io_adder_out[1]), .A2(n434), .Y(n254) );
  NAND2X0_LVT U470 ( .A1(n251), .A2(n435), .Y(n253) );
  NAND3X0_LVT U471 ( .A1(io_in2[1]), .A2(n122), .A3(io_in1[1]), .Y(n252) );
  NAND4X0_LVT U472 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .Y(n256) );
  AO21X1_LVT U473 ( .A1(n121), .A2(n_T_101[1]), .A3(n256), .Y(io_out[1]) );
  NAND2X0_LVT U474 ( .A1(n_T_101[61]), .A2(n441), .Y(n262) );
  AND2X1_LVT U475 ( .A1(io_in1[2]), .A2(n122), .Y(n258) );
  AOI22X1_LVT U476 ( .A1(io_in2[2]), .A2(n258), .A3(n257), .A4(n435), .Y(n261)
         );
  NAND2X0_LVT U477 ( .A1(n_T_101[2]), .A2(n121), .Y(n260) );
  NAND2X0_LVT U478 ( .A1(io_adder_out[2]), .A2(n434), .Y(n259) );
  NAND4X0_LVT U479 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .Y(io_out[2])
         );
  NAND2X0_LVT U480 ( .A1(n_T_101[3]), .A2(n121), .Y(n268) );
  NAND3X0_LVT U481 ( .A1(io_in2[3]), .A2(n122), .A3(io_in1[3]), .Y(n263) );
  OA21X1_LVT U482 ( .A1(n423), .A2(n264), .A3(n263), .Y(n267) );
  NAND2X0_LVT U483 ( .A1(n_T_101[60]), .A2(n441), .Y(n266) );
  NAND2X0_LVT U484 ( .A1(n434), .A2(io_adder_out[3]), .Y(n265) );
  NAND4X0_LVT U485 ( .A1(n268), .A2(n267), .A3(n266), .A4(n265), .Y(io_out[3])
         );
  NAND2X0_LVT U486 ( .A1(n_T_101[59]), .A2(n441), .Y(n274) );
  NAND3X0_LVT U487 ( .A1(io_in2[4]), .A2(n122), .A3(io_in1[4]), .Y(n269) );
  OA21X1_LVT U488 ( .A1(n423), .A2(n270), .A3(n269), .Y(n273) );
  NAND2X0_LVT U489 ( .A1(n_T_101[4]), .A2(n121), .Y(n272) );
  NAND2X0_LVT U490 ( .A1(io_adder_out[4]), .A2(n434), .Y(n271) );
  NAND4X0_LVT U491 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .Y(io_out[4])
         );
  NAND2X0_LVT U492 ( .A1(n_T_101[5]), .A2(n121), .Y(n280) );
  NAND3X0_LVT U493 ( .A1(io_in2[5]), .A2(n122), .A3(io_in1[5]), .Y(n275) );
  OA21X1_LVT U494 ( .A1(n423), .A2(n276), .A3(n275), .Y(n279) );
  NAND2X0_LVT U495 ( .A1(io_adder_out[5]), .A2(n434), .Y(n278) );
  NAND2X0_LVT U496 ( .A1(n_T_101[58]), .A2(n441), .Y(n277) );
  NAND4X0_LVT U497 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .Y(io_out[5])
         );
  NAND2X0_LVT U498 ( .A1(io_adder_out[6]), .A2(n434), .Y(n286) );
  NAND3X0_LVT U499 ( .A1(io_in2[6]), .A2(n122), .A3(io_in1[6]), .Y(n281) );
  OA21X1_LVT U500 ( .A1(n423), .A2(n282), .A3(n281), .Y(n285) );
  NAND2X0_LVT U501 ( .A1(n_T_101[57]), .A2(n441), .Y(n284) );
  NAND2X0_LVT U502 ( .A1(n_T_101[6]), .A2(n121), .Y(n283) );
  NAND4X0_LVT U503 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .Y(io_out[6])
         );
  NAND2X0_LVT U504 ( .A1(n_T_101[7]), .A2(n121), .Y(n292) );
  NAND2X0_LVT U505 ( .A1(io_adder_out[7]), .A2(n434), .Y(n291) );
  NAND3X0_LVT U506 ( .A1(io_in2[7]), .A2(n122), .A3(io_in1[7]), .Y(n287) );
  OA21X1_LVT U507 ( .A1(n423), .A2(n288), .A3(n287), .Y(n290) );
  NAND2X0_LVT U508 ( .A1(n_T_101[56]), .A2(n441), .Y(n289) );
  NAND4X0_LVT U509 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .Y(io_out[7])
         );
  NAND2X0_LVT U510 ( .A1(io_adder_out[8]), .A2(n434), .Y(n298) );
  NAND3X0_LVT U511 ( .A1(io_in2[8]), .A2(n122), .A3(io_in1[8]), .Y(n293) );
  OA21X1_LVT U512 ( .A1(n423), .A2(n294), .A3(n293), .Y(n297) );
  NAND2X0_LVT U513 ( .A1(n_T_101[55]), .A2(n441), .Y(n296) );
  NAND2X0_LVT U514 ( .A1(n_T_101[8]), .A2(n121), .Y(n295) );
  NAND4X0_LVT U515 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .Y(io_out[8])
         );
  NAND2X0_LVT U516 ( .A1(io_adder_out[9]), .A2(n434), .Y(n305) );
  NAND2X0_LVT U517 ( .A1(n_T_101[9]), .A2(n121), .Y(n304) );
  NAND2X0_LVT U518 ( .A1(io_in2[9]), .A2(n435), .Y(n301) );
  OA22X1_LVT U519 ( .A1(io_in2[9]), .A2(n423), .A3(n118), .A4(n299), .Y(n300)
         );
  MUX21X1_LVT U520 ( .A1(n301), .A2(n300), .S0(io_in1[9]), .Y(n303) );
  NAND2X0_LVT U521 ( .A1(n_T_101[54]), .A2(n441), .Y(n302) );
  NAND4X0_LVT U522 ( .A1(n305), .A2(n304), .A3(n303), .A4(n302), .Y(io_out[9])
         );
  NAND2X0_LVT U523 ( .A1(io_adder_out[10]), .A2(n434), .Y(n311) );
  NAND3X0_LVT U524 ( .A1(io_in2[10]), .A2(n122), .A3(io_in1[10]), .Y(n306) );
  OA21X1_LVT U525 ( .A1(n423), .A2(n307), .A3(n306), .Y(n310) );
  NAND2X0_LVT U526 ( .A1(n_T_101[53]), .A2(n441), .Y(n309) );
  NAND2X0_LVT U527 ( .A1(n_T_101[10]), .A2(n121), .Y(n308) );
  NAND4X0_LVT U528 ( .A1(n311), .A2(n310), .A3(n309), .A4(n308), .Y(io_out[10]) );
  NAND2X0_LVT U529 ( .A1(io_adder_out[11]), .A2(n434), .Y(n317) );
  NAND3X0_LVT U530 ( .A1(io_in2[11]), .A2(n122), .A3(io_in1[11]), .Y(n312) );
  OA21X1_LVT U531 ( .A1(n423), .A2(n313), .A3(n312), .Y(n316) );
  NAND2X0_LVT U532 ( .A1(n_T_101[11]), .A2(n121), .Y(n315) );
  NAND2X0_LVT U533 ( .A1(n_T_101[52]), .A2(n441), .Y(n314) );
  NAND4X0_LVT U534 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .Y(io_out[11]) );
  NAND2X0_LVT U535 ( .A1(io_adder_out[12]), .A2(n434), .Y(n323) );
  NAND3X0_LVT U536 ( .A1(io_in2[12]), .A2(n122), .A3(io_in1[12]), .Y(n318) );
  OA21X1_LVT U537 ( .A1(n423), .A2(n319), .A3(n318), .Y(n322) );
  NAND2X0_LVT U538 ( .A1(n_T_101[51]), .A2(n441), .Y(n321) );
  NAND2X0_LVT U539 ( .A1(n_T_101[12]), .A2(n121), .Y(n320) );
  NAND4X0_LVT U540 ( .A1(n323), .A2(n322), .A3(n321), .A4(n320), .Y(io_out[12]) );
  NAND2X0_LVT U541 ( .A1(io_adder_out[14]), .A2(n434), .Y(n330) );
  NAND3X0_LVT U542 ( .A1(io_in2[14]), .A2(n122), .A3(io_in1[14]), .Y(n325) );
  OA21X1_LVT U543 ( .A1(n423), .A2(n326), .A3(n325), .Y(n329) );
  NAND2X0_LVT U544 ( .A1(n_T_101[49]), .A2(n441), .Y(n328) );
  NAND2X0_LVT U545 ( .A1(n_T_101[14]), .A2(n121), .Y(n327) );
  NAND4X0_LVT U546 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .Y(io_out[14]) );
  NAND2X0_LVT U547 ( .A1(n_T_101[15]), .A2(n121), .Y(n335) );
  NAND2X0_LVT U548 ( .A1(n_T_101[48]), .A2(n441), .Y(n334) );
  OR2X1_LVT U549 ( .A1(n423), .A2(n331), .Y(n333) );
  NAND3X0_LVT U550 ( .A1(io_in2[15]), .A2(n122), .A3(io_in1[15]), .Y(n332) );
  NAND4X0_LVT U551 ( .A1(n335), .A2(n334), .A3(n333), .A4(n332), .Y(n336) );
  AO21X1_LVT U552 ( .A1(io_adder_out[15]), .A2(n434), .A3(n336), .Y(io_out[15]) );
  NAND2X0_LVT U553 ( .A1(io_adder_out[16]), .A2(n434), .Y(n342) );
  NAND3X0_LVT U554 ( .A1(io_in2[16]), .A2(n122), .A3(io_in1[16]), .Y(n337) );
  OA21X1_LVT U555 ( .A1(n423), .A2(n338), .A3(n337), .Y(n341) );
  NAND2X0_LVT U556 ( .A1(n_T_101[47]), .A2(n441), .Y(n340) );
  NAND2X0_LVT U557 ( .A1(n_T_101[16]), .A2(n121), .Y(n339) );
  NAND4X0_LVT U558 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .Y(io_out[16]) );
  NAND2X0_LVT U559 ( .A1(io_adder_out[17]), .A2(n434), .Y(n348) );
  NAND3X0_LVT U560 ( .A1(io_in2[17]), .A2(n122), .A3(io_in1[17]), .Y(n343) );
  OA21X1_LVT U561 ( .A1(n423), .A2(n344), .A3(n343), .Y(n347) );
  NAND2X0_LVT U562 ( .A1(n_T_101[17]), .A2(n121), .Y(n346) );
  NAND2X0_LVT U563 ( .A1(n_T_101[46]), .A2(n441), .Y(n345) );
  NAND4X0_LVT U564 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(io_out[17]) );
  NAND2X0_LVT U565 ( .A1(io_adder_out[18]), .A2(n434), .Y(n354) );
  NAND3X0_LVT U566 ( .A1(io_in2[18]), .A2(n122), .A3(io_in1[18]), .Y(n349) );
  OA21X1_LVT U567 ( .A1(n423), .A2(n350), .A3(n349), .Y(n353) );
  NAND2X0_LVT U568 ( .A1(n_T_101[45]), .A2(n441), .Y(n352) );
  NAND2X0_LVT U569 ( .A1(n_T_101[18]), .A2(n121), .Y(n351) );
  NAND4X0_LVT U570 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .Y(io_out[18]) );
  NAND2X0_LVT U571 ( .A1(io_adder_out[19]), .A2(n434), .Y(n360) );
  NAND3X0_LVT U572 ( .A1(io_in2[19]), .A2(n122), .A3(io_in1[19]), .Y(n355) );
  OA21X1_LVT U573 ( .A1(n423), .A2(n356), .A3(n355), .Y(n359) );
  NAND2X0_LVT U574 ( .A1(n_T_101[19]), .A2(n121), .Y(n358) );
  NAND2X0_LVT U575 ( .A1(n_T_101[44]), .A2(n441), .Y(n357) );
  NAND4X0_LVT U576 ( .A1(n360), .A2(n359), .A3(n358), .A4(n357), .Y(io_out[19]) );
  NAND2X0_LVT U577 ( .A1(io_adder_out[20]), .A2(n434), .Y(n366) );
  NAND3X0_LVT U578 ( .A1(io_in2[20]), .A2(n122), .A3(io_in1[20]), .Y(n361) );
  OA21X1_LVT U579 ( .A1(n423), .A2(n362), .A3(n361), .Y(n365) );
  NAND2X0_LVT U580 ( .A1(n_T_101[43]), .A2(n441), .Y(n364) );
  NAND2X0_LVT U581 ( .A1(n_T_101[20]), .A2(n121), .Y(n363) );
  NAND4X0_LVT U582 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .Y(io_out[20]) );
  NAND2X0_LVT U583 ( .A1(io_adder_out[21]), .A2(n434), .Y(n372) );
  NAND3X0_LVT U584 ( .A1(io_in2[21]), .A2(n122), .A3(io_in1[21]), .Y(n367) );
  OA21X1_LVT U585 ( .A1(n423), .A2(n368), .A3(n367), .Y(n371) );
  NAND2X0_LVT U586 ( .A1(n_T_101[21]), .A2(n121), .Y(n370) );
  NAND2X0_LVT U587 ( .A1(n_T_101[42]), .A2(n441), .Y(n369) );
  NAND4X0_LVT U588 ( .A1(n372), .A2(n371), .A3(n370), .A4(n369), .Y(io_out[21]) );
  NAND2X0_LVT U589 ( .A1(io_adder_out[22]), .A2(n434), .Y(n378) );
  NAND3X0_LVT U590 ( .A1(io_in2[22]), .A2(n122), .A3(io_in1[22]), .Y(n373) );
  OA21X1_LVT U591 ( .A1(n423), .A2(n374), .A3(n373), .Y(n377) );
  NAND2X0_LVT U592 ( .A1(n_T_101[41]), .A2(n441), .Y(n376) );
  NAND2X0_LVT U593 ( .A1(n_T_101[22]), .A2(n121), .Y(n375) );
  NAND4X0_LVT U594 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .Y(io_out[22]) );
  NAND2X0_LVT U595 ( .A1(io_adder_out[23]), .A2(n434), .Y(n384) );
  NAND3X0_LVT U596 ( .A1(io_in2[23]), .A2(n122), .A3(io_in1[23]), .Y(n379) );
  OA21X1_LVT U597 ( .A1(n423), .A2(n380), .A3(n379), .Y(n383) );
  NAND2X0_LVT U598 ( .A1(n_T_101[23]), .A2(n121), .Y(n382) );
  NAND2X0_LVT U599 ( .A1(n_T_101[40]), .A2(n441), .Y(n381) );
  NAND4X0_LVT U600 ( .A1(n384), .A2(n383), .A3(n382), .A4(n381), .Y(io_out[23]) );
  NAND2X0_LVT U601 ( .A1(io_adder_out[24]), .A2(n434), .Y(n390) );
  NAND3X0_LVT U602 ( .A1(io_in2[24]), .A2(n122), .A3(io_in1[24]), .Y(n385) );
  OA21X1_LVT U603 ( .A1(n423), .A2(n386), .A3(n385), .Y(n389) );
  NAND2X0_LVT U604 ( .A1(n_T_101[39]), .A2(n441), .Y(n388) );
  NAND2X0_LVT U605 ( .A1(n_T_101[24]), .A2(n121), .Y(n387) );
  NAND4X0_LVT U606 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .Y(io_out[24]) );
  NAND2X0_LVT U607 ( .A1(io_adder_out[25]), .A2(n434), .Y(n396) );
  NAND3X0_LVT U608 ( .A1(io_in2[25]), .A2(n122), .A3(io_in1[25]), .Y(n391) );
  OA21X1_LVT U609 ( .A1(n423), .A2(n392), .A3(n391), .Y(n395) );
  NAND2X0_LVT U610 ( .A1(n_T_101[25]), .A2(n121), .Y(n394) );
  NAND2X0_LVT U611 ( .A1(n_T_101[38]), .A2(n441), .Y(n393) );
  NAND4X0_LVT U612 ( .A1(n396), .A2(n395), .A3(n394), .A4(n393), .Y(io_out[25]) );
  NAND2X0_LVT U613 ( .A1(io_adder_out[26]), .A2(n434), .Y(n402) );
  NAND3X0_LVT U614 ( .A1(io_in2[26]), .A2(n122), .A3(io_in1[26]), .Y(n397) );
  OA21X1_LVT U615 ( .A1(n423), .A2(n398), .A3(n397), .Y(n401) );
  NAND2X0_LVT U616 ( .A1(n_T_101[37]), .A2(n441), .Y(n400) );
  NAND2X0_LVT U617 ( .A1(n_T_101[26]), .A2(n121), .Y(n399) );
  NAND4X0_LVT U618 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .Y(io_out[26]) );
  NAND2X0_LVT U619 ( .A1(io_adder_out[27]), .A2(n434), .Y(n408) );
  NAND3X0_LVT U620 ( .A1(io_in2[27]), .A2(n122), .A3(io_in1[27]), .Y(n403) );
  OA21X1_LVT U621 ( .A1(n423), .A2(n404), .A3(n403), .Y(n407) );
  NAND2X0_LVT U622 ( .A1(n_T_101[27]), .A2(n121), .Y(n406) );
  NAND2X0_LVT U623 ( .A1(n_T_101[36]), .A2(n441), .Y(n405) );
  NAND4X0_LVT U624 ( .A1(n408), .A2(n407), .A3(n406), .A4(n405), .Y(io_out[27]) );
  NAND2X0_LVT U625 ( .A1(io_adder_out[28]), .A2(n434), .Y(n414) );
  NAND3X0_LVT U626 ( .A1(io_in2[28]), .A2(n122), .A3(io_in1[28]), .Y(n409) );
  OA21X1_LVT U627 ( .A1(n423), .A2(n410), .A3(n409), .Y(n413) );
  NAND2X0_LVT U628 ( .A1(n_T_101[35]), .A2(n441), .Y(n412) );
  NAND2X0_LVT U629 ( .A1(n_T_101[28]), .A2(n121), .Y(n411) );
  NAND4X0_LVT U630 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .Y(io_out[28]) );
  NAND2X0_LVT U631 ( .A1(io_adder_out[29]), .A2(n434), .Y(n420) );
  NAND3X0_LVT U632 ( .A1(io_in2[29]), .A2(n122), .A3(io_in1[29]), .Y(n415) );
  OA21X1_LVT U633 ( .A1(n423), .A2(n416), .A3(n415), .Y(n419) );
  NAND2X0_LVT U634 ( .A1(n_T_101[29]), .A2(n121), .Y(n418) );
  NAND2X0_LVT U635 ( .A1(n_T_101[34]), .A2(n441), .Y(n417) );
  NAND4X0_LVT U636 ( .A1(n420), .A2(n419), .A3(n418), .A4(n417), .Y(io_out[29]) );
  NAND2X0_LVT U637 ( .A1(io_adder_out[30]), .A2(n434), .Y(n427) );
  NAND3X0_LVT U638 ( .A1(io_in2[30]), .A2(n122), .A3(io_in1[30]), .Y(n421) );
  OA21X1_LVT U639 ( .A1(n423), .A2(n422), .A3(n421), .Y(n426) );
  NAND2X0_LVT U640 ( .A1(n_T_101[33]), .A2(n441), .Y(n425) );
  NAND2X0_LVT U641 ( .A1(n_T_101[30]), .A2(n121), .Y(n424) );
  NAND4X0_LVT U642 ( .A1(n427), .A2(n426), .A3(n425), .A4(n424), .Y(io_out[30]) );
  NAND2X0_LVT U643 ( .A1(n_T_101[31]), .A2(n121), .Y(n432) );
  NAND2X0_LVT U644 ( .A1(n_T_101[32]), .A2(n441), .Y(n431) );
  NAND2X0_LVT U645 ( .A1(n428), .A2(n435), .Y(n430) );
  NAND3X0_LVT U646 ( .A1(io_in2[31]), .A2(n122), .A3(io_in1[31]), .Y(n429) );
  NAND4X0_LVT U647 ( .A1(n432), .A2(n431), .A3(n430), .A4(n429), .Y(n433) );
  AO21X1_LVT U648 ( .A1(n434), .A2(io_adder_out[31]), .A3(n433), .Y(io_out[31]) );
  NAND2X0_LVT U649 ( .A1(io_adder_out[32]), .A2(n602), .Y(n444) );
  AND2X1_LVT U650 ( .A1(n435), .A2(io_dw), .Y(n593) );
  NAND3X0_LVT U651 ( .A1(io_in2[32]), .A2(n603), .A3(io_in1[32]), .Y(n436) );
  OA21X1_LVT U652 ( .A1(n605), .A2(n437), .A3(n436), .Y(n438) );
  OA21X1_LVT U653 ( .A1(n117), .A2(n439), .A3(n438), .Y(n443) );
  NAND2X0_LVT U654 ( .A1(io_out[31]), .A2(n440), .Y(n606) );
  NAND2X0_LVT U655 ( .A1(n_T_101[31]), .A2(n598), .Y(n442) );
  NAND4X0_LVT U656 ( .A1(n444), .A2(n443), .A3(n115), .A4(n442), .Y(io_out[32]) );
  NAND2X0_LVT U657 ( .A1(io_adder_out[33]), .A2(n602), .Y(n451) );
  NAND3X0_LVT U658 ( .A1(io_in2[33]), .A2(n603), .A3(io_in1[33]), .Y(n445) );
  OA21X1_LVT U659 ( .A1(n605), .A2(n446), .A3(n445), .Y(n447) );
  OA21X1_LVT U660 ( .A1(n123), .A2(n448), .A3(n447), .Y(n450) );
  NAND2X0_LVT U661 ( .A1(n_T_101[33]), .A2(n124), .Y(n449) );
  NAND4X0_LVT U662 ( .A1(n115), .A2(n451), .A3(n450), .A4(n449), .Y(io_out[33]) );
  NAND3X0_LVT U663 ( .A1(io_in2[40]), .A2(n603), .A3(io_in1[40]), .Y(n458) );
  OA21X1_LVT U664 ( .A1(n605), .A2(n459), .A3(n458), .Y(n462) );
  NAND2X0_LVT U665 ( .A1(n_T_101[23]), .A2(n598), .Y(n461) );
  NAND2X0_LVT U666 ( .A1(n_T_101[40]), .A2(n124), .Y(n460) );
  NAND4X0_LVT U667 ( .A1(n606), .A2(n462), .A3(n461), .A4(n460), .Y(n463) );
  AO21X1_LVT U668 ( .A1(n602), .A2(n630), .A3(n463), .Y(io_out[40]) );
  NAND3X0_LVT U669 ( .A1(io_in2[41]), .A2(n603), .A3(io_in1[41]), .Y(n464) );
  OA21X1_LVT U670 ( .A1(n605), .A2(n465), .A3(n464), .Y(n468) );
  NAND2X0_LVT U671 ( .A1(n_T_101[41]), .A2(n124), .Y(n467) );
  NAND2X0_LVT U672 ( .A1(n_T_101[22]), .A2(n598), .Y(n466) );
  NAND4X0_LVT U673 ( .A1(n115), .A2(n468), .A3(n467), .A4(n466), .Y(n469) );
  AO21X1_LVT U674 ( .A1(n602), .A2(n629), .A3(n469), .Y(io_out[41]) );
  NAND3X0_LVT U675 ( .A1(io_in2[42]), .A2(n603), .A3(io_in1[42]), .Y(n470) );
  OA21X1_LVT U676 ( .A1(n605), .A2(n471), .A3(n470), .Y(n474) );
  NAND2X0_LVT U677 ( .A1(n_T_101[21]), .A2(n598), .Y(n473) );
  NAND2X0_LVT U678 ( .A1(n_T_101[42]), .A2(n124), .Y(n472) );
  NAND4X0_LVT U679 ( .A1(n115), .A2(n474), .A3(n473), .A4(n472), .Y(n475) );
  AO21X1_LVT U680 ( .A1(n602), .A2(n628), .A3(n475), .Y(io_out[42]) );
  NAND3X0_LVT U681 ( .A1(io_in2[43]), .A2(n603), .A3(io_in1[43]), .Y(n476) );
  OA21X1_LVT U682 ( .A1(n605), .A2(n477), .A3(n476), .Y(n480) );
  NAND2X0_LVT U683 ( .A1(n_T_101[43]), .A2(n124), .Y(n479) );
  NAND2X0_LVT U684 ( .A1(n_T_101[20]), .A2(n598), .Y(n478) );
  NAND4X0_LVT U685 ( .A1(n115), .A2(n480), .A3(n479), .A4(n478), .Y(n481) );
  AO21X1_LVT U686 ( .A1(n602), .A2(n627), .A3(n481), .Y(io_out[43]) );
  NAND3X0_LVT U687 ( .A1(io_in2[44]), .A2(n603), .A3(io_in1[44]), .Y(n482) );
  OA21X1_LVT U688 ( .A1(n605), .A2(n483), .A3(n482), .Y(n486) );
  NAND2X0_LVT U689 ( .A1(n_T_101[19]), .A2(n598), .Y(n485) );
  NAND2X0_LVT U690 ( .A1(n_T_101[44]), .A2(n124), .Y(n484) );
  NAND4X0_LVT U691 ( .A1(n115), .A2(n486), .A3(n485), .A4(n484), .Y(n487) );
  AO21X1_LVT U692 ( .A1(n602), .A2(n626), .A3(n487), .Y(io_out[44]) );
  NAND3X0_LVT U693 ( .A1(io_in2[45]), .A2(n603), .A3(io_in1[45]), .Y(n488) );
  OA21X1_LVT U694 ( .A1(n605), .A2(n489), .A3(n488), .Y(n492) );
  NAND2X0_LVT U695 ( .A1(n_T_101[45]), .A2(n124), .Y(n491) );
  NAND2X0_LVT U696 ( .A1(n_T_101[18]), .A2(n598), .Y(n490) );
  NAND4X0_LVT U697 ( .A1(n606), .A2(n492), .A3(n491), .A4(n490), .Y(n493) );
  AO21X1_LVT U698 ( .A1(n602), .A2(n625), .A3(n493), .Y(io_out[45]) );
  NAND3X0_LVT U699 ( .A1(io_in2[46]), .A2(n603), .A3(io_in1[46]), .Y(n494) );
  OA21X1_LVT U700 ( .A1(n605), .A2(n495), .A3(n494), .Y(n498) );
  NAND2X0_LVT U701 ( .A1(n_T_101[17]), .A2(n598), .Y(n497) );
  NAND2X0_LVT U702 ( .A1(n_T_101[46]), .A2(n124), .Y(n496) );
  NAND4X0_LVT U703 ( .A1(n606), .A2(n498), .A3(n497), .A4(n496), .Y(n499) );
  AO21X1_LVT U704 ( .A1(n602), .A2(n624), .A3(n499), .Y(io_out[46]) );
  NAND2X0_LVT U705 ( .A1(n623), .A2(n602), .Y(n506) );
  NAND3X0_LVT U706 ( .A1(io_in2[47]), .A2(n603), .A3(io_in1[47]), .Y(n500) );
  OA21X1_LVT U707 ( .A1(n605), .A2(n501), .A3(n500), .Y(n502) );
  OA21X1_LVT U708 ( .A1(n123), .A2(n503), .A3(n502), .Y(n505) );
  NAND2X0_LVT U709 ( .A1(n_T_101[47]), .A2(n124), .Y(n504) );
  NAND4X0_LVT U710 ( .A1(n606), .A2(n506), .A3(n505), .A4(n504), .Y(io_out[47]) );
  NAND3X0_LVT U711 ( .A1(io_in2[48]), .A2(n603), .A3(io_in1[48]), .Y(n507) );
  OA21X1_LVT U712 ( .A1(n605), .A2(n508), .A3(n507), .Y(n511) );
  NAND2X0_LVT U713 ( .A1(n_T_101[15]), .A2(n598), .Y(n510) );
  NAND2X0_LVT U714 ( .A1(n_T_101[48]), .A2(n124), .Y(n509) );
  NAND4X0_LVT U715 ( .A1(n606), .A2(n511), .A3(n510), .A4(n509), .Y(n512) );
  AO21X1_LVT U716 ( .A1(n602), .A2(n622), .A3(n512), .Y(io_out[48]) );
  NAND3X0_LVT U717 ( .A1(io_in2[49]), .A2(n603), .A3(io_in1[49]), .Y(n513) );
  OA21X1_LVT U718 ( .A1(n605), .A2(n514), .A3(n513), .Y(n517) );
  NAND2X0_LVT U719 ( .A1(n_T_101[49]), .A2(n124), .Y(n516) );
  NAND2X0_LVT U720 ( .A1(n_T_101[14]), .A2(n598), .Y(n515) );
  NAND4X0_LVT U721 ( .A1(n606), .A2(n517), .A3(n516), .A4(n515), .Y(n518) );
  AO21X1_LVT U722 ( .A1(n602), .A2(n621), .A3(n518), .Y(io_out[49]) );
  NAND3X0_LVT U723 ( .A1(io_in2[50]), .A2(n603), .A3(io_in1[50]), .Y(n519) );
  OA21X1_LVT U724 ( .A1(n605), .A2(n520), .A3(n519), .Y(n523) );
  NAND2X0_LVT U725 ( .A1(n_T_101[13]), .A2(n598), .Y(n522) );
  NAND2X0_LVT U726 ( .A1(n_T_101[50]), .A2(n124), .Y(n521) );
  NAND4X0_LVT U727 ( .A1(n606), .A2(n523), .A3(n522), .A4(n521), .Y(n524) );
  AO21X1_LVT U728 ( .A1(n602), .A2(n620), .A3(n524), .Y(io_out[50]) );
  NAND3X0_LVT U729 ( .A1(io_in2[51]), .A2(n603), .A3(io_in1[51]), .Y(n525) );
  OA21X1_LVT U730 ( .A1(n605), .A2(n526), .A3(n525), .Y(n529) );
  NAND2X0_LVT U731 ( .A1(n_T_101[51]), .A2(n124), .Y(n528) );
  NAND2X0_LVT U732 ( .A1(n_T_101[12]), .A2(n598), .Y(n527) );
  NAND4X0_LVT U733 ( .A1(n606), .A2(n529), .A3(n528), .A4(n527), .Y(n530) );
  AO21X1_LVT U734 ( .A1(n602), .A2(n619), .A3(n530), .Y(io_out[51]) );
  NAND3X0_LVT U735 ( .A1(io_in2[52]), .A2(n603), .A3(io_in1[52]), .Y(n531) );
  OA21X1_LVT U736 ( .A1(n605), .A2(n532), .A3(n531), .Y(n535) );
  NAND2X0_LVT U737 ( .A1(n_T_101[11]), .A2(n598), .Y(n534) );
  NAND2X0_LVT U738 ( .A1(n_T_101[52]), .A2(n124), .Y(n533) );
  NAND4X0_LVT U739 ( .A1(n606), .A2(n535), .A3(n534), .A4(n533), .Y(n536) );
  AO21X1_LVT U740 ( .A1(n602), .A2(n618), .A3(n536), .Y(io_out[52]) );
  NAND3X0_LVT U741 ( .A1(io_in2[53]), .A2(n603), .A3(io_in1[53]), .Y(n537) );
  OA21X1_LVT U742 ( .A1(n605), .A2(n538), .A3(n537), .Y(n541) );
  NAND2X0_LVT U743 ( .A1(n_T_101[53]), .A2(n124), .Y(n540) );
  NAND2X0_LVT U744 ( .A1(n_T_101[10]), .A2(n598), .Y(n539) );
  NAND4X0_LVT U745 ( .A1(n606), .A2(n541), .A3(n540), .A4(n539), .Y(n542) );
  AO21X1_LVT U746 ( .A1(n602), .A2(n617), .A3(n542), .Y(io_out[53]) );
  NAND3X0_LVT U747 ( .A1(io_in2[54]), .A2(n603), .A3(io_in1[54]), .Y(n543) );
  OA21X1_LVT U748 ( .A1(n605), .A2(n544), .A3(n543), .Y(n547) );
  NAND2X0_LVT U749 ( .A1(n_T_101[9]), .A2(n598), .Y(n546) );
  NAND2X0_LVT U750 ( .A1(n_T_101[54]), .A2(n124), .Y(n545) );
  NAND4X0_LVT U751 ( .A1(n606), .A2(n547), .A3(n546), .A4(n545), .Y(n548) );
  AO21X1_LVT U752 ( .A1(n602), .A2(n616), .A3(n548), .Y(io_out[54]) );
  NAND3X0_LVT U753 ( .A1(io_in2[55]), .A2(n603), .A3(io_in1[55]), .Y(n549) );
  OA21X1_LVT U754 ( .A1(n605), .A2(n550), .A3(n549), .Y(n553) );
  NAND2X0_LVT U755 ( .A1(n_T_101[55]), .A2(n124), .Y(n552) );
  NAND2X0_LVT U756 ( .A1(n_T_101[8]), .A2(n598), .Y(n551) );
  NAND4X0_LVT U757 ( .A1(n606), .A2(n553), .A3(n552), .A4(n551), .Y(n554) );
  AO21X1_LVT U758 ( .A1(n602), .A2(n615), .A3(n554), .Y(io_out[55]) );
  NAND3X0_LVT U759 ( .A1(io_in2[56]), .A2(n603), .A3(io_in1[56]), .Y(n555) );
  OA21X1_LVT U760 ( .A1(n605), .A2(n556), .A3(n555), .Y(n559) );
  NAND2X0_LVT U761 ( .A1(n_T_101[7]), .A2(n598), .Y(n558) );
  NAND2X0_LVT U762 ( .A1(n_T_101[56]), .A2(n124), .Y(n557) );
  NAND4X0_LVT U763 ( .A1(n115), .A2(n559), .A3(n558), .A4(n557), .Y(n560) );
  AO21X1_LVT U764 ( .A1(n602), .A2(n614), .A3(n560), .Y(io_out[56]) );
  NAND3X0_LVT U765 ( .A1(io_in2[57]), .A2(n603), .A3(io_in1[57]), .Y(n561) );
  OA21X1_LVT U766 ( .A1(n605), .A2(n562), .A3(n561), .Y(n565) );
  NAND2X0_LVT U767 ( .A1(n_T_101[57]), .A2(n124), .Y(n564) );
  NAND2X0_LVT U768 ( .A1(n_T_101[6]), .A2(n598), .Y(n563) );
  NAND4X0_LVT U769 ( .A1(n115), .A2(n565), .A3(n564), .A4(n563), .Y(n566) );
  AO21X1_LVT U770 ( .A1(n602), .A2(n613), .A3(n566), .Y(io_out[57]) );
  NAND3X0_LVT U771 ( .A1(io_in2[58]), .A2(n603), .A3(io_in1[58]), .Y(n567) );
  OA21X1_LVT U772 ( .A1(n605), .A2(n568), .A3(n567), .Y(n571) );
  NAND2X0_LVT U773 ( .A1(n_T_101[5]), .A2(n598), .Y(n570) );
  NAND2X0_LVT U774 ( .A1(n_T_101[58]), .A2(n124), .Y(n569) );
  NAND4X0_LVT U775 ( .A1(n115), .A2(n571), .A3(n570), .A4(n569), .Y(n572) );
  AO21X1_LVT U776 ( .A1(n602), .A2(n612), .A3(n572), .Y(io_out[58]) );
  NAND2X0_LVT U777 ( .A1(n611), .A2(n602), .Y(n579) );
  NAND2X0_LVT U778 ( .A1(n_T_101[59]), .A2(n124), .Y(n577) );
  NAND2X0_LVT U779 ( .A1(n_T_101[4]), .A2(n598), .Y(n576) );
  NAND2X0_LVT U780 ( .A1(n573), .A2(n593), .Y(n575) );
  NAND3X0_LVT U781 ( .A1(io_in2[59]), .A2(n603), .A3(io_in1[59]), .Y(n574) );
  AND4X1_LVT U782 ( .A1(n577), .A2(n576), .A3(n575), .A4(n574), .Y(n578) );
  NAND3X0_LVT U783 ( .A1(n579), .A2(n578), .A3(n115), .Y(io_out[59]) );
  NAND2X0_LVT U784 ( .A1(n610), .A2(n602), .Y(n586) );
  NAND2X0_LVT U785 ( .A1(n_T_101[3]), .A2(n598), .Y(n584) );
  NAND2X0_LVT U786 ( .A1(n_T_101[60]), .A2(n124), .Y(n583) );
  NAND2X0_LVT U787 ( .A1(n580), .A2(n593), .Y(n582) );
  NAND3X0_LVT U788 ( .A1(io_in2[60]), .A2(n603), .A3(io_in1[60]), .Y(n581) );
  AND4X1_LVT U789 ( .A1(n584), .A2(n583), .A3(n582), .A4(n581), .Y(n585) );
  NAND3X0_LVT U790 ( .A1(n586), .A2(n585), .A3(n115), .Y(io_out[60]) );
  NAND3X0_LVT U791 ( .A1(io_in2[61]), .A2(n603), .A3(io_in1[61]), .Y(n587) );
  OA21X1_LVT U792 ( .A1(n605), .A2(n588), .A3(n587), .Y(n591) );
  NAND2X0_LVT U793 ( .A1(n_T_101[61]), .A2(n124), .Y(n590) );
  NAND2X0_LVT U794 ( .A1(n_T_101[2]), .A2(n598), .Y(n589) );
  NAND4X0_LVT U795 ( .A1(n115), .A2(n591), .A3(n590), .A4(n589), .Y(n592) );
  AO21X1_LVT U796 ( .A1(n602), .A2(n609), .A3(n592), .Y(io_out[61]) );
  NAND2X0_LVT U797 ( .A1(n_T_101[62]), .A2(n124), .Y(n597) );
  NAND2X0_LVT U798 ( .A1(n594), .A2(n593), .Y(n596) );
  NAND3X0_LVT U799 ( .A1(io_in2[62]), .A2(n603), .A3(io_in1[62]), .Y(n595) );
  AND3X1_LVT U800 ( .A1(n597), .A2(n596), .A3(n595), .Y(n600) );
  NAND2X0_LVT U801 ( .A1(n_T_101[1]), .A2(n598), .Y(n599) );
  NAND3X0_LVT U802 ( .A1(n115), .A2(n600), .A3(n599), .Y(n601) );
  AO21X1_LVT U803 ( .A1(n602), .A2(n608), .A3(n601), .Y(io_out[62]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_MulDiv_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module MulDiv_DP_OP_279J39_124_314_J39_0 ( I1, I2, I3, O1 );
  input [8:0] I1;
  input [64:0] I2;
  input [64:0] I3;
  output [72:0] O1;
  wire   n551, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2527, n2528, n2529, n2530, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787;

  FADDX1_LVT U692 ( .A(n2171), .B(n2586), .CI(n1650), .CO(n551), .S(O1[1]) );
  FADDX1_LVT U699 ( .A(n1717), .B(n1653), .CI(n631), .CO(n627), .S(n628) );
  FADDX1_LVT U700 ( .A(n637), .B(n632), .CI(n635), .CO(n629), .S(n630) );
  FADDX1_LVT U701 ( .A(n1782), .B(n1654), .CI(n1718), .CO(n631), .S(n632) );
  FADDX1_LVT U702 ( .A(n643), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  FADDX1_LVT U703 ( .A(n1719), .B(n645), .CI(n638), .CO(n635), .S(n636) );
  FADDX1_LVT U704 ( .A(n1847), .B(n1655), .CI(n1783), .CO(n637), .S(n638) );
  FADDX1_LVT U705 ( .A(n651), .B(n649), .CI(n642), .CO(n639), .S(n640) );
  FADDX1_LVT U706 ( .A(n653), .B(n646), .CI(n644), .CO(n641), .S(n642) );
  FADDX1_LVT U707 ( .A(n1784), .B(n1720), .CI(n655), .CO(n643), .S(n644) );
  FADDX1_LVT U708 ( .A(n1912), .B(n1656), .CI(n1848), .CO(n645), .S(n646) );
  FADDX1_LVT U709 ( .A(n652), .B(n659), .CI(n650), .CO(n647), .S(n648) );
  FADDX1_LVT U710 ( .A(n654), .B(n663), .CI(n661), .CO(n649), .S(n650) );
  FADDX1_LVT U711 ( .A(n667), .B(n665), .CI(n656), .CO(n651), .S(n652) );
  FADDX1_LVT U712 ( .A(n1721), .B(n1785), .CI(n1849), .CO(n653), .S(n654) );
  FADDX1_LVT U713 ( .A(n1977), .B(n1657), .CI(n1913), .CO(n655), .S(n656) );
  FADDX1_LVT U714 ( .A(n662), .B(n671), .CI(n660), .CO(n657), .S(n658) );
  FADDX1_LVT U715 ( .A(n675), .B(n664), .CI(n673), .CO(n659), .S(n660) );
  FADDX1_LVT U716 ( .A(n668), .B(n666), .CI(n677), .CO(n661), .S(n662) );
  FADDX1_LVT U717 ( .A(n1786), .B(n681), .CI(n679), .CO(n663), .S(n664) );
  FADDX1_LVT U718 ( .A(n1722), .B(n1914), .CI(n1850), .CO(n665), .S(n666) );
  FADDX1_LVT U719 ( .A(n2042), .B(n1658), .CI(n1978), .CO(n667), .S(n668) );
  FADDX1_LVT U720 ( .A(n674), .B(n685), .CI(n672), .CO(n669), .S(n670) );
  FADDX1_LVT U721 ( .A(n689), .B(n676), .CI(n687), .CO(n671), .S(n672) );
  FADDX1_LVT U722 ( .A(n680), .B(n691), .CI(n678), .CO(n673), .S(n674) );
  FADDX1_LVT U723 ( .A(n695), .B(n693), .CI(n682), .CO(n675), .S(n676) );
  FADDX1_LVT U724 ( .A(n1915), .B(n1851), .CI(n697), .CO(n677), .S(n678) );
  FADDX1_LVT U725 ( .A(n1979), .B(n1723), .CI(n1787), .CO(n679), .S(n680) );
  FADDX1_LVT U726 ( .A(n2107), .B(n1659), .CI(n2043), .CO(n681), .S(n682) );
  FADDX1_LVT U727 ( .A(n688), .B(n701), .CI(n686), .CO(n683), .S(n684) );
  FADDX1_LVT U728 ( .A(n692), .B(n690), .CI(n703), .CO(n685), .S(n686) );
  FADDX1_LVT U729 ( .A(n696), .B(n707), .CI(n705), .CO(n687), .S(n688) );
  FADDX1_LVT U730 ( .A(n709), .B(n698), .CI(n694), .CO(n689), .S(n690) );
  FADDX1_LVT U731 ( .A(n1980), .B(n713), .CI(n711), .CO(n691), .S(n692) );
  FADDX1_LVT U732 ( .A(n2044), .B(n1852), .CI(n1916), .CO(n693), .S(n694) );
  FADDX1_LVT U733 ( .A(n2108), .B(n1724), .CI(n1788), .CO(n695), .S(n696) );
  FADDX1_LVT U734 ( .A(n2587), .B(n1660), .CI(n2172), .CO(n697), .S(n698) );
  FADDX1_LVT U735 ( .A(n704), .B(n717), .CI(n702), .CO(n699), .S(n700) );
  FADDX1_LVT U736 ( .A(n708), .B(n706), .CI(n719), .CO(n701), .S(n702) );
  FADDX1_LVT U737 ( .A(n712), .B(n723), .CI(n721), .CO(n703), .S(n704) );
  FADDX1_LVT U738 ( .A(n725), .B(n714), .CI(n710), .CO(n705), .S(n706) );
  FADDX1_LVT U739 ( .A(n1981), .B(n729), .CI(n727), .CO(n707), .S(n708) );
  FADDX1_LVT U740 ( .A(n2045), .B(n1853), .CI(n1917), .CO(n709), .S(n710) );
  FADDX1_LVT U741 ( .A(n2109), .B(n1725), .CI(n1789), .CO(n711), .S(n712) );
  FADDX1_LVT U742 ( .A(I3[63]), .B(n1661), .CI(n2173), .CO(n713), .S(n714) );
  FADDX1_LVT U743 ( .A(n720), .B(n733), .CI(n718), .CO(n715), .S(n716) );
  FADDX1_LVT U744 ( .A(n724), .B(n722), .CI(n735), .CO(n717), .S(n718) );
  FADDX1_LVT U745 ( .A(n728), .B(n739), .CI(n737), .CO(n719), .S(n720) );
  FADDX1_LVT U746 ( .A(n741), .B(n730), .CI(n726), .CO(n721), .S(n722) );
  FADDX1_LVT U747 ( .A(n1982), .B(n745), .CI(n743), .CO(n723), .S(n724) );
  FADDX1_LVT U748 ( .A(n2046), .B(n1854), .CI(n1918), .CO(n725), .S(n726) );
  FADDX1_LVT U749 ( .A(n2110), .B(n1726), .CI(n1790), .CO(n727), .S(n728) );
  FADDX1_LVT U750 ( .A(I3[62]), .B(n1662), .CI(n2174), .CO(n729), .S(n730) );
  FADDX1_LVT U751 ( .A(n736), .B(n749), .CI(n734), .CO(n731), .S(n732) );
  FADDX1_LVT U752 ( .A(n740), .B(n738), .CI(n751), .CO(n733), .S(n734) );
  FADDX1_LVT U753 ( .A(n744), .B(n755), .CI(n753), .CO(n735), .S(n736) );
  FADDX1_LVT U754 ( .A(n757), .B(n746), .CI(n742), .CO(n737), .S(n738) );
  FADDX1_LVT U755 ( .A(n1983), .B(n761), .CI(n759), .CO(n739), .S(n740) );
  FADDX1_LVT U756 ( .A(n2047), .B(n1855), .CI(n1919), .CO(n741), .S(n742) );
  FADDX1_LVT U757 ( .A(n2111), .B(n1727), .CI(n1791), .CO(n743), .S(n744) );
  FADDX1_LVT U758 ( .A(I3[61]), .B(n1663), .CI(n2175), .CO(n745), .S(n746) );
  FADDX1_LVT U759 ( .A(n752), .B(n765), .CI(n750), .CO(n747), .S(n748) );
  FADDX1_LVT U760 ( .A(n756), .B(n754), .CI(n767), .CO(n749), .S(n750) );
  FADDX1_LVT U761 ( .A(n760), .B(n771), .CI(n769), .CO(n751), .S(n752) );
  FADDX1_LVT U762 ( .A(n773), .B(n762), .CI(n758), .CO(n753), .S(n754) );
  FADDX1_LVT U763 ( .A(n1984), .B(n777), .CI(n775), .CO(n755), .S(n756) );
  FADDX1_LVT U764 ( .A(n2048), .B(n1856), .CI(n1920), .CO(n757), .S(n758) );
  FADDX1_LVT U765 ( .A(n2112), .B(n1728), .CI(n1792), .CO(n759), .S(n760) );
  FADDX1_LVT U766 ( .A(I3[60]), .B(n1664), .CI(n2176), .CO(n761), .S(n762) );
  FADDX1_LVT U767 ( .A(n768), .B(n781), .CI(n766), .CO(n763), .S(n764) );
  FADDX1_LVT U768 ( .A(n772), .B(n770), .CI(n783), .CO(n765), .S(n766) );
  FADDX1_LVT U769 ( .A(n776), .B(n787), .CI(n785), .CO(n767), .S(n768) );
  FADDX1_LVT U770 ( .A(n789), .B(n778), .CI(n774), .CO(n769), .S(n770) );
  FADDX1_LVT U771 ( .A(n1985), .B(n793), .CI(n791), .CO(n771), .S(n772) );
  FADDX1_LVT U772 ( .A(n2049), .B(n1857), .CI(n1921), .CO(n773), .S(n774) );
  FADDX1_LVT U773 ( .A(n2113), .B(n1729), .CI(n1793), .CO(n775), .S(n776) );
  FADDX1_LVT U774 ( .A(I3[59]), .B(n1665), .CI(n2177), .CO(n777), .S(n778) );
  FADDX1_LVT U775 ( .A(n784), .B(n797), .CI(n782), .CO(n779), .S(n780) );
  FADDX1_LVT U776 ( .A(n788), .B(n786), .CI(n799), .CO(n781), .S(n782) );
  FADDX1_LVT U777 ( .A(n792), .B(n803), .CI(n801), .CO(n783), .S(n784) );
  FADDX1_LVT U778 ( .A(n805), .B(n794), .CI(n790), .CO(n785), .S(n786) );
  FADDX1_LVT U779 ( .A(n1986), .B(n809), .CI(n807), .CO(n787), .S(n788) );
  FADDX1_LVT U780 ( .A(n2050), .B(n1858), .CI(n1922), .CO(n789), .S(n790) );
  FADDX1_LVT U781 ( .A(n2114), .B(n1730), .CI(n1794), .CO(n791), .S(n792) );
  FADDX1_LVT U782 ( .A(I3[58]), .B(n1666), .CI(n2178), .CO(n793), .S(n794) );
  FADDX1_LVT U783 ( .A(n800), .B(n813), .CI(n798), .CO(n795), .S(n796) );
  FADDX1_LVT U784 ( .A(n804), .B(n802), .CI(n815), .CO(n797), .S(n798) );
  FADDX1_LVT U785 ( .A(n808), .B(n819), .CI(n817), .CO(n799), .S(n800) );
  FADDX1_LVT U786 ( .A(n821), .B(n810), .CI(n806), .CO(n801), .S(n802) );
  FADDX1_LVT U787 ( .A(n1987), .B(n825), .CI(n823), .CO(n803), .S(n804) );
  FADDX1_LVT U788 ( .A(n2051), .B(n1859), .CI(n1923), .CO(n805), .S(n806) );
  FADDX1_LVT U789 ( .A(n2115), .B(n1731), .CI(n1795), .CO(n807), .S(n808) );
  FADDX1_LVT U790 ( .A(I3[57]), .B(n1667), .CI(n2179), .CO(n809), .S(n810) );
  FADDX1_LVT U791 ( .A(n816), .B(n829), .CI(n814), .CO(n811), .S(n812) );
  FADDX1_LVT U792 ( .A(n820), .B(n818), .CI(n831), .CO(n813), .S(n814) );
  FADDX1_LVT U793 ( .A(n824), .B(n835), .CI(n833), .CO(n815), .S(n816) );
  FADDX1_LVT U794 ( .A(n837), .B(n826), .CI(n822), .CO(n817), .S(n818) );
  FADDX1_LVT U795 ( .A(n1988), .B(n841), .CI(n839), .CO(n819), .S(n820) );
  FADDX1_LVT U796 ( .A(n2052), .B(n1860), .CI(n1924), .CO(n821), .S(n822) );
  FADDX1_LVT U797 ( .A(n2116), .B(n1732), .CI(n1796), .CO(n823), .S(n824) );
  FADDX1_LVT U798 ( .A(I3[56]), .B(n1668), .CI(n2180), .CO(n825), .S(n826) );
  FADDX1_LVT U799 ( .A(n832), .B(n845), .CI(n830), .CO(n827), .S(n828) );
  FADDX1_LVT U800 ( .A(n836), .B(n834), .CI(n847), .CO(n829), .S(n830) );
  FADDX1_LVT U801 ( .A(n840), .B(n851), .CI(n849), .CO(n831), .S(n832) );
  FADDX1_LVT U802 ( .A(n853), .B(n842), .CI(n838), .CO(n833), .S(n834) );
  FADDX1_LVT U803 ( .A(n1989), .B(n857), .CI(n855), .CO(n835), .S(n836) );
  FADDX1_LVT U804 ( .A(n2053), .B(n1861), .CI(n1925), .CO(n837), .S(n838) );
  FADDX1_LVT U805 ( .A(n2117), .B(n1733), .CI(n1797), .CO(n839), .S(n840) );
  FADDX1_LVT U806 ( .A(I3[55]), .B(n1669), .CI(n2181), .CO(n841), .S(n842) );
  FADDX1_LVT U807 ( .A(n848), .B(n861), .CI(n846), .CO(n843), .S(n844) );
  FADDX1_LVT U808 ( .A(n852), .B(n850), .CI(n863), .CO(n845), .S(n846) );
  FADDX1_LVT U809 ( .A(n856), .B(n867), .CI(n865), .CO(n847), .S(n848) );
  FADDX1_LVT U810 ( .A(n869), .B(n858), .CI(n854), .CO(n849), .S(n850) );
  FADDX1_LVT U811 ( .A(n1990), .B(n873), .CI(n871), .CO(n851), .S(n852) );
  FADDX1_LVT U812 ( .A(n2054), .B(n1862), .CI(n1926), .CO(n853), .S(n854) );
  FADDX1_LVT U813 ( .A(n2118), .B(n1734), .CI(n1798), .CO(n855), .S(n856) );
  FADDX1_LVT U814 ( .A(I3[54]), .B(n1670), .CI(n2182), .CO(n857), .S(n858) );
  FADDX1_LVT U815 ( .A(n864), .B(n877), .CI(n862), .CO(n859), .S(n860) );
  FADDX1_LVT U816 ( .A(n868), .B(n866), .CI(n879), .CO(n861), .S(n862) );
  FADDX1_LVT U817 ( .A(n872), .B(n883), .CI(n881), .CO(n863), .S(n864) );
  FADDX1_LVT U818 ( .A(n885), .B(n874), .CI(n870), .CO(n865), .S(n866) );
  FADDX1_LVT U819 ( .A(n1991), .B(n889), .CI(n887), .CO(n867), .S(n868) );
  FADDX1_LVT U820 ( .A(n2055), .B(n1863), .CI(n1927), .CO(n869), .S(n870) );
  FADDX1_LVT U821 ( .A(n2119), .B(n1735), .CI(n1799), .CO(n871), .S(n872) );
  FADDX1_LVT U822 ( .A(I3[53]), .B(n1671), .CI(n2183), .CO(n873), .S(n874) );
  FADDX1_LVT U823 ( .A(n880), .B(n893), .CI(n878), .CO(n875), .S(n876) );
  FADDX1_LVT U824 ( .A(n884), .B(n882), .CI(n895), .CO(n877), .S(n878) );
  FADDX1_LVT U825 ( .A(n888), .B(n899), .CI(n897), .CO(n879), .S(n880) );
  FADDX1_LVT U826 ( .A(n901), .B(n890), .CI(n886), .CO(n881), .S(n882) );
  FADDX1_LVT U827 ( .A(n1992), .B(n905), .CI(n903), .CO(n883), .S(n884) );
  FADDX1_LVT U828 ( .A(n2056), .B(n1864), .CI(n1928), .CO(n885), .S(n886) );
  FADDX1_LVT U829 ( .A(n2120), .B(n1736), .CI(n1800), .CO(n887), .S(n888) );
  FADDX1_LVT U830 ( .A(I3[52]), .B(n1672), .CI(n2184), .CO(n889), .S(n890) );
  FADDX1_LVT U831 ( .A(n896), .B(n909), .CI(n894), .CO(n891), .S(n892) );
  FADDX1_LVT U832 ( .A(n900), .B(n898), .CI(n911), .CO(n893), .S(n894) );
  FADDX1_LVT U833 ( .A(n904), .B(n915), .CI(n913), .CO(n895), .S(n896) );
  FADDX1_LVT U834 ( .A(n917), .B(n906), .CI(n902), .CO(n897), .S(n898) );
  FADDX1_LVT U835 ( .A(n1993), .B(n921), .CI(n919), .CO(n899), .S(n900) );
  FADDX1_LVT U836 ( .A(n2057), .B(n1865), .CI(n1929), .CO(n901), .S(n902) );
  FADDX1_LVT U837 ( .A(n2121), .B(n1737), .CI(n1801), .CO(n903), .S(n904) );
  FADDX1_LVT U838 ( .A(I3[51]), .B(n1673), .CI(n2185), .CO(n905), .S(n906) );
  FADDX1_LVT U839 ( .A(n912), .B(n925), .CI(n910), .CO(n907), .S(n908) );
  FADDX1_LVT U840 ( .A(n916), .B(n914), .CI(n927), .CO(n909), .S(n910) );
  FADDX1_LVT U841 ( .A(n920), .B(n931), .CI(n929), .CO(n911), .S(n912) );
  FADDX1_LVT U842 ( .A(n933), .B(n922), .CI(n918), .CO(n913), .S(n914) );
  FADDX1_LVT U843 ( .A(n1994), .B(n937), .CI(n935), .CO(n915), .S(n916) );
  FADDX1_LVT U844 ( .A(n2058), .B(n1866), .CI(n1930), .CO(n917), .S(n918) );
  FADDX1_LVT U845 ( .A(n2122), .B(n1738), .CI(n1802), .CO(n919), .S(n920) );
  FADDX1_LVT U846 ( .A(I3[50]), .B(n1674), .CI(n2186), .CO(n921), .S(n922) );
  FADDX1_LVT U847 ( .A(n928), .B(n941), .CI(n926), .CO(n923), .S(n924) );
  FADDX1_LVT U848 ( .A(n932), .B(n930), .CI(n943), .CO(n925), .S(n926) );
  FADDX1_LVT U849 ( .A(n936), .B(n947), .CI(n945), .CO(n927), .S(n928) );
  FADDX1_LVT U850 ( .A(n949), .B(n938), .CI(n934), .CO(n929), .S(n930) );
  FADDX1_LVT U851 ( .A(n1995), .B(n953), .CI(n951), .CO(n931), .S(n932) );
  FADDX1_LVT U852 ( .A(n2059), .B(n1867), .CI(n1931), .CO(n933), .S(n934) );
  FADDX1_LVT U853 ( .A(n2123), .B(n1739), .CI(n1803), .CO(n935), .S(n936) );
  FADDX1_LVT U854 ( .A(I3[49]), .B(n1675), .CI(n2187), .CO(n937), .S(n938) );
  FADDX1_LVT U855 ( .A(n944), .B(n957), .CI(n942), .CO(n939), .S(n940) );
  FADDX1_LVT U856 ( .A(n948), .B(n946), .CI(n959), .CO(n941), .S(n942) );
  FADDX1_LVT U857 ( .A(n952), .B(n963), .CI(n961), .CO(n943), .S(n944) );
  FADDX1_LVT U858 ( .A(n965), .B(n954), .CI(n950), .CO(n945), .S(n946) );
  FADDX1_LVT U859 ( .A(n1996), .B(n969), .CI(n967), .CO(n947), .S(n948) );
  FADDX1_LVT U860 ( .A(n2060), .B(n1868), .CI(n1932), .CO(n949), .S(n950) );
  FADDX1_LVT U861 ( .A(n2124), .B(n1740), .CI(n1804), .CO(n951), .S(n952) );
  FADDX1_LVT U862 ( .A(I3[48]), .B(n1676), .CI(n2188), .CO(n953), .S(n954) );
  FADDX1_LVT U863 ( .A(n960), .B(n973), .CI(n958), .CO(n955), .S(n956) );
  FADDX1_LVT U864 ( .A(n964), .B(n962), .CI(n975), .CO(n957), .S(n958) );
  FADDX1_LVT U865 ( .A(n968), .B(n979), .CI(n977), .CO(n959), .S(n960) );
  FADDX1_LVT U866 ( .A(n981), .B(n970), .CI(n966), .CO(n961), .S(n962) );
  FADDX1_LVT U867 ( .A(n1997), .B(n985), .CI(n983), .CO(n963), .S(n964) );
  FADDX1_LVT U868 ( .A(n2061), .B(n1869), .CI(n1933), .CO(n965), .S(n966) );
  FADDX1_LVT U869 ( .A(n2125), .B(n1741), .CI(n1805), .CO(n967), .S(n968) );
  FADDX1_LVT U870 ( .A(I3[47]), .B(n1677), .CI(n2189), .CO(n969), .S(n970) );
  FADDX1_LVT U871 ( .A(n976), .B(n989), .CI(n974), .CO(n971), .S(n972) );
  FADDX1_LVT U872 ( .A(n980), .B(n978), .CI(n991), .CO(n973), .S(n974) );
  FADDX1_LVT U873 ( .A(n984), .B(n995), .CI(n993), .CO(n975), .S(n976) );
  FADDX1_LVT U874 ( .A(n997), .B(n986), .CI(n982), .CO(n977), .S(n978) );
  FADDX1_LVT U875 ( .A(n1998), .B(n1001), .CI(n999), .CO(n979), .S(n980) );
  FADDX1_LVT U876 ( .A(n2062), .B(n1870), .CI(n1934), .CO(n981), .S(n982) );
  FADDX1_LVT U877 ( .A(n2126), .B(n1742), .CI(n1806), .CO(n983), .S(n984) );
  FADDX1_LVT U878 ( .A(I3[46]), .B(n1678), .CI(n2190), .CO(n985), .S(n986) );
  FADDX1_LVT U879 ( .A(n992), .B(n1005), .CI(n990), .CO(n987), .S(n988) );
  FADDX1_LVT U880 ( .A(n996), .B(n994), .CI(n1007), .CO(n989), .S(n990) );
  FADDX1_LVT U881 ( .A(n1000), .B(n1011), .CI(n1009), .CO(n991), .S(n992) );
  FADDX1_LVT U882 ( .A(n1013), .B(n1002), .CI(n998), .CO(n993), .S(n994) );
  FADDX1_LVT U883 ( .A(n1999), .B(n1017), .CI(n1015), .CO(n995), .S(n996) );
  FADDX1_LVT U884 ( .A(n2063), .B(n1871), .CI(n1935), .CO(n997), .S(n998) );
  FADDX1_LVT U885 ( .A(n2127), .B(n1743), .CI(n1807), .CO(n999), .S(n1000) );
  FADDX1_LVT U886 ( .A(I3[45]), .B(n1679), .CI(n2191), .CO(n1001), .S(n1002)
         );
  FADDX1_LVT U887 ( .A(n1008), .B(n1021), .CI(n1006), .CO(n1003), .S(n1004) );
  FADDX1_LVT U888 ( .A(n1012), .B(n1010), .CI(n1023), .CO(n1005), .S(n1006) );
  FADDX1_LVT U889 ( .A(n1016), .B(n1027), .CI(n1025), .CO(n1007), .S(n1008) );
  FADDX1_LVT U890 ( .A(n1029), .B(n1018), .CI(n1014), .CO(n1009), .S(n1010) );
  FADDX1_LVT U891 ( .A(n2000), .B(n1033), .CI(n1031), .CO(n1011), .S(n1012) );
  FADDX1_LVT U892 ( .A(n2064), .B(n1872), .CI(n1936), .CO(n1013), .S(n1014) );
  FADDX1_LVT U893 ( .A(n2128), .B(n1744), .CI(n1808), .CO(n1015), .S(n1016) );
  FADDX1_LVT U894 ( .A(I3[44]), .B(n1680), .CI(n2192), .CO(n1017), .S(n1018)
         );
  FADDX1_LVT U895 ( .A(n1024), .B(n1037), .CI(n1022), .CO(n1019), .S(n1020) );
  FADDX1_LVT U896 ( .A(n1028), .B(n1026), .CI(n1039), .CO(n1021), .S(n1022) );
  FADDX1_LVT U897 ( .A(n1032), .B(n1043), .CI(n1041), .CO(n1023), .S(n1024) );
  FADDX1_LVT U898 ( .A(n1045), .B(n1034), .CI(n1030), .CO(n1025), .S(n1026) );
  FADDX1_LVT U899 ( .A(n2001), .B(n1049), .CI(n1047), .CO(n1027), .S(n1028) );
  FADDX1_LVT U900 ( .A(n2065), .B(n1873), .CI(n1937), .CO(n1029), .S(n1030) );
  FADDX1_LVT U901 ( .A(n2129), .B(n1745), .CI(n1809), .CO(n1031), .S(n1032) );
  FADDX1_LVT U902 ( .A(I3[43]), .B(n1681), .CI(n2193), .CO(n1033), .S(n1034)
         );
  FADDX1_LVT U903 ( .A(n1040), .B(n1053), .CI(n1038), .CO(n1035), .S(n1036) );
  FADDX1_LVT U904 ( .A(n1044), .B(n1042), .CI(n1055), .CO(n1037), .S(n1038) );
  FADDX1_LVT U905 ( .A(n1048), .B(n1059), .CI(n1057), .CO(n1039), .S(n1040) );
  FADDX1_LVT U906 ( .A(n1061), .B(n1050), .CI(n1046), .CO(n1041), .S(n1042) );
  FADDX1_LVT U907 ( .A(n2002), .B(n1065), .CI(n1063), .CO(n1043), .S(n1044) );
  FADDX1_LVT U908 ( .A(n2066), .B(n1874), .CI(n1938), .CO(n1045), .S(n1046) );
  FADDX1_LVT U909 ( .A(n2130), .B(n1746), .CI(n1810), .CO(n1047), .S(n1048) );
  FADDX1_LVT U910 ( .A(I3[42]), .B(n1682), .CI(n2194), .CO(n1049), .S(n1050)
         );
  FADDX1_LVT U911 ( .A(n1056), .B(n1069), .CI(n1054), .CO(n1051), .S(n1052) );
  FADDX1_LVT U912 ( .A(n1060), .B(n1058), .CI(n1071), .CO(n1053), .S(n1054) );
  FADDX1_LVT U913 ( .A(n1064), .B(n1075), .CI(n1073), .CO(n1055), .S(n1056) );
  FADDX1_LVT U914 ( .A(n1077), .B(n1066), .CI(n1062), .CO(n1057), .S(n1058) );
  FADDX1_LVT U915 ( .A(n2003), .B(n1081), .CI(n1079), .CO(n1059), .S(n1060) );
  FADDX1_LVT U916 ( .A(n2067), .B(n1875), .CI(n1939), .CO(n1061), .S(n1062) );
  FADDX1_LVT U917 ( .A(n2131), .B(n1747), .CI(n1811), .CO(n1063), .S(n1064) );
  FADDX1_LVT U918 ( .A(I3[41]), .B(n1683), .CI(n2195), .CO(n1065), .S(n1066)
         );
  FADDX1_LVT U919 ( .A(n1072), .B(n1085), .CI(n1070), .CO(n1067), .S(n1068) );
  FADDX1_LVT U920 ( .A(n1076), .B(n1074), .CI(n1087), .CO(n1069), .S(n1070) );
  FADDX1_LVT U921 ( .A(n1080), .B(n1091), .CI(n1089), .CO(n1071), .S(n1072) );
  FADDX1_LVT U922 ( .A(n1093), .B(n1082), .CI(n1078), .CO(n1073), .S(n1074) );
  FADDX1_LVT U923 ( .A(n2004), .B(n1097), .CI(n1095), .CO(n1075), .S(n1076) );
  FADDX1_LVT U924 ( .A(n2068), .B(n1876), .CI(n1940), .CO(n1077), .S(n1078) );
  FADDX1_LVT U925 ( .A(n2132), .B(n1748), .CI(n1812), .CO(n1079), .S(n1080) );
  FADDX1_LVT U926 ( .A(I3[40]), .B(n1684), .CI(n2196), .CO(n1081), .S(n1082)
         );
  FADDX1_LVT U927 ( .A(n1088), .B(n1101), .CI(n1086), .CO(n1083), .S(n1084) );
  FADDX1_LVT U928 ( .A(n1092), .B(n1090), .CI(n1103), .CO(n1085), .S(n1086) );
  FADDX1_LVT U929 ( .A(n1096), .B(n1107), .CI(n1105), .CO(n1087), .S(n1088) );
  FADDX1_LVT U930 ( .A(n1109), .B(n1098), .CI(n1094), .CO(n1089), .S(n1090) );
  FADDX1_LVT U931 ( .A(n2005), .B(n1113), .CI(n1111), .CO(n1091), .S(n1092) );
  FADDX1_LVT U932 ( .A(n2069), .B(n1877), .CI(n1941), .CO(n1093), .S(n1094) );
  FADDX1_LVT U933 ( .A(n2133), .B(n1749), .CI(n1813), .CO(n1095), .S(n1096) );
  FADDX1_LVT U934 ( .A(I3[39]), .B(n1685), .CI(n2197), .CO(n1097), .S(n1098)
         );
  FADDX1_LVT U935 ( .A(n1104), .B(n1117), .CI(n1102), .CO(n1099), .S(n1100) );
  FADDX1_LVT U936 ( .A(n1108), .B(n1106), .CI(n1119), .CO(n1101), .S(n1102) );
  FADDX1_LVT U937 ( .A(n1112), .B(n1123), .CI(n1121), .CO(n1103), .S(n1104) );
  FADDX1_LVT U938 ( .A(n1125), .B(n1114), .CI(n1110), .CO(n1105), .S(n1106) );
  FADDX1_LVT U939 ( .A(n2006), .B(n1129), .CI(n1127), .CO(n1107), .S(n1108) );
  FADDX1_LVT U940 ( .A(n2070), .B(n1878), .CI(n1942), .CO(n1109), .S(n1110) );
  FADDX1_LVT U941 ( .A(n2134), .B(n1750), .CI(n1814), .CO(n1111), .S(n1112) );
  FADDX1_LVT U942 ( .A(I3[38]), .B(n1686), .CI(n2198), .CO(n1113), .S(n1114)
         );
  FADDX1_LVT U943 ( .A(n1120), .B(n1133), .CI(n1118), .CO(n1115), .S(n1116) );
  FADDX1_LVT U944 ( .A(n1124), .B(n1122), .CI(n1135), .CO(n1117), .S(n1118) );
  FADDX1_LVT U945 ( .A(n1128), .B(n1139), .CI(n1137), .CO(n1119), .S(n1120) );
  FADDX1_LVT U946 ( .A(n1141), .B(n1130), .CI(n1126), .CO(n1121), .S(n1122) );
  FADDX1_LVT U947 ( .A(n2007), .B(n1145), .CI(n1143), .CO(n1123), .S(n1124) );
  FADDX1_LVT U948 ( .A(n2071), .B(n1879), .CI(n1943), .CO(n1125), .S(n1126) );
  FADDX1_LVT U949 ( .A(n2135), .B(n1751), .CI(n1815), .CO(n1127), .S(n1128) );
  FADDX1_LVT U950 ( .A(I3[37]), .B(n1687), .CI(n2199), .CO(n1129), .S(n1130)
         );
  FADDX1_LVT U951 ( .A(n1136), .B(n1149), .CI(n1134), .CO(n1131), .S(n1132) );
  FADDX1_LVT U952 ( .A(n1140), .B(n1138), .CI(n1151), .CO(n1133), .S(n1134) );
  FADDX1_LVT U953 ( .A(n1144), .B(n1155), .CI(n1153), .CO(n1135), .S(n1136) );
  FADDX1_LVT U954 ( .A(n1157), .B(n1146), .CI(n1142), .CO(n1137), .S(n1138) );
  FADDX1_LVT U955 ( .A(n2008), .B(n1161), .CI(n1159), .CO(n1139), .S(n1140) );
  FADDX1_LVT U956 ( .A(n2072), .B(n1880), .CI(n1944), .CO(n1141), .S(n1142) );
  FADDX1_LVT U957 ( .A(n2136), .B(n1752), .CI(n1816), .CO(n1143), .S(n1144) );
  FADDX1_LVT U958 ( .A(I3[36]), .B(n1688), .CI(n2200), .CO(n1145), .S(n1146)
         );
  FADDX1_LVT U959 ( .A(n1152), .B(n1165), .CI(n1150), .CO(n1147), .S(n1148) );
  FADDX1_LVT U960 ( .A(n1156), .B(n1154), .CI(n1167), .CO(n1149), .S(n1150) );
  FADDX1_LVT U961 ( .A(n1160), .B(n1171), .CI(n1169), .CO(n1151), .S(n1152) );
  FADDX1_LVT U962 ( .A(n1173), .B(n1162), .CI(n1158), .CO(n1153), .S(n1154) );
  FADDX1_LVT U963 ( .A(n2009), .B(n1177), .CI(n1175), .CO(n1155), .S(n1156) );
  FADDX1_LVT U964 ( .A(n2073), .B(n1881), .CI(n1945), .CO(n1157), .S(n1158) );
  FADDX1_LVT U965 ( .A(n2137), .B(n1753), .CI(n1817), .CO(n1159), .S(n1160) );
  FADDX1_LVT U966 ( .A(I3[35]), .B(n1689), .CI(n2201), .CO(n1161), .S(n1162)
         );
  FADDX1_LVT U967 ( .A(n1168), .B(n1181), .CI(n1166), .CO(n1163), .S(n1164) );
  FADDX1_LVT U968 ( .A(n1172), .B(n1170), .CI(n1183), .CO(n1165), .S(n1166) );
  FADDX1_LVT U969 ( .A(n1176), .B(n1187), .CI(n1185), .CO(n1167), .S(n1168) );
  FADDX1_LVT U970 ( .A(n1189), .B(n1178), .CI(n1174), .CO(n1169), .S(n1170) );
  FADDX1_LVT U971 ( .A(n2010), .B(n1193), .CI(n1191), .CO(n1171), .S(n1172) );
  FADDX1_LVT U972 ( .A(n2074), .B(n1882), .CI(n1946), .CO(n1173), .S(n1174) );
  FADDX1_LVT U973 ( .A(n2138), .B(n1754), .CI(n1818), .CO(n1175), .S(n1176) );
  FADDX1_LVT U974 ( .A(I3[34]), .B(n1690), .CI(n2202), .CO(n1177), .S(n1178)
         );
  FADDX1_LVT U975 ( .A(n1184), .B(n1197), .CI(n1182), .CO(n1179), .S(n1180) );
  FADDX1_LVT U976 ( .A(n1188), .B(n1186), .CI(n1199), .CO(n1181), .S(n1182) );
  FADDX1_LVT U977 ( .A(n1192), .B(n1203), .CI(n1201), .CO(n1183), .S(n1184) );
  FADDX1_LVT U978 ( .A(n1205), .B(n1194), .CI(n1190), .CO(n1185), .S(n1186) );
  FADDX1_LVT U979 ( .A(n2011), .B(n1209), .CI(n1207), .CO(n1187), .S(n1188) );
  FADDX1_LVT U980 ( .A(n2075), .B(n1883), .CI(n1947), .CO(n1189), .S(n1190) );
  FADDX1_LVT U981 ( .A(n2139), .B(n1755), .CI(n1819), .CO(n1191), .S(n1192) );
  FADDX1_LVT U982 ( .A(I3[33]), .B(n1691), .CI(n2203), .CO(n1193), .S(n1194)
         );
  FADDX1_LVT U983 ( .A(n1200), .B(n1213), .CI(n1198), .CO(n1195), .S(n1196) );
  FADDX1_LVT U984 ( .A(n1204), .B(n1202), .CI(n1215), .CO(n1197), .S(n1198) );
  FADDX1_LVT U985 ( .A(n1208), .B(n1219), .CI(n1217), .CO(n1199), .S(n1200) );
  FADDX1_LVT U986 ( .A(n1221), .B(n1210), .CI(n1206), .CO(n1201), .S(n1202) );
  FADDX1_LVT U987 ( .A(n2012), .B(n1225), .CI(n1223), .CO(n1203), .S(n1204) );
  FADDX1_LVT U988 ( .A(n2076), .B(n1884), .CI(n1948), .CO(n1205), .S(n1206) );
  FADDX1_LVT U989 ( .A(n2140), .B(n1756), .CI(n1820), .CO(n1207), .S(n1208) );
  FADDX1_LVT U990 ( .A(I3[32]), .B(n1692), .CI(n2204), .CO(n1209), .S(n1210)
         );
  FADDX1_LVT U991 ( .A(n1216), .B(n1229), .CI(n1214), .CO(n1211), .S(n1212) );
  FADDX1_LVT U992 ( .A(n1220), .B(n1218), .CI(n1231), .CO(n1213), .S(n1214) );
  FADDX1_LVT U993 ( .A(n1224), .B(n1235), .CI(n1233), .CO(n1215), .S(n1216) );
  FADDX1_LVT U994 ( .A(n1237), .B(n1226), .CI(n1222), .CO(n1217), .S(n1218) );
  FADDX1_LVT U995 ( .A(n2013), .B(n1241), .CI(n1239), .CO(n1219), .S(n1220) );
  FADDX1_LVT U996 ( .A(n2077), .B(n1885), .CI(n1949), .CO(n1221), .S(n1222) );
  FADDX1_LVT U997 ( .A(n2141), .B(n1757), .CI(n1821), .CO(n1223), .S(n1224) );
  FADDX1_LVT U998 ( .A(I3[31]), .B(n1693), .CI(n2205), .CO(n1225), .S(n1226)
         );
  FADDX1_LVT U999 ( .A(n1232), .B(n1245), .CI(n1230), .CO(n1227), .S(n1228) );
  FADDX1_LVT U1000 ( .A(n1236), .B(n1234), .CI(n1247), .CO(n1229), .S(n1230)
         );
  FADDX1_LVT U1001 ( .A(n1240), .B(n1251), .CI(n1249), .CO(n1231), .S(n1232)
         );
  FADDX1_LVT U1002 ( .A(n1253), .B(n1242), .CI(n1238), .CO(n1233), .S(n1234)
         );
  FADDX1_LVT U1003 ( .A(n2014), .B(n1257), .CI(n1255), .CO(n1235), .S(n1236)
         );
  FADDX1_LVT U1004 ( .A(n2078), .B(n1886), .CI(n1950), .CO(n1237), .S(n1238)
         );
  FADDX1_LVT U1005 ( .A(n2142), .B(n1758), .CI(n1822), .CO(n1239), .S(n1240)
         );
  FADDX1_LVT U1006 ( .A(I3[30]), .B(n1694), .CI(n2206), .CO(n1241), .S(n1242)
         );
  FADDX1_LVT U1007 ( .A(n1248), .B(n1261), .CI(n1246), .CO(n1243), .S(n1244)
         );
  FADDX1_LVT U1008 ( .A(n1252), .B(n1250), .CI(n1263), .CO(n1245), .S(n1246)
         );
  FADDX1_LVT U1009 ( .A(n1256), .B(n1267), .CI(n1265), .CO(n1247), .S(n1248)
         );
  FADDX1_LVT U1010 ( .A(n1269), .B(n1258), .CI(n1254), .CO(n1249), .S(n1250)
         );
  FADDX1_LVT U1011 ( .A(n2015), .B(n1273), .CI(n1271), .CO(n1251), .S(n1252)
         );
  FADDX1_LVT U1012 ( .A(n2079), .B(n1887), .CI(n1951), .CO(n1253), .S(n1254)
         );
  FADDX1_LVT U1013 ( .A(n2143), .B(n1759), .CI(n1823), .CO(n1255), .S(n1256)
         );
  FADDX1_LVT U1014 ( .A(I3[29]), .B(n1695), .CI(n2207), .CO(n1257), .S(n1258)
         );
  FADDX1_LVT U1015 ( .A(n1264), .B(n1277), .CI(n1262), .CO(n1259), .S(n1260)
         );
  FADDX1_LVT U1016 ( .A(n1268), .B(n1266), .CI(n1279), .CO(n1261), .S(n1262)
         );
  FADDX1_LVT U1017 ( .A(n1272), .B(n1283), .CI(n1281), .CO(n1263), .S(n1264)
         );
  FADDX1_LVT U1018 ( .A(n1285), .B(n1274), .CI(n1270), .CO(n1265), .S(n1266)
         );
  FADDX1_LVT U1019 ( .A(n2016), .B(n1289), .CI(n1287), .CO(n1267), .S(n1268)
         );
  FADDX1_LVT U1020 ( .A(n2080), .B(n1888), .CI(n1952), .CO(n1269), .S(n1270)
         );
  FADDX1_LVT U1021 ( .A(n2144), .B(n1760), .CI(n1824), .CO(n1271), .S(n1272)
         );
  FADDX1_LVT U1022 ( .A(I3[28]), .B(n1696), .CI(n2208), .CO(n1273), .S(n1274)
         );
  FADDX1_LVT U1023 ( .A(n1280), .B(n1293), .CI(n1278), .CO(n1275), .S(n1276)
         );
  FADDX1_LVT U1024 ( .A(n1284), .B(n1282), .CI(n1295), .CO(n1277), .S(n1278)
         );
  FADDX1_LVT U1025 ( .A(n1288), .B(n1299), .CI(n1297), .CO(n1279), .S(n1280)
         );
  FADDX1_LVT U1026 ( .A(n1301), .B(n1290), .CI(n1286), .CO(n1281), .S(n1282)
         );
  FADDX1_LVT U1027 ( .A(n2017), .B(n1305), .CI(n1303), .CO(n1283), .S(n1284)
         );
  FADDX1_LVT U1028 ( .A(n2081), .B(n1889), .CI(n1953), .CO(n1285), .S(n1286)
         );
  FADDX1_LVT U1029 ( .A(n2145), .B(n1761), .CI(n1825), .CO(n1287), .S(n1288)
         );
  FADDX1_LVT U1030 ( .A(I3[27]), .B(n1697), .CI(n2209), .CO(n1289), .S(n1290)
         );
  FADDX1_LVT U1031 ( .A(n1296), .B(n1309), .CI(n1294), .CO(n1291), .S(n1292)
         );
  FADDX1_LVT U1032 ( .A(n1300), .B(n1298), .CI(n1311), .CO(n1293), .S(n1294)
         );
  FADDX1_LVT U1033 ( .A(n1304), .B(n1315), .CI(n1313), .CO(n1295), .S(n1296)
         );
  FADDX1_LVT U1034 ( .A(n1317), .B(n1306), .CI(n1302), .CO(n1297), .S(n1298)
         );
  FADDX1_LVT U1035 ( .A(n2018), .B(n1321), .CI(n1319), .CO(n1299), .S(n1300)
         );
  FADDX1_LVT U1036 ( .A(n2082), .B(n1890), .CI(n1954), .CO(n1301), .S(n1302)
         );
  FADDX1_LVT U1037 ( .A(n2146), .B(n1762), .CI(n1826), .CO(n1303), .S(n1304)
         );
  FADDX1_LVT U1038 ( .A(I3[26]), .B(n1698), .CI(n2210), .CO(n1305), .S(n1306)
         );
  FADDX1_LVT U1039 ( .A(n1312), .B(n1325), .CI(n1310), .CO(n1307), .S(n1308)
         );
  FADDX1_LVT U1040 ( .A(n1316), .B(n1314), .CI(n1327), .CO(n1309), .S(n1310)
         );
  FADDX1_LVT U1041 ( .A(n1320), .B(n1331), .CI(n1329), .CO(n1311), .S(n1312)
         );
  FADDX1_LVT U1042 ( .A(n1333), .B(n1322), .CI(n1318), .CO(n1313), .S(n1314)
         );
  FADDX1_LVT U1043 ( .A(n2019), .B(n1337), .CI(n1335), .CO(n1315), .S(n1316)
         );
  FADDX1_LVT U1044 ( .A(n2083), .B(n1891), .CI(n1955), .CO(n1317), .S(n1318)
         );
  FADDX1_LVT U1045 ( .A(n2147), .B(n1763), .CI(n1827), .CO(n1319), .S(n1320)
         );
  FADDX1_LVT U1046 ( .A(I3[25]), .B(n1699), .CI(n2211), .CO(n1321), .S(n1322)
         );
  FADDX1_LVT U1047 ( .A(n1328), .B(n1341), .CI(n1326), .CO(n1323), .S(n1324)
         );
  FADDX1_LVT U1048 ( .A(n1332), .B(n1330), .CI(n1343), .CO(n1325), .S(n1326)
         );
  FADDX1_LVT U1049 ( .A(n1336), .B(n1347), .CI(n1345), .CO(n1327), .S(n1328)
         );
  FADDX1_LVT U1050 ( .A(n1349), .B(n1338), .CI(n1334), .CO(n1329), .S(n1330)
         );
  FADDX1_LVT U1051 ( .A(n2020), .B(n1353), .CI(n1351), .CO(n1331), .S(n1332)
         );
  FADDX1_LVT U1052 ( .A(n2084), .B(n1892), .CI(n1956), .CO(n1333), .S(n1334)
         );
  FADDX1_LVT U1053 ( .A(n2148), .B(n1764), .CI(n1828), .CO(n1335), .S(n1336)
         );
  FADDX1_LVT U1054 ( .A(I3[24]), .B(n1700), .CI(n2212), .CO(n1337), .S(n1338)
         );
  FADDX1_LVT U1055 ( .A(n1344), .B(n1357), .CI(n1342), .CO(n1339), .S(n1340)
         );
  FADDX1_LVT U1056 ( .A(n1348), .B(n1346), .CI(n1359), .CO(n1341), .S(n1342)
         );
  FADDX1_LVT U1057 ( .A(n1352), .B(n1363), .CI(n1361), .CO(n1343), .S(n1344)
         );
  FADDX1_LVT U1058 ( .A(n1365), .B(n1354), .CI(n1350), .CO(n1345), .S(n1346)
         );
  FADDX1_LVT U1059 ( .A(n2021), .B(n1369), .CI(n1367), .CO(n1347), .S(n1348)
         );
  FADDX1_LVT U1060 ( .A(n2085), .B(n1893), .CI(n1957), .CO(n1349), .S(n1350)
         );
  FADDX1_LVT U1061 ( .A(n2149), .B(n1765), .CI(n1829), .CO(n1351), .S(n1352)
         );
  FADDX1_LVT U1062 ( .A(I3[23]), .B(n1701), .CI(n2213), .CO(n1353), .S(n1354)
         );
  FADDX1_LVT U1063 ( .A(n1360), .B(n1373), .CI(n1358), .CO(n1355), .S(n1356)
         );
  FADDX1_LVT U1064 ( .A(n1364), .B(n1362), .CI(n1375), .CO(n1357), .S(n1358)
         );
  FADDX1_LVT U1065 ( .A(n1368), .B(n1379), .CI(n1377), .CO(n1359), .S(n1360)
         );
  FADDX1_LVT U1066 ( .A(n1381), .B(n1370), .CI(n1366), .CO(n1361), .S(n1362)
         );
  FADDX1_LVT U1067 ( .A(n2022), .B(n1385), .CI(n1383), .CO(n1363), .S(n1364)
         );
  FADDX1_LVT U1068 ( .A(n2086), .B(n1894), .CI(n1958), .CO(n1365), .S(n1366)
         );
  FADDX1_LVT U1069 ( .A(n2150), .B(n1766), .CI(n1830), .CO(n1367), .S(n1368)
         );
  FADDX1_LVT U1070 ( .A(I3[22]), .B(n1702), .CI(n2214), .CO(n1369), .S(n1370)
         );
  FADDX1_LVT U1071 ( .A(n1376), .B(n1389), .CI(n1374), .CO(n1371), .S(n1372)
         );
  FADDX1_LVT U1072 ( .A(n1380), .B(n1378), .CI(n1391), .CO(n1373), .S(n1374)
         );
  FADDX1_LVT U1073 ( .A(n1384), .B(n1395), .CI(n1393), .CO(n1375), .S(n1376)
         );
  FADDX1_LVT U1074 ( .A(n1397), .B(n1386), .CI(n1382), .CO(n1377), .S(n1378)
         );
  FADDX1_LVT U1075 ( .A(n2023), .B(n1401), .CI(n1399), .CO(n1379), .S(n1380)
         );
  FADDX1_LVT U1076 ( .A(n2087), .B(n1895), .CI(n1959), .CO(n1381), .S(n1382)
         );
  FADDX1_LVT U1077 ( .A(n2151), .B(n1767), .CI(n1831), .CO(n1383), .S(n1384)
         );
  FADDX1_LVT U1078 ( .A(I3[21]), .B(n1703), .CI(n2215), .CO(n1385), .S(n1386)
         );
  FADDX1_LVT U1079 ( .A(n1392), .B(n1405), .CI(n1390), .CO(n1387), .S(n1388)
         );
  FADDX1_LVT U1080 ( .A(n1396), .B(n1394), .CI(n1407), .CO(n1389), .S(n1390)
         );
  FADDX1_LVT U1081 ( .A(n1400), .B(n1411), .CI(n1409), .CO(n1391), .S(n1392)
         );
  FADDX1_LVT U1082 ( .A(n1413), .B(n1402), .CI(n1398), .CO(n1393), .S(n1394)
         );
  FADDX1_LVT U1083 ( .A(n2024), .B(n1417), .CI(n1415), .CO(n1395), .S(n1396)
         );
  FADDX1_LVT U1084 ( .A(n2088), .B(n1896), .CI(n1960), .CO(n1397), .S(n1398)
         );
  FADDX1_LVT U1085 ( .A(n2152), .B(n1768), .CI(n1832), .CO(n1399), .S(n1400)
         );
  FADDX1_LVT U1086 ( .A(I3[20]), .B(n1704), .CI(n2216), .CO(n1401), .S(n1402)
         );
  FADDX1_LVT U1087 ( .A(n1408), .B(n1421), .CI(n1406), .CO(n1403), .S(n1404)
         );
  FADDX1_LVT U1088 ( .A(n1412), .B(n1410), .CI(n1423), .CO(n1405), .S(n1406)
         );
  FADDX1_LVT U1089 ( .A(n1416), .B(n1427), .CI(n1425), .CO(n1407), .S(n1408)
         );
  FADDX1_LVT U1090 ( .A(n1429), .B(n1418), .CI(n1414), .CO(n1409), .S(n1410)
         );
  FADDX1_LVT U1091 ( .A(n2025), .B(n1433), .CI(n1431), .CO(n1411), .S(n1412)
         );
  FADDX1_LVT U1092 ( .A(n2089), .B(n1897), .CI(n1961), .CO(n1413), .S(n1414)
         );
  FADDX1_LVT U1093 ( .A(n2153), .B(n1769), .CI(n1833), .CO(n1415), .S(n1416)
         );
  FADDX1_LVT U1094 ( .A(I3[19]), .B(n1705), .CI(n2217), .CO(n1417), .S(n1418)
         );
  FADDX1_LVT U1095 ( .A(n1424), .B(n1437), .CI(n1422), .CO(n1419), .S(n1420)
         );
  FADDX1_LVT U1096 ( .A(n1428), .B(n1426), .CI(n1439), .CO(n1421), .S(n1422)
         );
  FADDX1_LVT U1097 ( .A(n1432), .B(n1443), .CI(n1441), .CO(n1423), .S(n1424)
         );
  FADDX1_LVT U1098 ( .A(n1445), .B(n1434), .CI(n1430), .CO(n1425), .S(n1426)
         );
  FADDX1_LVT U1099 ( .A(n2026), .B(n1449), .CI(n1447), .CO(n1427), .S(n1428)
         );
  FADDX1_LVT U1100 ( .A(n2090), .B(n1898), .CI(n1962), .CO(n1429), .S(n1430)
         );
  FADDX1_LVT U1101 ( .A(n2154), .B(n1770), .CI(n1834), .CO(n1431), .S(n1432)
         );
  FADDX1_LVT U1102 ( .A(I3[18]), .B(n1706), .CI(n2218), .CO(n1433), .S(n1434)
         );
  FADDX1_LVT U1103 ( .A(n1440), .B(n1453), .CI(n1438), .CO(n1435), .S(n1436)
         );
  FADDX1_LVT U1104 ( .A(n1444), .B(n1442), .CI(n1455), .CO(n1437), .S(n1438)
         );
  FADDX1_LVT U1105 ( .A(n1448), .B(n1459), .CI(n1457), .CO(n1439), .S(n1440)
         );
  FADDX1_LVT U1106 ( .A(n1461), .B(n1450), .CI(n1446), .CO(n1441), .S(n1442)
         );
  FADDX1_LVT U1107 ( .A(n2027), .B(n1465), .CI(n1463), .CO(n1443), .S(n1444)
         );
  FADDX1_LVT U1108 ( .A(n2091), .B(n1899), .CI(n1963), .CO(n1445), .S(n1446)
         );
  FADDX1_LVT U1109 ( .A(n2155), .B(n1771), .CI(n1835), .CO(n1447), .S(n1448)
         );
  FADDX1_LVT U1110 ( .A(I3[17]), .B(n1707), .CI(n2219), .CO(n1449), .S(n1450)
         );
  FADDX1_LVT U1111 ( .A(n1456), .B(n1469), .CI(n1454), .CO(n1451), .S(n1452)
         );
  FADDX1_LVT U1112 ( .A(n1460), .B(n1458), .CI(n1471), .CO(n1453), .S(n1454)
         );
  FADDX1_LVT U1113 ( .A(n1464), .B(n1475), .CI(n1473), .CO(n1455), .S(n1456)
         );
  FADDX1_LVT U1114 ( .A(n1477), .B(n1466), .CI(n1462), .CO(n1457), .S(n1458)
         );
  FADDX1_LVT U1115 ( .A(n2028), .B(n1481), .CI(n1479), .CO(n1459), .S(n1460)
         );
  FADDX1_LVT U1116 ( .A(n2092), .B(n1900), .CI(n1964), .CO(n1461), .S(n1462)
         );
  FADDX1_LVT U1117 ( .A(n2156), .B(n1772), .CI(n1836), .CO(n1463), .S(n1464)
         );
  FADDX1_LVT U1118 ( .A(I3[16]), .B(n1708), .CI(n2220), .CO(n1465), .S(n1466)
         );
  FADDX1_LVT U1119 ( .A(n1472), .B(n1485), .CI(n1470), .CO(n1467), .S(n1468)
         );
  FADDX1_LVT U1120 ( .A(n1476), .B(n1474), .CI(n1487), .CO(n1469), .S(n1470)
         );
  FADDX1_LVT U1121 ( .A(n1480), .B(n1491), .CI(n1489), .CO(n1471), .S(n1472)
         );
  FADDX1_LVT U1122 ( .A(n1493), .B(n1482), .CI(n1478), .CO(n1473), .S(n1474)
         );
  FADDX1_LVT U1123 ( .A(n2029), .B(n1497), .CI(n1495), .CO(n1475), .S(n1476)
         );
  FADDX1_LVT U1124 ( .A(n2093), .B(n1901), .CI(n1965), .CO(n1477), .S(n1478)
         );
  FADDX1_LVT U1125 ( .A(n2157), .B(n1773), .CI(n1837), .CO(n1479), .S(n1480)
         );
  FADDX1_LVT U1126 ( .A(I3[15]), .B(n1709), .CI(n2221), .CO(n1481), .S(n1482)
         );
  FADDX1_LVT U1127 ( .A(n1488), .B(n1501), .CI(n1486), .CO(n1483), .S(n1484)
         );
  FADDX1_LVT U1128 ( .A(n1492), .B(n1490), .CI(n1503), .CO(n1485), .S(n1486)
         );
  FADDX1_LVT U1129 ( .A(n1496), .B(n1507), .CI(n1505), .CO(n1487), .S(n1488)
         );
  FADDX1_LVT U1130 ( .A(n1509), .B(n1498), .CI(n1494), .CO(n1489), .S(n1490)
         );
  FADDX1_LVT U1131 ( .A(n2030), .B(n1513), .CI(n1511), .CO(n1491), .S(n1492)
         );
  FADDX1_LVT U1132 ( .A(n2094), .B(n1902), .CI(n1966), .CO(n1493), .S(n1494)
         );
  FADDX1_LVT U1133 ( .A(n2158), .B(n1774), .CI(n1838), .CO(n1495), .S(n1496)
         );
  FADDX1_LVT U1134 ( .A(I3[14]), .B(n1710), .CI(n2222), .CO(n1497), .S(n1498)
         );
  FADDX1_LVT U1135 ( .A(n1504), .B(n1517), .CI(n1502), .CO(n1499), .S(n1500)
         );
  FADDX1_LVT U1136 ( .A(n1508), .B(n1506), .CI(n1519), .CO(n1501), .S(n1502)
         );
  FADDX1_LVT U1137 ( .A(n1512), .B(n1523), .CI(n1521), .CO(n1503), .S(n1504)
         );
  FADDX1_LVT U1138 ( .A(n1525), .B(n1514), .CI(n1510), .CO(n1505), .S(n1506)
         );
  FADDX1_LVT U1139 ( .A(n2031), .B(n1529), .CI(n1527), .CO(n1507), .S(n1508)
         );
  FADDX1_LVT U1140 ( .A(n2095), .B(n1903), .CI(n1967), .CO(n1509), .S(n1510)
         );
  FADDX1_LVT U1141 ( .A(n2159), .B(n1775), .CI(n1839), .CO(n1511), .S(n1512)
         );
  FADDX1_LVT U1142 ( .A(I3[13]), .B(n1711), .CI(n2223), .CO(n1513), .S(n1514)
         );
  FADDX1_LVT U1143 ( .A(n1520), .B(n1533), .CI(n1518), .CO(n1515), .S(n1516)
         );
  FADDX1_LVT U1144 ( .A(n1524), .B(n1522), .CI(n1535), .CO(n1517), .S(n1518)
         );
  FADDX1_LVT U1145 ( .A(n1528), .B(n1539), .CI(n1537), .CO(n1519), .S(n1520)
         );
  FADDX1_LVT U1146 ( .A(n1541), .B(n1530), .CI(n1526), .CO(n1521), .S(n1522)
         );
  FADDX1_LVT U1147 ( .A(n2032), .B(n1545), .CI(n1543), .CO(n1523), .S(n1524)
         );
  FADDX1_LVT U1148 ( .A(n2096), .B(n1904), .CI(n1968), .CO(n1525), .S(n1526)
         );
  FADDX1_LVT U1149 ( .A(n2160), .B(n1776), .CI(n1840), .CO(n1527), .S(n1528)
         );
  FADDX1_LVT U1150 ( .A(I3[12]), .B(n1712), .CI(n2224), .CO(n1529), .S(n1530)
         );
  FADDX1_LVT U1151 ( .A(n1536), .B(n1549), .CI(n1534), .CO(n1531), .S(n1532)
         );
  FADDX1_LVT U1152 ( .A(n1540), .B(n1538), .CI(n1551), .CO(n1533), .S(n1534)
         );
  FADDX1_LVT U1153 ( .A(n1544), .B(n1555), .CI(n1553), .CO(n1535), .S(n1536)
         );
  FADDX1_LVT U1154 ( .A(n1557), .B(n1546), .CI(n1542), .CO(n1537), .S(n1538)
         );
  FADDX1_LVT U1155 ( .A(n2033), .B(n1561), .CI(n1559), .CO(n1539), .S(n1540)
         );
  FADDX1_LVT U1156 ( .A(n2097), .B(n1905), .CI(n1969), .CO(n1541), .S(n1542)
         );
  FADDX1_LVT U1157 ( .A(n2161), .B(n1777), .CI(n1841), .CO(n1543), .S(n1544)
         );
  FADDX1_LVT U1158 ( .A(I3[11]), .B(n1713), .CI(n2225), .CO(n1545), .S(n1546)
         );
  FADDX1_LVT U1159 ( .A(n1565), .B(n1552), .CI(n1550), .CO(n1547), .S(n1548)
         );
  FADDX1_LVT U1160 ( .A(n1556), .B(n1554), .CI(n1567), .CO(n1549), .S(n1550)
         );
  FADDX1_LVT U1161 ( .A(n1560), .B(n1571), .CI(n1569), .CO(n1551), .S(n1552)
         );
  FADDX1_LVT U1162 ( .A(n1573), .B(n1562), .CI(n1558), .CO(n1553), .S(n1554)
         );
  FADDX1_LVT U1163 ( .A(n2034), .B(n1577), .CI(n1575), .CO(n1555), .S(n1556)
         );
  FADDX1_LVT U1164 ( .A(n2098), .B(n1906), .CI(n1970), .CO(n1557), .S(n1558)
         );
  FADDX1_LVT U1165 ( .A(n2162), .B(n1778), .CI(n1842), .CO(n1559), .S(n1560)
         );
  FADDX1_LVT U1166 ( .A(I3[10]), .B(n1714), .CI(n2226), .CO(n1561), .S(n1562)
         );
  FADDX1_LVT U1167 ( .A(n1581), .B(n1568), .CI(n1566), .CO(n1563), .S(n1564)
         );
  FADDX1_LVT U1168 ( .A(n1572), .B(n1583), .CI(n1570), .CO(n1565), .S(n1566)
         );
  FADDX1_LVT U1169 ( .A(n1576), .B(n1587), .CI(n1585), .CO(n1567), .S(n1568)
         );
  FADDX1_LVT U1170 ( .A(n1589), .B(n1578), .CI(n1574), .CO(n1569), .S(n1570)
         );
  FADDX1_LVT U1171 ( .A(n2035), .B(n1593), .CI(n1591), .CO(n1571), .S(n1572)
         );
  FADDX1_LVT U1172 ( .A(n2099), .B(n1907), .CI(n1971), .CO(n1573), .S(n1574)
         );
  FADDX1_LVT U1173 ( .A(n2163), .B(n1779), .CI(n1843), .CO(n1575), .S(n1576)
         );
  FADDX1_LVT U1174 ( .A(I3[9]), .B(n1715), .CI(n2227), .CO(n1577), .S(n1578)
         );
  FADDX1_LVT U1175 ( .A(n1597), .B(n1584), .CI(n1582), .CO(n1579), .S(n1580)
         );
  FADDX1_LVT U1176 ( .A(n1588), .B(n1599), .CI(n1586), .CO(n1581), .S(n1582)
         );
  FADDX1_LVT U1177 ( .A(n1590), .B(n1592), .CI(n1601), .CO(n1583), .S(n1584)
         );
  FADDX1_LVT U1178 ( .A(n1605), .B(n1603), .CI(n1594), .CO(n1585), .S(n1586)
         );
  FADDX1_LVT U1179 ( .A(n2100), .B(n2036), .CI(n1607), .CO(n1587), .S(n1588)
         );
  FADDX1_LVT U1180 ( .A(n2164), .B(n1908), .CI(n1972), .CO(n1589), .S(n1590)
         );
  FADDX1_LVT U1181 ( .A(n2228), .B(n1780), .CI(n1844), .CO(n1591), .S(n1592)
         );
  FADDX1_LVT U1184 ( .A(n1611), .B(n1600), .CI(n1598), .CO(n1595), .S(n1596)
         );
  FADDX1_LVT U1185 ( .A(n1606), .B(n1613), .CI(n1602), .CO(n1597), .S(n1598)
         );
  FADDX1_LVT U1186 ( .A(n1617), .B(n1615), .CI(n1604), .CO(n1599), .S(n1600)
         );
  FADDX1_LVT U1187 ( .A(n2037), .B(n1619), .CI(n1608), .CO(n1601), .S(n1602)
         );
  FADDX1_LVT U1188 ( .A(n1973), .B(n2101), .CI(n1909), .CO(n1603), .S(n1604)
         );
  FADDX1_LVT U1189 ( .A(n2229), .B(n1781), .CI(n2165), .CO(n1605), .S(n1606)
         );
  HADDX1_LVT U1190 ( .A0(I3[7]), .B0(n1845), .C1(n1607), .SO(n1608) );
  FADDX1_LVT U1191 ( .A(n1623), .B(n1614), .CI(n1612), .CO(n1609), .S(n1610)
         );
  FADDX1_LVT U1192 ( .A(n1616), .B(n1618), .CI(n1625), .CO(n1611), .S(n1612)
         );
  FADDX1_LVT U1193 ( .A(n1629), .B(n1620), .CI(n1627), .CO(n1613), .S(n1614)
         );
  FADDX1_LVT U1194 ( .A(n2102), .B(n1974), .CI(n2038), .CO(n1615), .S(n1616)
         );
  FADDX1_LVT U1195 ( .A(n2230), .B(n1846), .CI(n2166), .CO(n1617), .S(n1618)
         );
  HADDX1_LVT U1196 ( .A0(I3[6]), .B0(n1910), .C1(n1619), .SO(n1620) );
  FADDX1_LVT U1197 ( .A(n1633), .B(n1626), .CI(n1624), .CO(n1621), .S(n1622)
         );
  FADDX1_LVT U1198 ( .A(n1630), .B(n1635), .CI(n1628), .CO(n1623), .S(n1624)
         );
  FADDX1_LVT U1199 ( .A(n2103), .B(n2039), .CI(n1637), .CO(n1625), .S(n1626)
         );
  FADDX1_LVT U1200 ( .A(n2231), .B(n1911), .CI(n2167), .CO(n1627), .S(n1628)
         );
  HADDX1_LVT U1201 ( .A0(I3[5]), .B0(n1975), .C1(n1629), .SO(n1630) );
  FADDX1_LVT U1202 ( .A(n1641), .B(n1636), .CI(n1634), .CO(n1631), .S(n1632)
         );
  FADDX1_LVT U1203 ( .A(n2168), .B(n1643), .CI(n1638), .CO(n1633), .S(n1634)
         );
  FADDX1_LVT U1204 ( .A(n2232), .B(n1976), .CI(n2104), .CO(n1635), .S(n1636)
         );
  HADDX1_LVT U1205 ( .A0(I3[4]), .B0(n2040), .C1(n1637), .SO(n1638) );
  FADDX1_LVT U1206 ( .A(n1647), .B(n1644), .CI(n1642), .CO(n1639), .S(n1640)
         );
  FADDX1_LVT U1207 ( .A(n2233), .B(n2041), .CI(n2169), .CO(n1641), .S(n1642)
         );
  HADDX1_LVT U1208 ( .A0(I3[3]), .B0(n2105), .C1(n1643), .SO(n1644) );
  FADDX1_LVT U1209 ( .A(n2170), .B(n2106), .CI(n1649), .CO(n1645), .S(n1646)
         );
  HADDX1_LVT U1210 ( .A0(I3[2]), .B0(n2234), .C1(n1647), .SO(n1648) );
  HADDX1_LVT U1211 ( .A0(I3[1]), .B0(n2235), .C1(n1649), .SO(n1650) );
  AO221X1_LVT U1874 ( .A1(1'b1), .A2(n2547), .A3(n2761), .A4(n2759), .A5(n2758), .Y(n2549) );
  OA221X1_LVT U1875 ( .A1(n2714), .A2(1'b1), .A3(n2714), .A4(n2536), .A5(n2719), .Y(n2537) );
  AO221X1_LVT U1876 ( .A1(1'b1), .A2(n2530), .A3(n2625), .A4(n2619), .A5(n2620), .Y(n2532) );
  OR2X1_LVT U1877 ( .A1(n715), .A2(n700), .Y(n2527) );
  AND3X1_LVT U1878 ( .A1(n2621), .A2(n2623), .A3(n2527), .Y(n2528) );
  AOI22X1_LVT U1879 ( .A1(n715), .A2(n700), .A3(n2528), .A4(n2624), .Y(n2529)
         );
  AND3X1_LVT U1880 ( .A1(n2618), .A2(n2625), .A3(n2617), .Y(n2530) );
  NAND3X0_LVT U1882 ( .A1(n2626), .A2(n2528), .A3(n2532), .Y(n2533) );
  NAND3X0_LVT U1883 ( .A1(n2621), .A2(n2622), .A3(n2527), .Y(n2534) );
  NAND3X0_LVT U1884 ( .A1(n716), .A2(n731), .A3(n2527), .Y(n2535) );
  NAND4X0_LVT U1885 ( .A1(n2529), .A2(n2533), .A3(n2534), .A4(n2535), .Y(n2594) );
  OA221X1_LVT U1886 ( .A1(n2712), .A2(n2716), .A3(n2712), .A4(n2717), .A5(
        n2718), .Y(n2536) );
  OA22X1_LVT U1887 ( .A1(n1243), .A2(n1228), .A3(n2537), .A4(n2713), .Y(n2538)
         );
  OA22X1_LVT U1888 ( .A1(n2538), .A2(n2715), .A3(n1227), .A4(n1212), .Y(n2539)
         );
  AO21X1_LVT U1889 ( .A1(n1212), .A2(n1227), .A3(n2539), .Y(n2618) );
  OA221X1_LVT U1890 ( .A1(I3[0]), .A2(I2[0]), .A3(I3[0]), .A4(I1[0]), .A5(
        n2589), .Y(O1[0]) );
  AO222X1_LVT U1891 ( .A1(n1631), .A2(n1622), .A3(n1631), .A4(n2782), .A5(
        n1622), .A6(n2782), .Y(n2776) );
  AO21X1_LVT U1893 ( .A1(n2778), .A2(n2779), .A3(n2776), .Y(n2541) );
  OA22X1_LVT U1894 ( .A1(n1621), .A2(n1610), .A3(n1609), .A4(n1596), .Y(n2542)
         );
  OR2X1_LVT U1895 ( .A1(n1609), .A2(n1596), .Y(n2543) );
  AO222X1_LVT U1896 ( .A1(n2541), .A2(n2542), .A3(n2543), .A4(n2777), .A5(
        n1596), .A6(n1609), .Y(n2757) );
  OR2X1_LVT U1897 ( .A1(n1340), .A2(n2739), .Y(n2544) );
  AO22X1_LVT U1898 ( .A1(n2735), .A2(n2736), .A3(n2738), .A4(n2737), .Y(n2545)
         );
  AO221X1_LVT U1899 ( .A1(n2544), .A2(n1355), .A3(n2739), .A4(n1340), .A5(
        n2545), .Y(n2712) );
  AO21X1_LVT U1900 ( .A1(n2784), .A2(n551), .A3(n2785), .Y(n2546) );
  AO222X1_LVT U1901 ( .A1(n1645), .A2(n1640), .A3(n1645), .A4(n2546), .A5(
        n1640), .A6(n2546), .Y(n2778) );
  AND3X1_LVT U1902 ( .A1(n2757), .A2(n2761), .A3(n2756), .Y(n2547) );
  OA22X1_LVT U1904 ( .A1(n1499), .A2(n1484), .A3(n1483), .A4(n1468), .Y(n2550)
         );
  OR2X1_LVT U1905 ( .A1(n1483), .A2(n1468), .Y(n2551) );
  AO222X1_LVT U1906 ( .A1(n2549), .A2(n2550), .A3(n2551), .A4(n2760), .A5(
        n1468), .A6(n1483), .Y(n2716) );
  AO222X1_LVT U1907 ( .A1(n683), .A2(n670), .A3(n683), .A4(n2615), .A5(n670), 
        .A6(n2615), .Y(n2608) );
  OR2X1_LVT U1908 ( .A1(n828), .A2(n2647), .Y(n2552) );
  AO22X1_LVT U1909 ( .A1(n2643), .A2(n2644), .A3(n2646), .A4(n2645), .Y(n2553)
         );
  AO221X1_LVT U1910 ( .A1(n2552), .A2(n843), .A3(n2647), .A4(n828), .A5(n2553), 
        .Y(n2620) );
  AO22X1_LVT U1911 ( .A1(n2691), .A2(n2692), .A3(n2694), .A4(n2693), .Y(n2554)
         );
  OR2X1_LVT U1912 ( .A1(n1084), .A2(n2695), .Y(n2555) );
  AO221X1_LVT U1913 ( .A1(n2555), .A2(n1099), .A3(n2695), .A4(n1084), .A5(
        n2554), .Y(n2667) );
  AO222X1_LVT U1914 ( .A1(n1259), .A2(n1244), .A3(n1259), .A4(n2723), .A5(
        n1244), .A6(n2723), .Y(n2713) );
  AO222X1_LVT U1915 ( .A1(n1451), .A2(n1436), .A3(n1451), .A4(n2754), .A5(
        n1436), .A6(n2754), .Y(n2750) );
  AO222X1_LVT U1916 ( .A1(n1515), .A2(n1500), .A3(n1515), .A4(n2765), .A5(
        n1500), .A6(n2765), .Y(n2758) );
  AO222X1_LVT U1917 ( .A1(n1579), .A2(n1564), .A3(n1579), .A4(n2774), .A5(
        n1564), .A6(n2774), .Y(n2770) );
  AO222X1_LVT U1918 ( .A1(n747), .A2(n732), .A3(n747), .A4(n2630), .A5(n732), 
        .A6(n2630), .Y(n2622) );
  AO222X1_LVT U1919 ( .A1(n811), .A2(n796), .A3(n811), .A4(n2640), .A5(n796), 
        .A6(n2640), .Y(n2636) );
  AO222X1_LVT U1920 ( .A1(n875), .A2(n860), .A3(n875), .A4(n2653), .A5(n860), 
        .A6(n2653), .Y(n2644) );
  AO222X1_LVT U1921 ( .A1(n939), .A2(n924), .A3(n939), .A4(n2662), .A5(n924), 
        .A6(n2662), .Y(n2658) );
  AO222X1_LVT U1922 ( .A1(n1003), .A2(n988), .A3(n1003), .A4(n2679), .A5(n988), 
        .A6(n2679), .Y(n2672) );
  AO222X1_LVT U1923 ( .A1(n1067), .A2(n1052), .A3(n1067), .A4(n2689), .A5(
        n1052), .A6(n2689), .Y(n2685) );
  AO222X1_LVT U1924 ( .A1(n1131), .A2(n1116), .A3(n1131), .A4(n2701), .A5(
        n1116), .A6(n2701), .Y(n2692) );
  AO222X1_LVT U1925 ( .A1(n1195), .A2(n1180), .A3(n1195), .A4(n2710), .A5(
        n1180), .A6(n2710), .Y(n2706) );
  AO222X1_LVT U1926 ( .A1(n1323), .A2(n1308), .A3(n1323), .A4(n2733), .A5(
        n1308), .A6(n2733), .Y(n2729) );
  AO222X1_LVT U1927 ( .A1(n1387), .A2(n1372), .A3(n1387), .A4(n2745), .A5(
        n1372), .A6(n2745), .Y(n2736) );
  AO222X1_LVT U1928 ( .A1(n639), .A2(n634), .A3(n647), .A4(n640), .A5(n2602), 
        .A6(n2601), .Y(n2556) );
  AND2X1_LVT U1929 ( .A1(n2603), .A2(n2556), .Y(n2598) );
  NBUFFX2_LVT U1930 ( .A(I2[14]), .Y(n2563) );
  NBUFFX2_LVT U1931 ( .A(I2[6]), .Y(n2558) );
  NBUFFX2_LVT U1932 ( .A(I2[61]), .Y(n2582) );
  NBUFFX2_LVT U1933 ( .A(I2[46]), .Y(n2574) );
  NBUFFX2_LVT U1934 ( .A(I2[38]), .Y(n2571) );
  NBUFFX2_LVT U1935 ( .A(I2[54]), .Y(n2577) );
  NBUFFX2_LVT U1936 ( .A(I2[22]), .Y(n2565) );
  NBUFFX2_LVT U1937 ( .A(I2[63]), .Y(n2583) );
  NBUFFX2_LVT U1938 ( .A(I2[60]), .Y(n2581) );
  NBUFFX2_LVT U1939 ( .A(I2[57]), .Y(n2580) );
  NBUFFX2_LVT U1940 ( .A(I2[56]), .Y(n2579) );
  NBUFFX2_LVT U1941 ( .A(I2[55]), .Y(n2578) );
  NBUFFX2_LVT U1942 ( .A(I2[52]), .Y(n2575) );
  NBUFFX2_LVT U1943 ( .A(I2[53]), .Y(n2576) );
  NBUFFX2_LVT U1944 ( .A(I2[44]), .Y(n2572) );
  NBUFFX2_LVT U1945 ( .A(I2[45]), .Y(n2573) );
  NBUFFX2_LVT U1946 ( .A(I2[9]), .Y(n2560) );
  NBUFFX2_LVT U1947 ( .A(I2[12]), .Y(n2561) );
  NBUFFX2_LVT U1948 ( .A(I2[13]), .Y(n2562) );
  NBUFFX2_LVT U1949 ( .A(I2[20]), .Y(n2564) );
  NBUFFX2_LVT U1950 ( .A(I2[37]), .Y(n2570) );
  NBUFFX2_LVT U1951 ( .A(I2[28]), .Y(n2566) );
  NBUFFX2_LVT U1952 ( .A(I2[31]), .Y(n2568) );
  NBUFFX2_LVT U1953 ( .A(I2[30]), .Y(n2567) );
  NBUFFX2_LVT U1954 ( .A(I2[36]), .Y(n2569) );
  NBUFFX2_LVT U1955 ( .A(I2[7]), .Y(n2559) );
  NBUFFX2_LVT U1956 ( .A(I2[4]), .Y(n2557) );
  NBUFFX2_LVT U1957 ( .A(I1[5]), .Y(n2584) );
  NBUFFX2_LVT U1958 ( .A(I1[7]), .Y(n2585) );
  INVX1_LVT U1959 ( .A(n2589), .Y(n2586) );
  INVX1_LVT U1960 ( .A(I3[64]), .Y(n2587) );
  INVX1_LVT U1961 ( .A(I3[8]), .Y(n2588) );
  FADDX1_LVT U1962 ( .A(n2590), .B(n627), .CI(n2591), .S(O1[72]) );
  AND2X1_LVT U1963 ( .A1(I1[8]), .A2(I2[64]), .Y(n2591) );
  OA222X1_LVT U1964 ( .A1(n2592), .A2(n2593), .A3(n2592), .A4(n2594), .A5(
        n2592), .A6(n2595), .Y(n2590) );
  AO22X1_LVT U1965 ( .A1(n2596), .A2(n2595), .A3(n628), .A4(n629), .Y(n2592)
         );
  OR2X1_LVT U1966 ( .A1(n628), .A2(n629), .Y(n2595) );
  FADDX1_LVT U1967 ( .A(n2597), .B(n628), .CI(n629), .S(O1[71]) );
  AO21X1_LVT U1968 ( .A1(n2594), .A2(n2593), .A3(n2596), .Y(n2597) );
  AO222X1_LVT U1969 ( .A1(n630), .A2(n633), .A3(n630), .A4(n2598), .A5(n633), 
        .A6(n2598), .Y(n2596) );
  OA21X1_LVT U1970 ( .A1(n630), .A2(n633), .A3(n2599), .Y(n2593) );
  FADDX1_LVT U1971 ( .A(n2600), .B(n630), .CI(n633), .S(O1[70]) );
  AO21X1_LVT U1972 ( .A1(n2599), .A2(n2594), .A3(n2598), .Y(n2600) );
  AND3X1_LVT U1973 ( .A1(n2604), .A2(n2602), .A3(n2603), .Y(n2599) );
  OR2X1_LVT U1974 ( .A1(n639), .A2(n634), .Y(n2603) );
  FADDX1_LVT U1975 ( .A(n639), .B(n634), .CI(n2605), .S(O1[69]) );
  AO22X1_LVT U1976 ( .A1(n647), .A2(n640), .A3(n2606), .A4(n2602), .Y(n2605)
         );
  OR2X1_LVT U1977 ( .A1(n647), .A2(n640), .Y(n2602) );
  FADDX1_LVT U1978 ( .A(n647), .B(n640), .CI(n2606), .S(O1[68]) );
  AO21X1_LVT U1979 ( .A1(n2594), .A2(n2604), .A3(n2601), .Y(n2606) );
  AO221X1_LVT U1980 ( .A1(n657), .A2(n648), .A3(n2607), .A4(n2608), .A5(n2609), 
        .Y(n2601) );
  AND3X1_LVT U1981 ( .A1(n669), .A2(n658), .A3(n2610), .Y(n2609) );
  OA21X1_LVT U1982 ( .A1(n648), .A2(n657), .A3(n2611), .Y(n2607) );
  AND3X1_LVT U1983 ( .A1(n2612), .A2(n2611), .A3(n2610), .Y(n2604) );
  OR2X1_LVT U1984 ( .A1(n657), .A2(n648), .Y(n2610) );
  FADDX1_LVT U1985 ( .A(n657), .B(n648), .CI(n2613), .S(O1[67]) );
  AO22X1_LVT U1986 ( .A1(n669), .A2(n658), .A3(n2614), .A4(n2611), .Y(n2613)
         );
  OR2X1_LVT U1987 ( .A1(n669), .A2(n658), .Y(n2611) );
  FADDX1_LVT U1988 ( .A(n669), .B(n658), .CI(n2614), .S(O1[66]) );
  AO21X1_LVT U1989 ( .A1(n2612), .A2(n2594), .A3(n2608), .Y(n2614) );
  OA22X1_LVT U1990 ( .A1(n683), .A2(n670), .A3(n699), .A4(n684), .Y(n2612) );
  FADDX1_LVT U1991 ( .A(n683), .B(n670), .CI(n2616), .S(O1[65]) );
  OA22X1_LVT U1992 ( .A1(n699), .A2(n684), .A3(n2615), .A4(n2594), .Y(n2616)
         );
  AND2X1_LVT U1993 ( .A1(n699), .A2(n684), .Y(n2615) );
  FADDX1_LVT U1994 ( .A(n699), .B(n684), .CI(n2594), .S(O1[64]) );
  FADDX1_LVT U1995 ( .A(n715), .B(n700), .CI(n2627), .S(O1[63]) );
  AO22X1_LVT U1996 ( .A1(n731), .A2(n716), .A3(n2628), .A4(n2621), .Y(n2627)
         );
  OR2X1_LVT U1997 ( .A1(n731), .A2(n716), .Y(n2621) );
  FADDX1_LVT U1998 ( .A(n731), .B(n716), .CI(n2628), .S(O1[62]) );
  AO21X1_LVT U1999 ( .A1(n2623), .A2(n2629), .A3(n2622), .Y(n2628) );
  OA22X1_LVT U2000 ( .A1(n747), .A2(n732), .A3(n763), .A4(n748), .Y(n2623) );
  FADDX1_LVT U2001 ( .A(n747), .B(n732), .CI(n2631), .S(O1[61]) );
  AO221X1_LVT U2002 ( .A1(n2629), .A2(n763), .A3(n2629), .A4(n748), .A5(n2630), 
        .Y(n2631) );
  AND2X1_LVT U2003 ( .A1(n763), .A2(n748), .Y(n2630) );
  FADDX1_LVT U2004 ( .A(n763), .B(n748), .CI(n2629), .S(O1[60]) );
  AO21X1_LVT U2005 ( .A1(n2626), .A2(n2632), .A3(n2624), .Y(n2629) );
  AO222X1_LVT U2006 ( .A1(n779), .A2(n764), .A3(n2633), .A4(n2634), .A5(n2635), 
        .A6(n2636), .Y(n2624) );
  OR2X1_LVT U2007 ( .A1(n764), .A2(n779), .Y(n2634) );
  AND2X1_LVT U2008 ( .A1(n2635), .A2(n2637), .Y(n2626) );
  OA22X1_LVT U2009 ( .A1(n779), .A2(n764), .A3(n795), .A4(n780), .Y(n2635) );
  FADDX1_LVT U2010 ( .A(n779), .B(n764), .CI(n2638), .S(O1[59]) );
  OA22X1_LVT U2011 ( .A1(n2633), .A2(n2639), .A3(n795), .A4(n780), .Y(n2638)
         );
  AND2X1_LVT U2012 ( .A1(n795), .A2(n780), .Y(n2633) );
  FADDX1_LVT U2013 ( .A(n795), .B(n780), .CI(n2639), .S(O1[58]) );
  AO21X1_LVT U2014 ( .A1(n2637), .A2(n2632), .A3(n2636), .Y(n2639) );
  OA22X1_LVT U2015 ( .A1(n811), .A2(n796), .A3(n827), .A4(n812), .Y(n2637) );
  FADDX1_LVT U2016 ( .A(n811), .B(n796), .CI(n2641), .S(O1[57]) );
  OA22X1_LVT U2017 ( .A1(n2640), .A2(n2632), .A3(n827), .A4(n812), .Y(n2641)
         );
  AND2X1_LVT U2018 ( .A1(n827), .A2(n812), .Y(n2640) );
  FADDX1_LVT U2019 ( .A(n827), .B(n812), .CI(n2632), .S(O1[56]) );
  AO21X1_LVT U2020 ( .A1(n2625), .A2(n2642), .A3(n2620), .Y(n2632) );
  AND2X1_LVT U2021 ( .A1(n2646), .A2(n2648), .Y(n2625) );
  AND2X1_LVT U2022 ( .A1(n2643), .A2(n2649), .Y(n2646) );
  OA22X1_LVT U2023 ( .A1(n843), .A2(n828), .A3(n859), .A4(n844), .Y(n2643) );
  FADDX1_LVT U2024 ( .A(n843), .B(n828), .CI(n2650), .S(O1[55]) );
  OA22X1_LVT U2025 ( .A1(n2647), .A2(n2651), .A3(n859), .A4(n844), .Y(n2650)
         );
  AND2X1_LVT U2026 ( .A1(n859), .A2(n844), .Y(n2647) );
  FADDX1_LVT U2027 ( .A(n859), .B(n844), .CI(n2651), .S(O1[54]) );
  AO21X1_LVT U2028 ( .A1(n2649), .A2(n2652), .A3(n2644), .Y(n2651) );
  OA22X1_LVT U2029 ( .A1(n875), .A2(n860), .A3(n891), .A4(n876), .Y(n2649) );
  FADDX1_LVT U2030 ( .A(n875), .B(n860), .CI(n2654), .S(O1[53]) );
  OA22X1_LVT U2031 ( .A1(n2653), .A2(n2652), .A3(n891), .A4(n876), .Y(n2654)
         );
  AND2X1_LVT U2032 ( .A1(n891), .A2(n876), .Y(n2653) );
  FADDX1_LVT U2033 ( .A(n891), .B(n876), .CI(n2652), .S(O1[52]) );
  AO21X1_LVT U2034 ( .A1(n2648), .A2(n2642), .A3(n2645), .Y(n2652) );
  AO222X1_LVT U2035 ( .A1(n907), .A2(n892), .A3(n2655), .A4(n2656), .A5(n2657), 
        .A6(n2658), .Y(n2645) );
  OR2X1_LVT U2036 ( .A1(n892), .A2(n907), .Y(n2656) );
  AND2X1_LVT U2037 ( .A1(n2657), .A2(n2659), .Y(n2648) );
  OA22X1_LVT U2038 ( .A1(n907), .A2(n892), .A3(n923), .A4(n908), .Y(n2657) );
  FADDX1_LVT U2039 ( .A(n907), .B(n892), .CI(n2660), .S(O1[51]) );
  OA22X1_LVT U2040 ( .A1(n2655), .A2(n2661), .A3(n923), .A4(n908), .Y(n2660)
         );
  AND2X1_LVT U2041 ( .A1(n923), .A2(n908), .Y(n2655) );
  FADDX1_LVT U2042 ( .A(n923), .B(n908), .CI(n2661), .S(O1[50]) );
  AO21X1_LVT U2043 ( .A1(n2659), .A2(n2642), .A3(n2658), .Y(n2661) );
  OA22X1_LVT U2044 ( .A1(n939), .A2(n924), .A3(n955), .A4(n940), .Y(n2659) );
  FADDX1_LVT U2045 ( .A(n939), .B(n924), .CI(n2663), .S(O1[49]) );
  OA22X1_LVT U2046 ( .A1(n2662), .A2(n2642), .A3(n955), .A4(n940), .Y(n2663)
         );
  AND2X1_LVT U2047 ( .A1(n955), .A2(n940), .Y(n2662) );
  FADDX1_LVT U2048 ( .A(n955), .B(n940), .CI(n2642), .S(O1[48]) );
  AO21X1_LVT U2049 ( .A1(n2617), .A2(n2618), .A3(n2619), .Y(n2642) );
  AO221X1_LVT U2050 ( .A1(n2664), .A2(n2665), .A3(n2666), .A4(n2667), .A5(
        n2668), .Y(n2619) );
  AO222X1_LVT U2051 ( .A1(n971), .A2(n956), .A3(n2669), .A4(n2670), .A5(n2671), 
        .A6(n2672), .Y(n2668) );
  OR2X1_LVT U2052 ( .A1(n956), .A2(n971), .Y(n2670) );
  AND2X1_LVT U2053 ( .A1(n2666), .A2(n2673), .Y(n2617) );
  AND2X1_LVT U2054 ( .A1(n2674), .A2(n2665), .Y(n2666) );
  AND2X1_LVT U2055 ( .A1(n2671), .A2(n2675), .Y(n2665) );
  OA22X1_LVT U2056 ( .A1(n971), .A2(n956), .A3(n987), .A4(n972), .Y(n2671) );
  FADDX1_LVT U2057 ( .A(n971), .B(n956), .CI(n2676), .S(O1[47]) );
  OA22X1_LVT U2058 ( .A1(n2669), .A2(n2677), .A3(n987), .A4(n972), .Y(n2676)
         );
  AND2X1_LVT U2059 ( .A1(n987), .A2(n972), .Y(n2669) );
  FADDX1_LVT U2060 ( .A(n987), .B(n972), .CI(n2677), .S(O1[46]) );
  AO21X1_LVT U2061 ( .A1(n2675), .A2(n2678), .A3(n2672), .Y(n2677) );
  OA22X1_LVT U2062 ( .A1(n1003), .A2(n988), .A3(n1019), .A4(n1004), .Y(n2675)
         );
  FADDX1_LVT U2063 ( .A(n1003), .B(n988), .CI(n2680), .S(O1[45]) );
  OA22X1_LVT U2064 ( .A1(n2679), .A2(n2678), .A3(n1019), .A4(n1004), .Y(n2680)
         );
  AND2X1_LVT U2065 ( .A1(n1019), .A2(n1004), .Y(n2679) );
  FADDX1_LVT U2066 ( .A(n1019), .B(n1004), .CI(n2678), .S(O1[44]) );
  AO21X1_LVT U2067 ( .A1(n2674), .A2(n2681), .A3(n2664), .Y(n2678) );
  AO222X1_LVT U2068 ( .A1(n1035), .A2(n1020), .A3(n2682), .A4(n2683), .A5(
        n2684), .A6(n2685), .Y(n2664) );
  OR2X1_LVT U2069 ( .A1(n1020), .A2(n1035), .Y(n2683) );
  AND2X1_LVT U2070 ( .A1(n2684), .A2(n2686), .Y(n2674) );
  OA22X1_LVT U2071 ( .A1(n1035), .A2(n1020), .A3(n1051), .A4(n1036), .Y(n2684)
         );
  FADDX1_LVT U2072 ( .A(n1035), .B(n1020), .CI(n2687), .S(O1[43]) );
  OA22X1_LVT U2073 ( .A1(n2682), .A2(n2688), .A3(n1051), .A4(n1036), .Y(n2687)
         );
  AND2X1_LVT U2074 ( .A1(n1051), .A2(n1036), .Y(n2682) );
  FADDX1_LVT U2075 ( .A(n1051), .B(n1036), .CI(n2688), .S(O1[42]) );
  AO21X1_LVT U2076 ( .A1(n2686), .A2(n2681), .A3(n2685), .Y(n2688) );
  OA22X1_LVT U2077 ( .A1(n1067), .A2(n1052), .A3(n1083), .A4(n1068), .Y(n2686)
         );
  FADDX1_LVT U2078 ( .A(n1067), .B(n1052), .CI(n2690), .S(O1[41]) );
  OA22X1_LVT U2079 ( .A1(n2689), .A2(n2681), .A3(n1083), .A4(n1068), .Y(n2690)
         );
  AND2X1_LVT U2080 ( .A1(n1083), .A2(n1068), .Y(n2689) );
  FADDX1_LVT U2081 ( .A(n1083), .B(n1068), .CI(n2681), .S(O1[40]) );
  AO21X1_LVT U2082 ( .A1(n2673), .A2(n2618), .A3(n2667), .Y(n2681) );
  AND2X1_LVT U2083 ( .A1(n2694), .A2(n2696), .Y(n2673) );
  AND2X1_LVT U2084 ( .A1(n2691), .A2(n2697), .Y(n2694) );
  OA22X1_LVT U2085 ( .A1(n1099), .A2(n1084), .A3(n1115), .A4(n1100), .Y(n2691)
         );
  FADDX1_LVT U2086 ( .A(n1099), .B(n1084), .CI(n2698), .S(O1[39]) );
  OA22X1_LVT U2087 ( .A1(n2695), .A2(n2699), .A3(n1115), .A4(n1100), .Y(n2698)
         );
  AND2X1_LVT U2088 ( .A1(n1115), .A2(n1100), .Y(n2695) );
  FADDX1_LVT U2089 ( .A(n1115), .B(n1100), .CI(n2699), .S(O1[38]) );
  AO21X1_LVT U2090 ( .A1(n2697), .A2(n2700), .A3(n2692), .Y(n2699) );
  OA22X1_LVT U2091 ( .A1(n1131), .A2(n1116), .A3(n1147), .A4(n1132), .Y(n2697)
         );
  FADDX1_LVT U2092 ( .A(n1131), .B(n1116), .CI(n2702), .S(O1[37]) );
  OA22X1_LVT U2093 ( .A1(n2701), .A2(n2700), .A3(n1147), .A4(n1132), .Y(n2702)
         );
  AND2X1_LVT U2094 ( .A1(n1147), .A2(n1132), .Y(n2701) );
  FADDX1_LVT U2095 ( .A(n1147), .B(n1132), .CI(n2700), .S(O1[36]) );
  AO21X1_LVT U2096 ( .A1(n2696), .A2(n2618), .A3(n2693), .Y(n2700) );
  AO222X1_LVT U2097 ( .A1(n1163), .A2(n1148), .A3(n2703), .A4(n2704), .A5(
        n2705), .A6(n2706), .Y(n2693) );
  OR2X1_LVT U2098 ( .A1(n1148), .A2(n1163), .Y(n2704) );
  AND2X1_LVT U2099 ( .A1(n2705), .A2(n2707), .Y(n2696) );
  OA22X1_LVT U2100 ( .A1(n1163), .A2(n1148), .A3(n1179), .A4(n1164), .Y(n2705)
         );
  FADDX1_LVT U2101 ( .A(n1163), .B(n1148), .CI(n2708), .S(O1[35]) );
  OA22X1_LVT U2102 ( .A1(n2703), .A2(n2709), .A3(n1179), .A4(n1164), .Y(n2708)
         );
  AND2X1_LVT U2103 ( .A1(n1179), .A2(n1164), .Y(n2703) );
  FADDX1_LVT U2104 ( .A(n1179), .B(n1164), .CI(n2709), .S(O1[34]) );
  AO21X1_LVT U2105 ( .A1(n2707), .A2(n2618), .A3(n2706), .Y(n2709) );
  OA22X1_LVT U2106 ( .A1(n1195), .A2(n1180), .A3(n1211), .A4(n1196), .Y(n2707)
         );
  FADDX1_LVT U2107 ( .A(n1195), .B(n1180), .CI(n2711), .S(O1[33]) );
  AO221X1_LVT U2108 ( .A1(n2618), .A2(n1211), .A3(n2618), .A4(n1196), .A5(
        n2710), .Y(n2711) );
  AND2X1_LVT U2109 ( .A1(n1211), .A2(n1196), .Y(n2710) );
  FADDX1_LVT U2110 ( .A(n1211), .B(n1196), .CI(n2618), .S(O1[32]) );
  FADDX1_LVT U2111 ( .A(n1227), .B(n1212), .CI(n2720), .S(O1[31]) );
  AO221X1_LVT U2112 ( .A1(n2721), .A2(n1243), .A3(n2721), .A4(n1228), .A5(
        n2715), .Y(n2720) );
  AND2X1_LVT U2113 ( .A1(n1243), .A2(n1228), .Y(n2715) );
  FADDX1_LVT U2114 ( .A(n1243), .B(n1228), .CI(n2721), .S(O1[30]) );
  AO21X1_LVT U2115 ( .A1(n2719), .A2(n2722), .A3(n2713), .Y(n2721) );
  OA22X1_LVT U2116 ( .A1(n1259), .A2(n1244), .A3(n1275), .A4(n1260), .Y(n2719)
         );
  FADDX1_LVT U2117 ( .A(n1259), .B(n1244), .CI(n2724), .S(O1[29]) );
  AO221X1_LVT U2118 ( .A1(n2722), .A2(n1275), .A3(n2722), .A4(n1260), .A5(
        n2723), .Y(n2724) );
  AND2X1_LVT U2119 ( .A1(n1275), .A2(n1260), .Y(n2723) );
  FADDX1_LVT U2120 ( .A(n1275), .B(n1260), .CI(n2722), .S(O1[28]) );
  AO21X1_LVT U2121 ( .A1(n2718), .A2(n2725), .A3(n2714), .Y(n2722) );
  AO222X1_LVT U2122 ( .A1(n1291), .A2(n1276), .A3(n2726), .A4(n2727), .A5(
        n2728), .A6(n2729), .Y(n2714) );
  OR2X1_LVT U2123 ( .A1(n1276), .A2(n1291), .Y(n2727) );
  AND2X1_LVT U2124 ( .A1(n2728), .A2(n2730), .Y(n2718) );
  OA22X1_LVT U2125 ( .A1(n1291), .A2(n1276), .A3(n1307), .A4(n1292), .Y(n2728)
         );
  FADDX1_LVT U2126 ( .A(n1291), .B(n1276), .CI(n2731), .S(O1[27]) );
  AO221X1_LVT U2127 ( .A1(n2732), .A2(n1307), .A3(n2732), .A4(n1292), .A5(
        n2726), .Y(n2731) );
  AND2X1_LVT U2128 ( .A1(n1307), .A2(n1292), .Y(n2726) );
  FADDX1_LVT U2129 ( .A(n1307), .B(n1292), .CI(n2732), .S(O1[26]) );
  AO21X1_LVT U2130 ( .A1(n2730), .A2(n2725), .A3(n2729), .Y(n2732) );
  OA22X1_LVT U2131 ( .A1(n1323), .A2(n1308), .A3(n1339), .A4(n1324), .Y(n2730)
         );
  FADDX1_LVT U2132 ( .A(n1323), .B(n1308), .CI(n2734), .S(O1[25]) );
  AO221X1_LVT U2133 ( .A1(n2725), .A2(n1339), .A3(n2725), .A4(n1324), .A5(
        n2733), .Y(n2734) );
  AND2X1_LVT U2134 ( .A1(n1339), .A2(n1324), .Y(n2733) );
  FADDX1_LVT U2135 ( .A(n1339), .B(n1324), .CI(n2725), .S(O1[24]) );
  AO21X1_LVT U2136 ( .A1(n2717), .A2(n2716), .A3(n2712), .Y(n2725) );
  AND2X1_LVT U2137 ( .A1(n2740), .A2(n2738), .Y(n2717) );
  AND2X1_LVT U2138 ( .A1(n2735), .A2(n2741), .Y(n2738) );
  OA22X1_LVT U2139 ( .A1(n1355), .A2(n1340), .A3(n1371), .A4(n1356), .Y(n2735)
         );
  FADDX1_LVT U2140 ( .A(n1355), .B(n1340), .CI(n2742), .S(O1[23]) );
  AO221X1_LVT U2141 ( .A1(n2743), .A2(n1371), .A3(n2743), .A4(n1356), .A5(
        n2739), .Y(n2742) );
  AND2X1_LVT U2142 ( .A1(n1371), .A2(n1356), .Y(n2739) );
  FADDX1_LVT U2143 ( .A(n1371), .B(n1356), .CI(n2743), .S(O1[22]) );
  AO21X1_LVT U2144 ( .A1(n2741), .A2(n2744), .A3(n2736), .Y(n2743) );
  OA22X1_LVT U2145 ( .A1(n1387), .A2(n1372), .A3(n1403), .A4(n1388), .Y(n2741)
         );
  FADDX1_LVT U2146 ( .A(n1387), .B(n1372), .CI(n2746), .S(O1[21]) );
  AO221X1_LVT U2147 ( .A1(n2744), .A2(n1403), .A3(n2744), .A4(n1388), .A5(
        n2745), .Y(n2746) );
  AND2X1_LVT U2148 ( .A1(n1403), .A2(n1388), .Y(n2745) );
  FADDX1_LVT U2149 ( .A(n1403), .B(n1388), .CI(n2744), .S(O1[20]) );
  AO21X1_LVT U2150 ( .A1(n2716), .A2(n2740), .A3(n2737), .Y(n2744) );
  AO222X1_LVT U2151 ( .A1(n1419), .A2(n1404), .A3(n2747), .A4(n2748), .A5(
        n2749), .A6(n2750), .Y(n2737) );
  OR2X1_LVT U2152 ( .A1(n1404), .A2(n1419), .Y(n2748) );
  AND2X1_LVT U2153 ( .A1(n2749), .A2(n2751), .Y(n2740) );
  OA22X1_LVT U2154 ( .A1(n1419), .A2(n1404), .A3(n1435), .A4(n1420), .Y(n2749)
         );
  FADDX1_LVT U2155 ( .A(n1419), .B(n1404), .CI(n2752), .S(O1[19]) );
  AO221X1_LVT U2156 ( .A1(n2753), .A2(n1435), .A3(n2753), .A4(n1420), .A5(
        n2747), .Y(n2752) );
  AND2X1_LVT U2157 ( .A1(n1435), .A2(n1420), .Y(n2747) );
  FADDX1_LVT U2158 ( .A(n1435), .B(n1420), .CI(n2753), .S(O1[18]) );
  AO21X1_LVT U2159 ( .A1(n2751), .A2(n2716), .A3(n2750), .Y(n2753) );
  OA22X1_LVT U2160 ( .A1(n1451), .A2(n1436), .A3(n1467), .A4(n1452), .Y(n2751)
         );
  FADDX1_LVT U2161 ( .A(n1451), .B(n1436), .CI(n2755), .S(O1[17]) );
  OA22X1_LVT U2162 ( .A1(n2716), .A2(n2754), .A3(n1467), .A4(n1452), .Y(n2755)
         );
  AND2X1_LVT U2163 ( .A1(n1467), .A2(n1452), .Y(n2754) );
  FADDX1_LVT U2164 ( .A(n2716), .B(n1467), .CI(n1452), .S(O1[16]) );
  FADDX1_LVT U2165 ( .A(n1483), .B(n1468), .CI(n2762), .S(O1[15]) );
  OA22X1_LVT U2166 ( .A1(n2760), .A2(n2763), .A3(n1499), .A4(n1484), .Y(n2762)
         );
  AND2X1_LVT U2167 ( .A1(n1499), .A2(n1484), .Y(n2760) );
  FADDX1_LVT U2168 ( .A(n1499), .B(n1484), .CI(n2763), .S(O1[14]) );
  AO21X1_LVT U2169 ( .A1(n2761), .A2(n2764), .A3(n2758), .Y(n2763) );
  OA22X1_LVT U2170 ( .A1(n1515), .A2(n1500), .A3(n1531), .A4(n1516), .Y(n2761)
         );
  FADDX1_LVT U2171 ( .A(n1515), .B(n1500), .CI(n2766), .S(O1[13]) );
  OA22X1_LVT U2172 ( .A1(n2765), .A2(n2764), .A3(n1531), .A4(n1516), .Y(n2766)
         );
  AND2X1_LVT U2173 ( .A1(n1531), .A2(n1516), .Y(n2765) );
  FADDX1_LVT U2174 ( .A(n1531), .B(n1516), .CI(n2764), .S(O1[12]) );
  AO21X1_LVT U2175 ( .A1(n2756), .A2(n2757), .A3(n2759), .Y(n2764) );
  AO222X1_LVT U2176 ( .A1(n1547), .A2(n1532), .A3(n2767), .A4(n2768), .A5(
        n2769), .A6(n2770), .Y(n2759) );
  OR2X1_LVT U2177 ( .A1(n1532), .A2(n1547), .Y(n2768) );
  AND2X1_LVT U2178 ( .A1(n2769), .A2(n2771), .Y(n2756) );
  OA22X1_LVT U2179 ( .A1(n1547), .A2(n1532), .A3(n1548), .A4(n1563), .Y(n2769)
         );
  FADDX1_LVT U2180 ( .A(n1547), .B(n1532), .CI(n2772), .S(O1[11]) );
  OA22X1_LVT U2181 ( .A1(n2767), .A2(n2773), .A3(n1548), .A4(n1563), .Y(n2772)
         );
  AND2X1_LVT U2182 ( .A1(n1548), .A2(n1563), .Y(n2767) );
  FADDX1_LVT U2183 ( .A(n1548), .B(n1563), .CI(n2773), .S(O1[10]) );
  AO21X1_LVT U2184 ( .A1(n2771), .A2(n2757), .A3(n2770), .Y(n2773) );
  OA22X1_LVT U2185 ( .A1(n1579), .A2(n1564), .A3(n1580), .A4(n1595), .Y(n2771)
         );
  FADDX1_LVT U2186 ( .A(n1579), .B(n1564), .CI(n2775), .S(O1[9]) );
  AO221X1_LVT U2187 ( .A1(n2757), .A2(n1580), .A3(n2757), .A4(n1595), .A5(
        n2774), .Y(n2775) );
  AND2X1_LVT U2188 ( .A1(n1580), .A2(n1595), .Y(n2774) );
  FADDX1_LVT U2189 ( .A(n1580), .B(n1595), .CI(n2757), .S(O1[8]) );
  FADDX1_LVT U2190 ( .A(n1609), .B(n1596), .CI(n2780), .S(O1[7]) );
  AO221X1_LVT U2191 ( .A1(n2781), .A2(n1621), .A3(n2781), .A4(n1610), .A5(
        n2777), .Y(n2780) );
  AND2X1_LVT U2192 ( .A1(n1621), .A2(n1610), .Y(n2777) );
  FADDX1_LVT U2193 ( .A(n1621), .B(n1610), .CI(n2781), .S(O1[6]) );
  AO21X1_LVT U2194 ( .A1(n2779), .A2(n2778), .A3(n2776), .Y(n2781) );
  OA22X1_LVT U2195 ( .A1(n1639), .A2(n1632), .A3(n1631), .A4(n1622), .Y(n2779)
         );
  FADDX1_LVT U2196 ( .A(n1631), .B(n1622), .CI(n2783), .S(O1[5]) );
  OA22X1_LVT U2197 ( .A1(n2778), .A2(n2782), .A3(n1639), .A4(n1632), .Y(n2783)
         );
  AND2X1_LVT U2198 ( .A1(n1639), .A2(n1632), .Y(n2782) );
  FADDX1_LVT U2199 ( .A(n2778), .B(n1639), .CI(n1632), .S(O1[4]) );
  FADDX1_LVT U2200 ( .A(n1645), .B(n1640), .CI(n2786), .S(O1[3]) );
  AO21X1_LVT U2201 ( .A1(n551), .A2(n2784), .A3(n2785), .Y(n2786) );
  AND2X1_LVT U2202 ( .A1(n1646), .A2(n1648), .Y(n2785) );
  OR2X1_LVT U2203 ( .A1(n1646), .A2(n1648), .Y(n2784) );
  FADDX1_LVT U2204 ( .A(n551), .B(n1646), .CI(n1648), .S(O1[2]) );
  NAND3X0_LVT U2205 ( .A1(I2[0]), .A2(I1[0]), .A3(I3[0]), .Y(n2589) );
  AND2X1_LVT U2206 ( .A1(I1[0]), .A2(I2[1]), .Y(n2235) );
  AND2X1_LVT U2207 ( .A1(I1[0]), .A2(I2[2]), .Y(n2234) );
  AND2X1_LVT U2208 ( .A1(I1[0]), .A2(I2[3]), .Y(n2233) );
  AND2X1_LVT U2209 ( .A1(I1[0]), .A2(n2557), .Y(n2232) );
  AND2X1_LVT U2210 ( .A1(I1[0]), .A2(I2[5]), .Y(n2231) );
  AND2X1_LVT U2211 ( .A1(I1[0]), .A2(n2558), .Y(n2230) );
  AND2X1_LVT U2212 ( .A1(I1[0]), .A2(n2559), .Y(n2229) );
  AND2X1_LVT U2213 ( .A1(I1[0]), .A2(I2[8]), .Y(n2228) );
  AND2X1_LVT U2214 ( .A1(I1[0]), .A2(n2560), .Y(n2227) );
  AND2X1_LVT U2215 ( .A1(I1[0]), .A2(I2[10]), .Y(n2226) );
  AND2X1_LVT U2216 ( .A1(I1[0]), .A2(I2[11]), .Y(n2225) );
  AND2X1_LVT U2217 ( .A1(I1[0]), .A2(n2561), .Y(n2224) );
  AND2X1_LVT U2218 ( .A1(I1[0]), .A2(n2562), .Y(n2223) );
  AND2X1_LVT U2219 ( .A1(I1[0]), .A2(n2563), .Y(n2222) );
  AND2X1_LVT U2220 ( .A1(I1[0]), .A2(I2[15]), .Y(n2221) );
  AND2X1_LVT U2221 ( .A1(I1[0]), .A2(I2[16]), .Y(n2220) );
  AND2X1_LVT U2222 ( .A1(I1[0]), .A2(I2[17]), .Y(n2219) );
  AND2X1_LVT U2223 ( .A1(I1[0]), .A2(I2[18]), .Y(n2218) );
  AND2X1_LVT U2224 ( .A1(I1[0]), .A2(I2[19]), .Y(n2217) );
  AND2X1_LVT U2225 ( .A1(I1[0]), .A2(n2564), .Y(n2216) );
  AND2X1_LVT U2226 ( .A1(I1[0]), .A2(I2[21]), .Y(n2215) );
  AND2X1_LVT U2227 ( .A1(I1[0]), .A2(n2565), .Y(n2214) );
  AND2X1_LVT U2228 ( .A1(I1[0]), .A2(I2[23]), .Y(n2213) );
  AND2X1_LVT U2229 ( .A1(I1[0]), .A2(I2[24]), .Y(n2212) );
  AND2X1_LVT U2230 ( .A1(I1[0]), .A2(I2[25]), .Y(n2211) );
  AND2X1_LVT U2231 ( .A1(I1[0]), .A2(I2[26]), .Y(n2210) );
  AND2X1_LVT U2232 ( .A1(I1[0]), .A2(I2[27]), .Y(n2209) );
  AND2X1_LVT U2233 ( .A1(I1[0]), .A2(n2566), .Y(n2208) );
  AND2X1_LVT U2234 ( .A1(I1[0]), .A2(I2[29]), .Y(n2207) );
  AND2X1_LVT U2235 ( .A1(I1[0]), .A2(n2567), .Y(n2206) );
  AND2X1_LVT U2236 ( .A1(I1[0]), .A2(n2568), .Y(n2205) );
  AND2X1_LVT U2237 ( .A1(I1[0]), .A2(I2[32]), .Y(n2204) );
  AND2X1_LVT U2238 ( .A1(I1[0]), .A2(I2[33]), .Y(n2203) );
  AND2X1_LVT U2239 ( .A1(I1[0]), .A2(I2[34]), .Y(n2202) );
  AND2X1_LVT U2240 ( .A1(I1[0]), .A2(I2[35]), .Y(n2201) );
  AND2X1_LVT U2241 ( .A1(I1[0]), .A2(n2569), .Y(n2200) );
  AND2X1_LVT U2242 ( .A1(I1[0]), .A2(n2570), .Y(n2199) );
  AND2X1_LVT U2243 ( .A1(I1[0]), .A2(n2571), .Y(n2198) );
  AND2X1_LVT U2244 ( .A1(I1[0]), .A2(I2[39]), .Y(n2197) );
  AND2X1_LVT U2245 ( .A1(I1[0]), .A2(I2[40]), .Y(n2196) );
  AND2X1_LVT U2246 ( .A1(I1[0]), .A2(I2[41]), .Y(n2195) );
  AND2X1_LVT U2247 ( .A1(I1[0]), .A2(I2[42]), .Y(n2194) );
  AND2X1_LVT U2248 ( .A1(I1[0]), .A2(I2[43]), .Y(n2193) );
  AND2X1_LVT U2249 ( .A1(I1[0]), .A2(n2572), .Y(n2192) );
  AND2X1_LVT U2250 ( .A1(I1[0]), .A2(n2573), .Y(n2191) );
  AND2X1_LVT U2251 ( .A1(I1[0]), .A2(n2574), .Y(n2190) );
  AND2X1_LVT U2252 ( .A1(I1[0]), .A2(I2[47]), .Y(n2189) );
  AND2X1_LVT U2253 ( .A1(I1[0]), .A2(I2[48]), .Y(n2188) );
  AND2X1_LVT U2254 ( .A1(I1[0]), .A2(I2[49]), .Y(n2187) );
  AND2X1_LVT U2255 ( .A1(I1[0]), .A2(I2[50]), .Y(n2186) );
  AND2X1_LVT U2256 ( .A1(I1[0]), .A2(I2[51]), .Y(n2185) );
  AND2X1_LVT U2257 ( .A1(I1[0]), .A2(n2575), .Y(n2184) );
  AND2X1_LVT U2258 ( .A1(I1[0]), .A2(n2576), .Y(n2183) );
  AND2X1_LVT U2259 ( .A1(I1[0]), .A2(n2577), .Y(n2182) );
  AND2X1_LVT U2260 ( .A1(I1[0]), .A2(n2578), .Y(n2181) );
  AND2X1_LVT U2261 ( .A1(I1[0]), .A2(n2579), .Y(n2180) );
  AND2X1_LVT U2262 ( .A1(I1[0]), .A2(n2580), .Y(n2179) );
  AND2X1_LVT U2263 ( .A1(I1[0]), .A2(I2[58]), .Y(n2178) );
  AND2X1_LVT U2264 ( .A1(I1[0]), .A2(I2[59]), .Y(n2177) );
  AND2X1_LVT U2265 ( .A1(I1[0]), .A2(n2581), .Y(n2176) );
  AND2X1_LVT U2266 ( .A1(I1[0]), .A2(n2582), .Y(n2175) );
  AND2X1_LVT U2267 ( .A1(I1[0]), .A2(I2[62]), .Y(n2174) );
  AND2X1_LVT U2268 ( .A1(I1[0]), .A2(n2583), .Y(n2173) );
  NAND2X0_LVT U2269 ( .A1(I2[64]), .A2(I1[0]), .Y(n2172) );
  AND2X1_LVT U2270 ( .A1(I2[0]), .A2(I1[1]), .Y(n2171) );
  AND2X1_LVT U2271 ( .A1(I2[1]), .A2(I1[1]), .Y(n2170) );
  AND2X1_LVT U2272 ( .A1(I2[2]), .A2(I1[1]), .Y(n2169) );
  AND2X1_LVT U2273 ( .A1(I2[3]), .A2(I1[1]), .Y(n2168) );
  AND2X1_LVT U2274 ( .A1(n2557), .A2(I1[1]), .Y(n2167) );
  AND2X1_LVT U2275 ( .A1(I2[5]), .A2(I1[1]), .Y(n2166) );
  AND2X1_LVT U2276 ( .A1(n2558), .A2(I1[1]), .Y(n2165) );
  AND2X1_LVT U2277 ( .A1(n2559), .A2(I1[1]), .Y(n2164) );
  AND2X1_LVT U2278 ( .A1(I2[8]), .A2(I1[1]), .Y(n2163) );
  AND2X1_LVT U2279 ( .A1(n2560), .A2(I1[1]), .Y(n2162) );
  AND2X1_LVT U2280 ( .A1(I2[10]), .A2(I1[1]), .Y(n2161) );
  AND2X1_LVT U2281 ( .A1(I2[11]), .A2(I1[1]), .Y(n2160) );
  AND2X1_LVT U2282 ( .A1(n2561), .A2(I1[1]), .Y(n2159) );
  AND2X1_LVT U2283 ( .A1(n2562), .A2(I1[1]), .Y(n2158) );
  AND2X1_LVT U2284 ( .A1(n2563), .A2(I1[1]), .Y(n2157) );
  AND2X1_LVT U2285 ( .A1(I2[15]), .A2(I1[1]), .Y(n2156) );
  AND2X1_LVT U2286 ( .A1(I2[16]), .A2(I1[1]), .Y(n2155) );
  AND2X1_LVT U2287 ( .A1(I2[17]), .A2(I1[1]), .Y(n2154) );
  AND2X1_LVT U2288 ( .A1(I2[18]), .A2(I1[1]), .Y(n2153) );
  AND2X1_LVT U2289 ( .A1(I2[19]), .A2(I1[1]), .Y(n2152) );
  AND2X1_LVT U2290 ( .A1(n2564), .A2(I1[1]), .Y(n2151) );
  AND2X1_LVT U2291 ( .A1(I2[21]), .A2(I1[1]), .Y(n2150) );
  AND2X1_LVT U2292 ( .A1(n2565), .A2(I1[1]), .Y(n2149) );
  AND2X1_LVT U2293 ( .A1(I2[23]), .A2(I1[1]), .Y(n2148) );
  AND2X1_LVT U2294 ( .A1(I2[24]), .A2(I1[1]), .Y(n2147) );
  AND2X1_LVT U2295 ( .A1(I2[25]), .A2(I1[1]), .Y(n2146) );
  AND2X1_LVT U2296 ( .A1(I2[26]), .A2(I1[1]), .Y(n2145) );
  AND2X1_LVT U2297 ( .A1(I2[27]), .A2(I1[1]), .Y(n2144) );
  AND2X1_LVT U2298 ( .A1(n2566), .A2(I1[1]), .Y(n2143) );
  AND2X1_LVT U2299 ( .A1(I2[29]), .A2(I1[1]), .Y(n2142) );
  AND2X1_LVT U2300 ( .A1(n2567), .A2(I1[1]), .Y(n2141) );
  AND2X1_LVT U2301 ( .A1(n2568), .A2(I1[1]), .Y(n2140) );
  AND2X1_LVT U2302 ( .A1(I2[32]), .A2(I1[1]), .Y(n2139) );
  AND2X1_LVT U2303 ( .A1(I2[33]), .A2(I1[1]), .Y(n2138) );
  AND2X1_LVT U2304 ( .A1(I2[34]), .A2(I1[1]), .Y(n2137) );
  AND2X1_LVT U2305 ( .A1(I2[35]), .A2(I1[1]), .Y(n2136) );
  AND2X1_LVT U2306 ( .A1(n2569), .A2(I1[1]), .Y(n2135) );
  AND2X1_LVT U2307 ( .A1(n2570), .A2(I1[1]), .Y(n2134) );
  AND2X1_LVT U2308 ( .A1(n2571), .A2(I1[1]), .Y(n2133) );
  AND2X1_LVT U2309 ( .A1(I2[39]), .A2(I1[1]), .Y(n2132) );
  AND2X1_LVT U2310 ( .A1(I2[40]), .A2(I1[1]), .Y(n2131) );
  AND2X1_LVT U2311 ( .A1(I2[41]), .A2(I1[1]), .Y(n2130) );
  AND2X1_LVT U2312 ( .A1(I2[42]), .A2(I1[1]), .Y(n2129) );
  AND2X1_LVT U2313 ( .A1(I2[43]), .A2(I1[1]), .Y(n2128) );
  AND2X1_LVT U2314 ( .A1(n2572), .A2(I1[1]), .Y(n2127) );
  AND2X1_LVT U2315 ( .A1(n2573), .A2(I1[1]), .Y(n2126) );
  AND2X1_LVT U2316 ( .A1(n2574), .A2(I1[1]), .Y(n2125) );
  AND2X1_LVT U2317 ( .A1(I2[47]), .A2(I1[1]), .Y(n2124) );
  AND2X1_LVT U2318 ( .A1(I2[48]), .A2(I1[1]), .Y(n2123) );
  AND2X1_LVT U2319 ( .A1(I2[49]), .A2(I1[1]), .Y(n2122) );
  AND2X1_LVT U2320 ( .A1(I2[50]), .A2(I1[1]), .Y(n2121) );
  AND2X1_LVT U2321 ( .A1(I2[51]), .A2(I1[1]), .Y(n2120) );
  AND2X1_LVT U2322 ( .A1(n2575), .A2(I1[1]), .Y(n2119) );
  AND2X1_LVT U2323 ( .A1(n2576), .A2(I1[1]), .Y(n2118) );
  AND2X1_LVT U2324 ( .A1(n2577), .A2(I1[1]), .Y(n2117) );
  AND2X1_LVT U2325 ( .A1(n2578), .A2(I1[1]), .Y(n2116) );
  AND2X1_LVT U2326 ( .A1(n2579), .A2(I1[1]), .Y(n2115) );
  AND2X1_LVT U2327 ( .A1(n2580), .A2(I1[1]), .Y(n2114) );
  AND2X1_LVT U2328 ( .A1(I2[58]), .A2(I1[1]), .Y(n2113) );
  AND2X1_LVT U2329 ( .A1(I2[59]), .A2(I1[1]), .Y(n2112) );
  AND2X1_LVT U2330 ( .A1(n2581), .A2(I1[1]), .Y(n2111) );
  AND2X1_LVT U2331 ( .A1(n2582), .A2(I1[1]), .Y(n2110) );
  AND2X1_LVT U2332 ( .A1(I2[62]), .A2(I1[1]), .Y(n2109) );
  AND2X1_LVT U2333 ( .A1(n2583), .A2(I1[1]), .Y(n2108) );
  NAND2X0_LVT U2334 ( .A1(I2[64]), .A2(I1[1]), .Y(n2107) );
  AND2X1_LVT U2335 ( .A1(I2[0]), .A2(I1[2]), .Y(n2106) );
  AND2X1_LVT U2336 ( .A1(I2[1]), .A2(I1[2]), .Y(n2105) );
  AND2X1_LVT U2337 ( .A1(I2[2]), .A2(I1[2]), .Y(n2104) );
  AND2X1_LVT U2338 ( .A1(I2[3]), .A2(I1[2]), .Y(n2103) );
  AND2X1_LVT U2339 ( .A1(n2557), .A2(I1[2]), .Y(n2102) );
  AND2X1_LVT U2340 ( .A1(I2[5]), .A2(I1[2]), .Y(n2101) );
  AND2X1_LVT U2341 ( .A1(n2558), .A2(I1[2]), .Y(n2100) );
  AND2X1_LVT U2342 ( .A1(n2559), .A2(I1[2]), .Y(n2099) );
  AND2X1_LVT U2343 ( .A1(I2[8]), .A2(I1[2]), .Y(n2098) );
  AND2X1_LVT U2344 ( .A1(n2560), .A2(I1[2]), .Y(n2097) );
  AND2X1_LVT U2345 ( .A1(I2[10]), .A2(I1[2]), .Y(n2096) );
  AND2X1_LVT U2346 ( .A1(I2[11]), .A2(I1[2]), .Y(n2095) );
  AND2X1_LVT U2347 ( .A1(n2561), .A2(I1[2]), .Y(n2094) );
  AND2X1_LVT U2348 ( .A1(n2562), .A2(I1[2]), .Y(n2093) );
  AND2X1_LVT U2349 ( .A1(n2563), .A2(I1[2]), .Y(n2092) );
  AND2X1_LVT U2350 ( .A1(I2[15]), .A2(I1[2]), .Y(n2091) );
  AND2X1_LVT U2351 ( .A1(I2[16]), .A2(I1[2]), .Y(n2090) );
  AND2X1_LVT U2352 ( .A1(I2[17]), .A2(I1[2]), .Y(n2089) );
  AND2X1_LVT U2353 ( .A1(I2[18]), .A2(I1[2]), .Y(n2088) );
  AND2X1_LVT U2354 ( .A1(I2[19]), .A2(I1[2]), .Y(n2087) );
  AND2X1_LVT U2355 ( .A1(n2564), .A2(I1[2]), .Y(n2086) );
  AND2X1_LVT U2356 ( .A1(I2[21]), .A2(I1[2]), .Y(n2085) );
  AND2X1_LVT U2357 ( .A1(n2565), .A2(I1[2]), .Y(n2084) );
  AND2X1_LVT U2358 ( .A1(I2[23]), .A2(I1[2]), .Y(n2083) );
  AND2X1_LVT U2359 ( .A1(I2[24]), .A2(I1[2]), .Y(n2082) );
  AND2X1_LVT U2360 ( .A1(I2[25]), .A2(I1[2]), .Y(n2081) );
  AND2X1_LVT U2361 ( .A1(I2[26]), .A2(I1[2]), .Y(n2080) );
  AND2X1_LVT U2362 ( .A1(I2[27]), .A2(I1[2]), .Y(n2079) );
  AND2X1_LVT U2363 ( .A1(n2566), .A2(I1[2]), .Y(n2078) );
  AND2X1_LVT U2364 ( .A1(I2[29]), .A2(I1[2]), .Y(n2077) );
  AND2X1_LVT U2365 ( .A1(n2567), .A2(I1[2]), .Y(n2076) );
  AND2X1_LVT U2366 ( .A1(n2568), .A2(I1[2]), .Y(n2075) );
  AND2X1_LVT U2367 ( .A1(I2[32]), .A2(I1[2]), .Y(n2074) );
  AND2X1_LVT U2368 ( .A1(I2[33]), .A2(I1[2]), .Y(n2073) );
  AND2X1_LVT U2369 ( .A1(I2[34]), .A2(I1[2]), .Y(n2072) );
  AND2X1_LVT U2370 ( .A1(I2[35]), .A2(I1[2]), .Y(n2071) );
  AND2X1_LVT U2371 ( .A1(n2569), .A2(I1[2]), .Y(n2070) );
  AND2X1_LVT U2372 ( .A1(n2570), .A2(I1[2]), .Y(n2069) );
  AND2X1_LVT U2373 ( .A1(n2571), .A2(I1[2]), .Y(n2068) );
  AND2X1_LVT U2374 ( .A1(I2[39]), .A2(I1[2]), .Y(n2067) );
  AND2X1_LVT U2375 ( .A1(I2[40]), .A2(I1[2]), .Y(n2066) );
  AND2X1_LVT U2376 ( .A1(I2[41]), .A2(I1[2]), .Y(n2065) );
  AND2X1_LVT U2377 ( .A1(I2[42]), .A2(I1[2]), .Y(n2064) );
  AND2X1_LVT U2378 ( .A1(I2[43]), .A2(I1[2]), .Y(n2063) );
  AND2X1_LVT U2379 ( .A1(n2572), .A2(I1[2]), .Y(n2062) );
  AND2X1_LVT U2380 ( .A1(n2573), .A2(I1[2]), .Y(n2061) );
  AND2X1_LVT U2381 ( .A1(n2574), .A2(I1[2]), .Y(n2060) );
  AND2X1_LVT U2382 ( .A1(I2[47]), .A2(I1[2]), .Y(n2059) );
  AND2X1_LVT U2383 ( .A1(I2[48]), .A2(I1[2]), .Y(n2058) );
  AND2X1_LVT U2384 ( .A1(I2[49]), .A2(I1[2]), .Y(n2057) );
  AND2X1_LVT U2385 ( .A1(I2[50]), .A2(I1[2]), .Y(n2056) );
  AND2X1_LVT U2386 ( .A1(I2[51]), .A2(I1[2]), .Y(n2055) );
  AND2X1_LVT U2387 ( .A1(n2575), .A2(I1[2]), .Y(n2054) );
  AND2X1_LVT U2388 ( .A1(n2576), .A2(I1[2]), .Y(n2053) );
  AND2X1_LVT U2389 ( .A1(n2577), .A2(I1[2]), .Y(n2052) );
  AND2X1_LVT U2390 ( .A1(n2578), .A2(I1[2]), .Y(n2051) );
  AND2X1_LVT U2391 ( .A1(n2579), .A2(I1[2]), .Y(n2050) );
  AND2X1_LVT U2392 ( .A1(n2580), .A2(I1[2]), .Y(n2049) );
  AND2X1_LVT U2393 ( .A1(I2[58]), .A2(I1[2]), .Y(n2048) );
  AND2X1_LVT U2394 ( .A1(I2[59]), .A2(I1[2]), .Y(n2047) );
  AND2X1_LVT U2395 ( .A1(n2581), .A2(I1[2]), .Y(n2046) );
  AND2X1_LVT U2396 ( .A1(n2582), .A2(I1[2]), .Y(n2045) );
  AND2X1_LVT U2397 ( .A1(I2[62]), .A2(I1[2]), .Y(n2044) );
  AND2X1_LVT U2398 ( .A1(n2583), .A2(I1[2]), .Y(n2043) );
  NAND2X0_LVT U2399 ( .A1(I2[64]), .A2(I1[2]), .Y(n2042) );
  AND2X1_LVT U2400 ( .A1(I2[0]), .A2(I1[3]), .Y(n2041) );
  AND2X1_LVT U2401 ( .A1(I2[1]), .A2(I1[3]), .Y(n2040) );
  AND2X1_LVT U2402 ( .A1(I2[2]), .A2(I1[3]), .Y(n2039) );
  AND2X1_LVT U2403 ( .A1(I2[3]), .A2(I1[3]), .Y(n2038) );
  AND2X1_LVT U2404 ( .A1(n2557), .A2(I1[3]), .Y(n2037) );
  AND2X1_LVT U2405 ( .A1(I2[5]), .A2(I1[3]), .Y(n2036) );
  AND2X1_LVT U2406 ( .A1(n2558), .A2(I1[3]), .Y(n2035) );
  AND2X1_LVT U2407 ( .A1(n2559), .A2(I1[3]), .Y(n2034) );
  AND2X1_LVT U2408 ( .A1(I2[8]), .A2(I1[3]), .Y(n2033) );
  AND2X1_LVT U2409 ( .A1(n2560), .A2(I1[3]), .Y(n2032) );
  AND2X1_LVT U2410 ( .A1(I2[10]), .A2(I1[3]), .Y(n2031) );
  AND2X1_LVT U2411 ( .A1(I2[11]), .A2(I1[3]), .Y(n2030) );
  AND2X1_LVT U2412 ( .A1(n2561), .A2(I1[3]), .Y(n2029) );
  AND2X1_LVT U2413 ( .A1(n2562), .A2(I1[3]), .Y(n2028) );
  AND2X1_LVT U2414 ( .A1(n2563), .A2(I1[3]), .Y(n2027) );
  AND2X1_LVT U2415 ( .A1(I2[15]), .A2(I1[3]), .Y(n2026) );
  AND2X1_LVT U2416 ( .A1(I2[16]), .A2(I1[3]), .Y(n2025) );
  AND2X1_LVT U2417 ( .A1(I2[17]), .A2(I1[3]), .Y(n2024) );
  AND2X1_LVT U2418 ( .A1(I2[18]), .A2(I1[3]), .Y(n2023) );
  AND2X1_LVT U2419 ( .A1(I2[19]), .A2(I1[3]), .Y(n2022) );
  AND2X1_LVT U2420 ( .A1(n2564), .A2(I1[3]), .Y(n2021) );
  AND2X1_LVT U2421 ( .A1(I2[21]), .A2(I1[3]), .Y(n2020) );
  AND2X1_LVT U2422 ( .A1(n2565), .A2(I1[3]), .Y(n2019) );
  AND2X1_LVT U2423 ( .A1(I2[23]), .A2(I1[3]), .Y(n2018) );
  AND2X1_LVT U2424 ( .A1(I2[24]), .A2(I1[3]), .Y(n2017) );
  AND2X1_LVT U2425 ( .A1(I2[25]), .A2(I1[3]), .Y(n2016) );
  AND2X1_LVT U2426 ( .A1(I2[26]), .A2(I1[3]), .Y(n2015) );
  AND2X1_LVT U2427 ( .A1(I2[27]), .A2(I1[3]), .Y(n2014) );
  AND2X1_LVT U2428 ( .A1(n2566), .A2(I1[3]), .Y(n2013) );
  AND2X1_LVT U2429 ( .A1(I2[29]), .A2(I1[3]), .Y(n2012) );
  AND2X1_LVT U2430 ( .A1(n2567), .A2(I1[3]), .Y(n2011) );
  AND2X1_LVT U2431 ( .A1(n2568), .A2(I1[3]), .Y(n2010) );
  AND2X1_LVT U2432 ( .A1(I2[32]), .A2(I1[3]), .Y(n2009) );
  AND2X1_LVT U2433 ( .A1(I2[33]), .A2(I1[3]), .Y(n2008) );
  AND2X1_LVT U2434 ( .A1(I2[34]), .A2(I1[3]), .Y(n2007) );
  AND2X1_LVT U2435 ( .A1(I2[35]), .A2(I1[3]), .Y(n2006) );
  AND2X1_LVT U2436 ( .A1(n2569), .A2(I1[3]), .Y(n2005) );
  AND2X1_LVT U2437 ( .A1(n2570), .A2(I1[3]), .Y(n2004) );
  AND2X1_LVT U2438 ( .A1(n2571), .A2(I1[3]), .Y(n2003) );
  AND2X1_LVT U2439 ( .A1(I2[39]), .A2(I1[3]), .Y(n2002) );
  AND2X1_LVT U2440 ( .A1(I2[40]), .A2(I1[3]), .Y(n2001) );
  AND2X1_LVT U2441 ( .A1(I2[41]), .A2(I1[3]), .Y(n2000) );
  AND2X1_LVT U2442 ( .A1(I2[42]), .A2(I1[3]), .Y(n1999) );
  AND2X1_LVT U2443 ( .A1(I2[43]), .A2(I1[3]), .Y(n1998) );
  AND2X1_LVT U2444 ( .A1(n2572), .A2(I1[3]), .Y(n1997) );
  AND2X1_LVT U2445 ( .A1(n2573), .A2(I1[3]), .Y(n1996) );
  AND2X1_LVT U2446 ( .A1(n2574), .A2(I1[3]), .Y(n1995) );
  AND2X1_LVT U2447 ( .A1(I2[47]), .A2(I1[3]), .Y(n1994) );
  AND2X1_LVT U2448 ( .A1(I2[48]), .A2(I1[3]), .Y(n1993) );
  AND2X1_LVT U2449 ( .A1(I2[49]), .A2(I1[3]), .Y(n1992) );
  AND2X1_LVT U2450 ( .A1(I2[50]), .A2(I1[3]), .Y(n1991) );
  AND2X1_LVT U2451 ( .A1(I2[51]), .A2(I1[3]), .Y(n1990) );
  AND2X1_LVT U2452 ( .A1(n2575), .A2(I1[3]), .Y(n1989) );
  AND2X1_LVT U2453 ( .A1(n2576), .A2(I1[3]), .Y(n1988) );
  AND2X1_LVT U2454 ( .A1(n2577), .A2(I1[3]), .Y(n1987) );
  AND2X1_LVT U2455 ( .A1(n2578), .A2(I1[3]), .Y(n1986) );
  AND2X1_LVT U2456 ( .A1(n2579), .A2(I1[3]), .Y(n1985) );
  AND2X1_LVT U2457 ( .A1(n2580), .A2(I1[3]), .Y(n1984) );
  AND2X1_LVT U2458 ( .A1(I2[58]), .A2(I1[3]), .Y(n1983) );
  AND2X1_LVT U2459 ( .A1(I2[59]), .A2(I1[3]), .Y(n1982) );
  AND2X1_LVT U2460 ( .A1(n2581), .A2(I1[3]), .Y(n1981) );
  AND2X1_LVT U2461 ( .A1(n2582), .A2(I1[3]), .Y(n1980) );
  AND2X1_LVT U2462 ( .A1(I2[62]), .A2(I1[3]), .Y(n1979) );
  AND2X1_LVT U2463 ( .A1(n2583), .A2(I1[3]), .Y(n1978) );
  NAND2X0_LVT U2464 ( .A1(I2[64]), .A2(I1[3]), .Y(n1977) );
  AND2X1_LVT U2465 ( .A1(I2[0]), .A2(I1[4]), .Y(n1976) );
  AND2X1_LVT U2466 ( .A1(I2[1]), .A2(I1[4]), .Y(n1975) );
  AND2X1_LVT U2467 ( .A1(I2[2]), .A2(I1[4]), .Y(n1974) );
  AND2X1_LVT U2468 ( .A1(I2[3]), .A2(I1[4]), .Y(n1973) );
  AND2X1_LVT U2469 ( .A1(n2557), .A2(I1[4]), .Y(n1972) );
  AND2X1_LVT U2470 ( .A1(I2[5]), .A2(I1[4]), .Y(n1971) );
  AND2X1_LVT U2471 ( .A1(n2558), .A2(I1[4]), .Y(n1970) );
  AND2X1_LVT U2472 ( .A1(n2559), .A2(I1[4]), .Y(n1969) );
  AND2X1_LVT U2473 ( .A1(I2[8]), .A2(I1[4]), .Y(n1968) );
  AND2X1_LVT U2474 ( .A1(n2560), .A2(I1[4]), .Y(n1967) );
  AND2X1_LVT U2475 ( .A1(I2[10]), .A2(I1[4]), .Y(n1966) );
  AND2X1_LVT U2476 ( .A1(I2[11]), .A2(I1[4]), .Y(n1965) );
  AND2X1_LVT U2477 ( .A1(n2561), .A2(I1[4]), .Y(n1964) );
  AND2X1_LVT U2478 ( .A1(n2562), .A2(I1[4]), .Y(n1963) );
  AND2X1_LVT U2479 ( .A1(n2563), .A2(I1[4]), .Y(n1962) );
  AND2X1_LVT U2480 ( .A1(I2[15]), .A2(I1[4]), .Y(n1961) );
  AND2X1_LVT U2481 ( .A1(I2[16]), .A2(I1[4]), .Y(n1960) );
  AND2X1_LVT U2482 ( .A1(I2[17]), .A2(I1[4]), .Y(n1959) );
  AND2X1_LVT U2483 ( .A1(I2[18]), .A2(I1[4]), .Y(n1958) );
  AND2X1_LVT U2484 ( .A1(I2[19]), .A2(I1[4]), .Y(n1957) );
  AND2X1_LVT U2485 ( .A1(n2564), .A2(I1[4]), .Y(n1956) );
  AND2X1_LVT U2486 ( .A1(I2[21]), .A2(I1[4]), .Y(n1955) );
  AND2X1_LVT U2487 ( .A1(n2565), .A2(I1[4]), .Y(n1954) );
  AND2X1_LVT U2488 ( .A1(I2[23]), .A2(I1[4]), .Y(n1953) );
  AND2X1_LVT U2489 ( .A1(I2[24]), .A2(I1[4]), .Y(n1952) );
  AND2X1_LVT U2490 ( .A1(I2[25]), .A2(I1[4]), .Y(n1951) );
  AND2X1_LVT U2491 ( .A1(I2[26]), .A2(I1[4]), .Y(n1950) );
  AND2X1_LVT U2492 ( .A1(I2[27]), .A2(I1[4]), .Y(n1949) );
  AND2X1_LVT U2493 ( .A1(n2566), .A2(I1[4]), .Y(n1948) );
  AND2X1_LVT U2494 ( .A1(I2[29]), .A2(I1[4]), .Y(n1947) );
  AND2X1_LVT U2495 ( .A1(n2567), .A2(I1[4]), .Y(n1946) );
  AND2X1_LVT U2496 ( .A1(n2568), .A2(I1[4]), .Y(n1945) );
  AND2X1_LVT U2497 ( .A1(I2[32]), .A2(I1[4]), .Y(n1944) );
  AND2X1_LVT U2498 ( .A1(I2[33]), .A2(I1[4]), .Y(n1943) );
  AND2X1_LVT U2499 ( .A1(I2[34]), .A2(I1[4]), .Y(n1942) );
  AND2X1_LVT U2500 ( .A1(I2[35]), .A2(I1[4]), .Y(n1941) );
  AND2X1_LVT U2501 ( .A1(n2569), .A2(I1[4]), .Y(n1940) );
  AND2X1_LVT U2502 ( .A1(n2570), .A2(I1[4]), .Y(n1939) );
  AND2X1_LVT U2503 ( .A1(n2571), .A2(I1[4]), .Y(n1938) );
  AND2X1_LVT U2504 ( .A1(I2[39]), .A2(I1[4]), .Y(n1937) );
  AND2X1_LVT U2505 ( .A1(I2[40]), .A2(I1[4]), .Y(n1936) );
  AND2X1_LVT U2506 ( .A1(I2[41]), .A2(I1[4]), .Y(n1935) );
  AND2X1_LVT U2507 ( .A1(I2[42]), .A2(I1[4]), .Y(n1934) );
  AND2X1_LVT U2508 ( .A1(I2[43]), .A2(I1[4]), .Y(n1933) );
  AND2X1_LVT U2509 ( .A1(n2572), .A2(I1[4]), .Y(n1932) );
  AND2X1_LVT U2510 ( .A1(n2573), .A2(I1[4]), .Y(n1931) );
  AND2X1_LVT U2511 ( .A1(n2574), .A2(I1[4]), .Y(n1930) );
  AND2X1_LVT U2512 ( .A1(I2[47]), .A2(I1[4]), .Y(n1929) );
  AND2X1_LVT U2513 ( .A1(I2[48]), .A2(I1[4]), .Y(n1928) );
  AND2X1_LVT U2514 ( .A1(I2[49]), .A2(I1[4]), .Y(n1927) );
  AND2X1_LVT U2515 ( .A1(I2[50]), .A2(I1[4]), .Y(n1926) );
  AND2X1_LVT U2516 ( .A1(I2[51]), .A2(I1[4]), .Y(n1925) );
  AND2X1_LVT U2517 ( .A1(n2575), .A2(I1[4]), .Y(n1924) );
  AND2X1_LVT U2518 ( .A1(n2576), .A2(I1[4]), .Y(n1923) );
  AND2X1_LVT U2519 ( .A1(n2577), .A2(I1[4]), .Y(n1922) );
  AND2X1_LVT U2520 ( .A1(n2578), .A2(I1[4]), .Y(n1921) );
  AND2X1_LVT U2521 ( .A1(n2579), .A2(I1[4]), .Y(n1920) );
  AND2X1_LVT U2522 ( .A1(n2580), .A2(I1[4]), .Y(n1919) );
  AND2X1_LVT U2523 ( .A1(I2[58]), .A2(I1[4]), .Y(n1918) );
  AND2X1_LVT U2524 ( .A1(I2[59]), .A2(I1[4]), .Y(n1917) );
  AND2X1_LVT U2525 ( .A1(n2581), .A2(I1[4]), .Y(n1916) );
  AND2X1_LVT U2526 ( .A1(n2582), .A2(I1[4]), .Y(n1915) );
  AND2X1_LVT U2527 ( .A1(I2[62]), .A2(I1[4]), .Y(n1914) );
  AND2X1_LVT U2528 ( .A1(n2583), .A2(I1[4]), .Y(n1913) );
  NAND2X0_LVT U2529 ( .A1(I2[64]), .A2(I1[4]), .Y(n1912) );
  AND2X1_LVT U2530 ( .A1(I2[0]), .A2(I1[5]), .Y(n1911) );
  AND2X1_LVT U2531 ( .A1(I2[1]), .A2(I1[5]), .Y(n1910) );
  AND2X1_LVT U2532 ( .A1(I2[2]), .A2(I1[5]), .Y(n1909) );
  AND2X1_LVT U2533 ( .A1(I2[3]), .A2(I1[5]), .Y(n1908) );
  AND2X1_LVT U2534 ( .A1(n2557), .A2(n2584), .Y(n1907) );
  AND2X1_LVT U2535 ( .A1(I2[5]), .A2(n2584), .Y(n1906) );
  AND2X1_LVT U2536 ( .A1(n2558), .A2(n2584), .Y(n1905) );
  AND2X1_LVT U2537 ( .A1(n2559), .A2(n2584), .Y(n1904) );
  AND2X1_LVT U2538 ( .A1(I2[8]), .A2(n2584), .Y(n1903) );
  AND2X1_LVT U2539 ( .A1(n2560), .A2(n2584), .Y(n1902) );
  AND2X1_LVT U2540 ( .A1(I2[10]), .A2(n2584), .Y(n1901) );
  AND2X1_LVT U2541 ( .A1(I2[11]), .A2(n2584), .Y(n1900) );
  AND2X1_LVT U2542 ( .A1(n2561), .A2(I1[5]), .Y(n1899) );
  AND2X1_LVT U2543 ( .A1(n2562), .A2(n2584), .Y(n1898) );
  AND2X1_LVT U2544 ( .A1(n2563), .A2(n2584), .Y(n1897) );
  AND2X1_LVT U2545 ( .A1(I2[15]), .A2(n2584), .Y(n1896) );
  AND2X1_LVT U2546 ( .A1(I2[16]), .A2(n2584), .Y(n1895) );
  AND2X1_LVT U2547 ( .A1(I2[17]), .A2(I1[5]), .Y(n1894) );
  AND2X1_LVT U2548 ( .A1(I2[18]), .A2(n2584), .Y(n1893) );
  AND2X1_LVT U2549 ( .A1(I2[19]), .A2(n2584), .Y(n1892) );
  AND2X1_LVT U2550 ( .A1(n2564), .A2(n2584), .Y(n1891) );
  AND2X1_LVT U2551 ( .A1(I2[21]), .A2(n2584), .Y(n1890) );
  AND2X1_LVT U2552 ( .A1(n2565), .A2(I1[5]), .Y(n1889) );
  AND2X1_LVT U2553 ( .A1(I2[23]), .A2(I1[5]), .Y(n1888) );
  AND2X1_LVT U2554 ( .A1(I2[24]), .A2(n2584), .Y(n1887) );
  AND2X1_LVT U2555 ( .A1(I2[25]), .A2(n2584), .Y(n1886) );
  AND2X1_LVT U2556 ( .A1(I2[26]), .A2(n2584), .Y(n1885) );
  AND2X1_LVT U2557 ( .A1(I2[27]), .A2(n2584), .Y(n1884) );
  AND2X1_LVT U2558 ( .A1(n2566), .A2(n2584), .Y(n1883) );
  AND2X1_LVT U2559 ( .A1(I2[29]), .A2(n2584), .Y(n1882) );
  AND2X1_LVT U2560 ( .A1(n2567), .A2(n2584), .Y(n1881) );
  AND2X1_LVT U2561 ( .A1(n2568), .A2(n2584), .Y(n1880) );
  AND2X1_LVT U2562 ( .A1(I2[32]), .A2(n2584), .Y(n1879) );
  AND2X1_LVT U2563 ( .A1(I2[33]), .A2(n2584), .Y(n1878) );
  AND2X1_LVT U2564 ( .A1(I2[34]), .A2(n2584), .Y(n1877) );
  AND2X1_LVT U2565 ( .A1(I2[35]), .A2(n2584), .Y(n1876) );
  AND2X1_LVT U2566 ( .A1(n2569), .A2(n2584), .Y(n1875) );
  AND2X1_LVT U2567 ( .A1(n2570), .A2(n2584), .Y(n1874) );
  AND2X1_LVT U2568 ( .A1(n2571), .A2(n2584), .Y(n1873) );
  AND2X1_LVT U2569 ( .A1(I2[39]), .A2(n2584), .Y(n1872) );
  AND2X1_LVT U2570 ( .A1(I2[40]), .A2(n2584), .Y(n1871) );
  AND2X1_LVT U2571 ( .A1(I2[41]), .A2(n2584), .Y(n1870) );
  AND2X1_LVT U2572 ( .A1(I2[42]), .A2(n2584), .Y(n1869) );
  AND2X1_LVT U2573 ( .A1(I2[43]), .A2(n2584), .Y(n1868) );
  AND2X1_LVT U2574 ( .A1(n2572), .A2(n2584), .Y(n1867) );
  AND2X1_LVT U2575 ( .A1(n2573), .A2(n2584), .Y(n1866) );
  AND2X1_LVT U2576 ( .A1(n2574), .A2(n2584), .Y(n1865) );
  AND2X1_LVT U2577 ( .A1(I2[47]), .A2(n2584), .Y(n1864) );
  AND2X1_LVT U2578 ( .A1(I2[48]), .A2(n2584), .Y(n1863) );
  AND2X1_LVT U2579 ( .A1(I2[49]), .A2(n2584), .Y(n1862) );
  AND2X1_LVT U2580 ( .A1(I2[50]), .A2(n2584), .Y(n1861) );
  AND2X1_LVT U2581 ( .A1(I2[51]), .A2(n2584), .Y(n1860) );
  AND2X1_LVT U2582 ( .A1(n2575), .A2(n2584), .Y(n1859) );
  AND2X1_LVT U2583 ( .A1(n2576), .A2(n2584), .Y(n1858) );
  AND2X1_LVT U2584 ( .A1(n2577), .A2(n2584), .Y(n1857) );
  AND2X1_LVT U2585 ( .A1(n2578), .A2(n2584), .Y(n1856) );
  AND2X1_LVT U2586 ( .A1(n2579), .A2(n2584), .Y(n1855) );
  AND2X1_LVT U2587 ( .A1(n2580), .A2(n2584), .Y(n1854) );
  AND2X1_LVT U2588 ( .A1(I2[58]), .A2(n2584), .Y(n1853) );
  AND2X1_LVT U2589 ( .A1(I2[59]), .A2(n2584), .Y(n1852) );
  AND2X1_LVT U2590 ( .A1(n2581), .A2(n2584), .Y(n1851) );
  AND2X1_LVT U2591 ( .A1(n2582), .A2(n2584), .Y(n1850) );
  AND2X1_LVT U2592 ( .A1(I2[62]), .A2(n2584), .Y(n1849) );
  AND2X1_LVT U2593 ( .A1(n2583), .A2(n2584), .Y(n1848) );
  NAND2X0_LVT U2594 ( .A1(I2[64]), .A2(n2584), .Y(n1847) );
  AND2X1_LVT U2595 ( .A1(I2[0]), .A2(I1[6]), .Y(n1846) );
  AND2X1_LVT U2596 ( .A1(I2[1]), .A2(I1[6]), .Y(n1845) );
  AND2X1_LVT U2597 ( .A1(I2[2]), .A2(I1[6]), .Y(n1844) );
  AND2X1_LVT U2598 ( .A1(I2[3]), .A2(I1[6]), .Y(n1843) );
  AND2X1_LVT U2599 ( .A1(n2557), .A2(I1[6]), .Y(n1842) );
  AND2X1_LVT U2600 ( .A1(I2[5]), .A2(I1[6]), .Y(n1841) );
  AND2X1_LVT U2601 ( .A1(n2558), .A2(I1[6]), .Y(n1840) );
  AND2X1_LVT U2602 ( .A1(n2559), .A2(I1[6]), .Y(n1839) );
  AND2X1_LVT U2603 ( .A1(I2[8]), .A2(I1[6]), .Y(n1838) );
  AND2X1_LVT U2604 ( .A1(n2560), .A2(I1[6]), .Y(n1837) );
  AND2X1_LVT U2605 ( .A1(I2[10]), .A2(I1[6]), .Y(n1836) );
  AND2X1_LVT U2606 ( .A1(I2[11]), .A2(I1[6]), .Y(n1835) );
  AND2X1_LVT U2607 ( .A1(n2561), .A2(I1[6]), .Y(n1834) );
  AND2X1_LVT U2608 ( .A1(n2562), .A2(I1[6]), .Y(n1833) );
  AND2X1_LVT U2609 ( .A1(n2563), .A2(I1[6]), .Y(n1832) );
  AND2X1_LVT U2610 ( .A1(I2[15]), .A2(I1[6]), .Y(n1831) );
  AND2X1_LVT U2611 ( .A1(I2[16]), .A2(I1[6]), .Y(n1830) );
  AND2X1_LVT U2612 ( .A1(I2[17]), .A2(I1[6]), .Y(n1829) );
  AND2X1_LVT U2613 ( .A1(I2[18]), .A2(I1[6]), .Y(n1828) );
  AND2X1_LVT U2614 ( .A1(I2[19]), .A2(I1[6]), .Y(n1827) );
  AND2X1_LVT U2615 ( .A1(n2564), .A2(I1[6]), .Y(n1826) );
  AND2X1_LVT U2616 ( .A1(I2[21]), .A2(I1[6]), .Y(n1825) );
  AND2X1_LVT U2617 ( .A1(n2565), .A2(I1[6]), .Y(n1824) );
  AND2X1_LVT U2618 ( .A1(I2[23]), .A2(I1[6]), .Y(n1823) );
  AND2X1_LVT U2619 ( .A1(I2[24]), .A2(I1[6]), .Y(n1822) );
  AND2X1_LVT U2620 ( .A1(I2[25]), .A2(I1[6]), .Y(n1821) );
  AND2X1_LVT U2621 ( .A1(I2[26]), .A2(I1[6]), .Y(n1820) );
  AND2X1_LVT U2622 ( .A1(I2[27]), .A2(I1[6]), .Y(n1819) );
  AND2X1_LVT U2623 ( .A1(n2566), .A2(I1[6]), .Y(n1818) );
  AND2X1_LVT U2624 ( .A1(I2[29]), .A2(I1[6]), .Y(n1817) );
  AND2X1_LVT U2625 ( .A1(n2567), .A2(I1[6]), .Y(n1816) );
  AND2X1_LVT U2626 ( .A1(n2568), .A2(I1[6]), .Y(n1815) );
  AND2X1_LVT U2627 ( .A1(I2[32]), .A2(I1[6]), .Y(n1814) );
  AND2X1_LVT U2628 ( .A1(I2[33]), .A2(I1[6]), .Y(n1813) );
  AND2X1_LVT U2629 ( .A1(I2[34]), .A2(I1[6]), .Y(n1812) );
  AND2X1_LVT U2630 ( .A1(I2[35]), .A2(I1[6]), .Y(n1811) );
  AND2X1_LVT U2631 ( .A1(n2569), .A2(I1[6]), .Y(n1810) );
  AND2X1_LVT U2632 ( .A1(n2570), .A2(I1[6]), .Y(n1809) );
  AND2X1_LVT U2633 ( .A1(n2571), .A2(I1[6]), .Y(n1808) );
  AND2X1_LVT U2634 ( .A1(I2[39]), .A2(I1[6]), .Y(n1807) );
  AND2X1_LVT U2635 ( .A1(I2[40]), .A2(I1[6]), .Y(n1806) );
  AND2X1_LVT U2636 ( .A1(I2[41]), .A2(I1[6]), .Y(n1805) );
  AND2X1_LVT U2637 ( .A1(I2[42]), .A2(I1[6]), .Y(n1804) );
  AND2X1_LVT U2638 ( .A1(I2[43]), .A2(I1[6]), .Y(n1803) );
  AND2X1_LVT U2639 ( .A1(n2572), .A2(I1[6]), .Y(n1802) );
  AND2X1_LVT U2640 ( .A1(n2573), .A2(I1[6]), .Y(n1801) );
  AND2X1_LVT U2641 ( .A1(n2574), .A2(I1[6]), .Y(n1800) );
  AND2X1_LVT U2642 ( .A1(I2[47]), .A2(I1[6]), .Y(n1799) );
  AND2X1_LVT U2643 ( .A1(I2[48]), .A2(I1[6]), .Y(n1798) );
  AND2X1_LVT U2644 ( .A1(I2[49]), .A2(I1[6]), .Y(n1797) );
  AND2X1_LVT U2645 ( .A1(I2[50]), .A2(I1[6]), .Y(n1796) );
  AND2X1_LVT U2646 ( .A1(I2[51]), .A2(I1[6]), .Y(n1795) );
  AND2X1_LVT U2647 ( .A1(n2575), .A2(I1[6]), .Y(n1794) );
  AND2X1_LVT U2648 ( .A1(n2576), .A2(I1[6]), .Y(n1793) );
  AND2X1_LVT U2649 ( .A1(n2577), .A2(I1[6]), .Y(n1792) );
  AND2X1_LVT U2650 ( .A1(n2578), .A2(I1[6]), .Y(n1791) );
  AND2X1_LVT U2651 ( .A1(n2579), .A2(I1[6]), .Y(n1790) );
  AND2X1_LVT U2652 ( .A1(n2580), .A2(I1[6]), .Y(n1789) );
  AND2X1_LVT U2653 ( .A1(I2[58]), .A2(I1[6]), .Y(n1788) );
  AND2X1_LVT U2654 ( .A1(I2[59]), .A2(I1[6]), .Y(n1787) );
  AND2X1_LVT U2655 ( .A1(n2581), .A2(I1[6]), .Y(n1786) );
  AND2X1_LVT U2656 ( .A1(n2582), .A2(I1[6]), .Y(n1785) );
  AND2X1_LVT U2657 ( .A1(I2[62]), .A2(I1[6]), .Y(n1784) );
  AND2X1_LVT U2658 ( .A1(n2583), .A2(I1[6]), .Y(n1783) );
  NAND2X0_LVT U2659 ( .A1(I2[64]), .A2(I1[6]), .Y(n1782) );
  AND2X1_LVT U2660 ( .A1(I2[0]), .A2(I1[7]), .Y(n1781) );
  AND2X1_LVT U2661 ( .A1(I2[1]), .A2(I1[7]), .Y(n1780) );
  AND2X1_LVT U2662 ( .A1(I2[2]), .A2(I1[7]), .Y(n1779) );
  AND2X1_LVT U2663 ( .A1(I2[3]), .A2(I1[7]), .Y(n1778) );
  AND2X1_LVT U2664 ( .A1(n2557), .A2(n2585), .Y(n1777) );
  AND2X1_LVT U2665 ( .A1(I2[5]), .A2(n2585), .Y(n1776) );
  AND2X1_LVT U2666 ( .A1(n2558), .A2(n2585), .Y(n1775) );
  AND2X1_LVT U2667 ( .A1(n2559), .A2(n2585), .Y(n1774) );
  AND2X1_LVT U2668 ( .A1(I2[8]), .A2(n2585), .Y(n1773) );
  AND2X1_LVT U2669 ( .A1(n2560), .A2(n2585), .Y(n1772) );
  AND2X1_LVT U2670 ( .A1(I2[10]), .A2(n2585), .Y(n1771) );
  AND2X1_LVT U2671 ( .A1(I2[11]), .A2(n2585), .Y(n1770) );
  AND2X1_LVT U2672 ( .A1(n2561), .A2(I1[7]), .Y(n1769) );
  AND2X1_LVT U2673 ( .A1(n2562), .A2(n2585), .Y(n1768) );
  AND2X1_LVT U2674 ( .A1(n2563), .A2(n2585), .Y(n1767) );
  AND2X1_LVT U2675 ( .A1(I2[15]), .A2(n2585), .Y(n1766) );
  AND2X1_LVT U2676 ( .A1(I2[16]), .A2(n2585), .Y(n1765) );
  AND2X1_LVT U2677 ( .A1(I2[17]), .A2(I1[7]), .Y(n1764) );
  AND2X1_LVT U2678 ( .A1(I2[18]), .A2(n2585), .Y(n1763) );
  AND2X1_LVT U2679 ( .A1(I2[19]), .A2(n2585), .Y(n1762) );
  AND2X1_LVT U2680 ( .A1(n2564), .A2(I1[7]), .Y(n1761) );
  AND2X1_LVT U2681 ( .A1(I2[21]), .A2(n2585), .Y(n1760) );
  AND2X1_LVT U2682 ( .A1(n2565), .A2(I1[7]), .Y(n1759) );
  AND2X1_LVT U2683 ( .A1(I2[23]), .A2(I1[7]), .Y(n1758) );
  AND2X1_LVT U2684 ( .A1(I2[24]), .A2(n2585), .Y(n1757) );
  AND2X1_LVT U2685 ( .A1(I2[25]), .A2(n2585), .Y(n1756) );
  AND2X1_LVT U2686 ( .A1(I2[26]), .A2(n2585), .Y(n1755) );
  AND2X1_LVT U2687 ( .A1(I2[27]), .A2(n2585), .Y(n1754) );
  AND2X1_LVT U2688 ( .A1(n2566), .A2(n2585), .Y(n1753) );
  AND2X1_LVT U2689 ( .A1(I2[29]), .A2(n2585), .Y(n1752) );
  AND2X1_LVT U2690 ( .A1(n2567), .A2(n2585), .Y(n1751) );
  AND2X1_LVT U2691 ( .A1(n2568), .A2(n2585), .Y(n1750) );
  AND2X1_LVT U2692 ( .A1(I2[32]), .A2(n2585), .Y(n1749) );
  AND2X1_LVT U2693 ( .A1(I2[33]), .A2(n2585), .Y(n1748) );
  AND2X1_LVT U2694 ( .A1(I2[34]), .A2(n2585), .Y(n1747) );
  AND2X1_LVT U2695 ( .A1(I2[35]), .A2(n2585), .Y(n1746) );
  AND2X1_LVT U2696 ( .A1(n2569), .A2(n2585), .Y(n1745) );
  AND2X1_LVT U2697 ( .A1(n2570), .A2(n2585), .Y(n1744) );
  AND2X1_LVT U2698 ( .A1(n2571), .A2(n2585), .Y(n1743) );
  AND2X1_LVT U2699 ( .A1(I2[39]), .A2(n2585), .Y(n1742) );
  AND2X1_LVT U2700 ( .A1(I2[40]), .A2(n2585), .Y(n1741) );
  AND2X1_LVT U2701 ( .A1(I2[41]), .A2(n2585), .Y(n1740) );
  AND2X1_LVT U2702 ( .A1(I2[42]), .A2(n2585), .Y(n1739) );
  AND2X1_LVT U2703 ( .A1(I2[43]), .A2(n2585), .Y(n1738) );
  AND2X1_LVT U2704 ( .A1(n2572), .A2(n2585), .Y(n1737) );
  AND2X1_LVT U2705 ( .A1(n2573), .A2(n2585), .Y(n1736) );
  AND2X1_LVT U2706 ( .A1(n2574), .A2(n2585), .Y(n1735) );
  AND2X1_LVT U2707 ( .A1(I2[47]), .A2(n2585), .Y(n1734) );
  AND2X1_LVT U2708 ( .A1(I2[48]), .A2(n2585), .Y(n1733) );
  AND2X1_LVT U2709 ( .A1(I2[49]), .A2(n2585), .Y(n1732) );
  AND2X1_LVT U2710 ( .A1(I2[50]), .A2(n2585), .Y(n1731) );
  AND2X1_LVT U2711 ( .A1(I2[51]), .A2(n2585), .Y(n1730) );
  AND2X1_LVT U2712 ( .A1(n2575), .A2(n2585), .Y(n1729) );
  AND2X1_LVT U2713 ( .A1(n2576), .A2(n2585), .Y(n1728) );
  AND2X1_LVT U2714 ( .A1(n2577), .A2(n2585), .Y(n1727) );
  AND2X1_LVT U2715 ( .A1(n2578), .A2(n2585), .Y(n1726) );
  AND2X1_LVT U2716 ( .A1(n2579), .A2(n2585), .Y(n1725) );
  AND2X1_LVT U2717 ( .A1(n2580), .A2(n2585), .Y(n1724) );
  AND2X1_LVT U2718 ( .A1(I2[58]), .A2(n2585), .Y(n1723) );
  AND2X1_LVT U2719 ( .A1(I2[59]), .A2(n2585), .Y(n1722) );
  AND2X1_LVT U2720 ( .A1(n2581), .A2(n2585), .Y(n1721) );
  AND2X1_LVT U2721 ( .A1(n2582), .A2(n2585), .Y(n1720) );
  AND2X1_LVT U2722 ( .A1(I2[62]), .A2(n2585), .Y(n1719) );
  AND2X1_LVT U2723 ( .A1(n2583), .A2(n2585), .Y(n1718) );
  NAND2X0_LVT U2724 ( .A1(I2[64]), .A2(n2585), .Y(n1717) );
  NAND2X0_LVT U2725 ( .A1(I1[8]), .A2(I2[1]), .Y(n1715) );
  NAND2X0_LVT U2726 ( .A1(I1[8]), .A2(I2[2]), .Y(n1714) );
  NAND2X0_LVT U2727 ( .A1(I1[8]), .A2(I2[3]), .Y(n1713) );
  NAND2X0_LVT U2728 ( .A1(I1[8]), .A2(n2557), .Y(n1712) );
  NAND2X0_LVT U2729 ( .A1(I1[8]), .A2(I2[5]), .Y(n1711) );
  NAND2X0_LVT U2730 ( .A1(I1[8]), .A2(n2558), .Y(n1710) );
  NAND2X0_LVT U2731 ( .A1(I1[8]), .A2(n2559), .Y(n1709) );
  NAND2X0_LVT U2732 ( .A1(I1[8]), .A2(I2[8]), .Y(n1708) );
  NAND2X0_LVT U2733 ( .A1(I1[8]), .A2(n2560), .Y(n1707) );
  NAND2X0_LVT U2734 ( .A1(I1[8]), .A2(I2[10]), .Y(n1706) );
  NAND2X0_LVT U2735 ( .A1(I1[8]), .A2(I2[11]), .Y(n1705) );
  NAND2X0_LVT U2736 ( .A1(I1[8]), .A2(n2561), .Y(n1704) );
  NAND2X0_LVT U2737 ( .A1(I1[8]), .A2(n2562), .Y(n1703) );
  NAND2X0_LVT U2738 ( .A1(I1[8]), .A2(n2563), .Y(n1702) );
  NAND2X0_LVT U2739 ( .A1(I1[8]), .A2(I2[15]), .Y(n1701) );
  NAND2X0_LVT U2740 ( .A1(I1[8]), .A2(I2[16]), .Y(n1700) );
  NAND2X0_LVT U2741 ( .A1(I1[8]), .A2(I2[17]), .Y(n1699) );
  NAND2X0_LVT U2742 ( .A1(I1[8]), .A2(I2[18]), .Y(n1698) );
  NAND2X0_LVT U2743 ( .A1(I1[8]), .A2(I2[19]), .Y(n1697) );
  NAND2X0_LVT U2744 ( .A1(I1[8]), .A2(n2564), .Y(n1696) );
  NAND2X0_LVT U2745 ( .A1(I1[8]), .A2(I2[21]), .Y(n1695) );
  NAND2X0_LVT U2746 ( .A1(I1[8]), .A2(n2565), .Y(n1694) );
  NAND2X0_LVT U2747 ( .A1(I1[8]), .A2(I2[23]), .Y(n1693) );
  NAND2X0_LVT U2748 ( .A1(I1[8]), .A2(I2[24]), .Y(n1692) );
  NAND2X0_LVT U2749 ( .A1(I1[8]), .A2(I2[25]), .Y(n1691) );
  NAND2X0_LVT U2750 ( .A1(I1[8]), .A2(I2[26]), .Y(n1690) );
  NAND2X0_LVT U2751 ( .A1(I1[8]), .A2(I2[27]), .Y(n1689) );
  NAND2X0_LVT U2752 ( .A1(I1[8]), .A2(n2566), .Y(n1688) );
  NAND2X0_LVT U2753 ( .A1(I1[8]), .A2(I2[29]), .Y(n1687) );
  NAND2X0_LVT U2754 ( .A1(I1[8]), .A2(n2567), .Y(n1686) );
  NAND2X0_LVT U2755 ( .A1(I1[8]), .A2(n2568), .Y(n1685) );
  NAND2X0_LVT U2756 ( .A1(I1[8]), .A2(I2[32]), .Y(n1684) );
  NAND2X0_LVT U2757 ( .A1(I1[8]), .A2(I2[33]), .Y(n1683) );
  NAND2X0_LVT U2758 ( .A1(I1[8]), .A2(I2[34]), .Y(n1682) );
  NAND2X0_LVT U2759 ( .A1(I1[8]), .A2(I2[35]), .Y(n1681) );
  NAND2X0_LVT U2760 ( .A1(I1[8]), .A2(n2569), .Y(n1680) );
  NAND2X0_LVT U2761 ( .A1(I1[8]), .A2(n2570), .Y(n1679) );
  NAND2X0_LVT U2762 ( .A1(I1[8]), .A2(n2571), .Y(n1678) );
  NAND2X0_LVT U2763 ( .A1(I1[8]), .A2(I2[39]), .Y(n1677) );
  NAND2X0_LVT U2764 ( .A1(I1[8]), .A2(I2[40]), .Y(n1676) );
  NAND2X0_LVT U2765 ( .A1(I1[8]), .A2(I2[41]), .Y(n1675) );
  NAND2X0_LVT U2766 ( .A1(I1[8]), .A2(I2[42]), .Y(n1674) );
  NAND2X0_LVT U2767 ( .A1(I1[8]), .A2(I2[43]), .Y(n1673) );
  NAND2X0_LVT U2768 ( .A1(I1[8]), .A2(n2572), .Y(n1672) );
  NAND2X0_LVT U2769 ( .A1(I1[8]), .A2(n2573), .Y(n1671) );
  NAND2X0_LVT U2770 ( .A1(I1[8]), .A2(n2574), .Y(n1670) );
  NAND2X0_LVT U2771 ( .A1(I1[8]), .A2(I2[47]), .Y(n1669) );
  NAND2X0_LVT U2772 ( .A1(I1[8]), .A2(I2[48]), .Y(n1668) );
  NAND2X0_LVT U2773 ( .A1(I1[8]), .A2(I2[49]), .Y(n1667) );
  NAND2X0_LVT U2774 ( .A1(I1[8]), .A2(I2[50]), .Y(n1666) );
  NAND2X0_LVT U2775 ( .A1(I1[8]), .A2(I2[51]), .Y(n1665) );
  NAND2X0_LVT U2776 ( .A1(I1[8]), .A2(n2575), .Y(n1664) );
  NAND2X0_LVT U2777 ( .A1(I1[8]), .A2(n2576), .Y(n1663) );
  NAND2X0_LVT U2778 ( .A1(I1[8]), .A2(n2577), .Y(n1662) );
  NAND2X0_LVT U2779 ( .A1(I1[8]), .A2(n2578), .Y(n1661) );
  NAND2X0_LVT U2780 ( .A1(I1[8]), .A2(n2579), .Y(n1660) );
  NAND2X0_LVT U2781 ( .A1(I1[8]), .A2(n2580), .Y(n1659) );
  NAND2X0_LVT U2782 ( .A1(I1[8]), .A2(I2[58]), .Y(n1658) );
  NAND2X0_LVT U2783 ( .A1(I1[8]), .A2(I2[59]), .Y(n1657) );
  NAND2X0_LVT U2784 ( .A1(I1[8]), .A2(n2581), .Y(n1656) );
  NAND2X0_LVT U2785 ( .A1(I1[8]), .A2(n2582), .Y(n1655) );
  NAND2X0_LVT U2786 ( .A1(I1[8]), .A2(I2[62]), .Y(n1654) );
  NAND2X0_LVT U2787 ( .A1(I1[8]), .A2(n2583), .Y(n1653) );
  HADDX1_LVT U2788 ( .A0(I3[8]), .B0(n2787), .SO(n1594) );
  NAND2X0_LVT U2789 ( .A1(n2787), .A2(n2588), .Y(n1593) );
  AND2X1_LVT U2790 ( .A1(I1[8]), .A2(I2[0]), .Y(n2787) );
endmodule


module MulDiv_DW_leftsh_J39_0 ( A, SH, B );
  input [126:0] A;
  input [5:0] SH;
  output [126:0] B;
  wire   n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038;

  AO22X1_LVT U544 ( .A1(SH[5]), .A2(n777), .A3(n704), .A4(n680), .Y(B[56]) );
  AO22X1_LVT U545 ( .A1(SH[5]), .A2(n805), .A3(n721), .A4(n680), .Y(B[48]) );
  AND2X1_LVT U546 ( .A1(n680), .A2(n821), .Y(B[12]) );
  AO22X1_LVT U547 ( .A1(SH[5]), .A2(n754), .A3(n680), .A4(n689), .Y(B[64]) );
  AO22X1_LVT U548 ( .A1(SH[5]), .A2(n701), .A3(n737), .A4(n680), .Y(B[40]) );
  AND2X1_LVT U549 ( .A1(n777), .A2(n680), .Y(B[24]) );
  AND2X1_LVT U550 ( .A1(n680), .A2(n875), .Y(B[2]) );
  AND2X1_LVT U551 ( .A1(n805), .A2(n680), .Y(B[16]) );
  AND2X1_LVT U552 ( .A1(n680), .A2(n800), .Y(B[4]) );
  AND2X1_LVT U553 ( .A1(n885), .A2(n680), .Y(B[0]) );
  AND2X1_LVT U554 ( .A1(n680), .A2(n880), .Y(B[1]) );
  AO22X1_LVT U555 ( .A1(SH[5]), .A2(n885), .A3(n754), .A4(n680), .Y(B[32]) );
  AO22X1_LVT U556 ( .A1(SH[5]), .A2(n789), .A3(n713), .A4(n680), .Y(B[52]) );
  INVX1_LVT U557 ( .A(SH[2]), .Y(n683) );
  INVX1_LVT U558 ( .A(SH[3]), .Y(n682) );
  INVX1_LVT U559 ( .A(SH[4]), .Y(n681) );
  INVX1_LVT U560 ( .A(SH[5]), .Y(n680) );
  INVX1_LVT U561 ( .A(SH[0]), .Y(n679) );
  INVX1_LVT U562 ( .A(SH[1]), .Y(n684) );
  AND2X1_LVT U563 ( .A1(n685), .A2(n680), .Y(B[9]) );
  AND2X1_LVT U564 ( .A1(SH[5]), .A2(n686), .Y(B[99]) );
  AND2X1_LVT U565 ( .A1(SH[5]), .A2(n687), .Y(B[98]) );
  AND2X1_LVT U566 ( .A1(SH[5]), .A2(n688), .Y(B[97]) );
  AND2X1_LVT U567 ( .A1(SH[5]), .A2(n689), .Y(B[96]) );
  AND2X1_LVT U568 ( .A1(SH[5]), .A2(n690), .Y(B[95]) );
  OA222X1_LVT U569 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n691), .A5(n680), 
        .A6(n692), .Y(B[94]) );
  AO22X1_LVT U570 ( .A1(SH[5]), .A2(n693), .A3(n680), .A4(n694), .Y(B[93]) );
  OA222X1_LVT U571 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n695), .A5(n680), 
        .A6(n696), .Y(B[92]) );
  OA222X1_LVT U572 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n697), .A5(n680), 
        .A6(n698), .Y(B[91]) );
  AO22X1_LVT U573 ( .A1(SH[5]), .A2(n699), .A3(n680), .A4(n700), .Y(B[90]) );
  AND2X1_LVT U574 ( .A1(n701), .A2(n680), .Y(B[8]) );
  AO22X1_LVT U575 ( .A1(SH[5]), .A2(n702), .A3(n680), .A4(n703), .Y(B[89]) );
  AO22X1_LVT U576 ( .A1(SH[5]), .A2(n704), .A3(n680), .A4(n705), .Y(B[88]) );
  AO22X1_LVT U577 ( .A1(SH[5]), .A2(n706), .A3(n680), .A4(n707), .Y(B[87]) );
  OA222X1_LVT U578 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n708), .A5(n680), 
        .A6(n709), .Y(B[86]) );
  OA222X1_LVT U579 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n710), .A5(n680), 
        .A6(n711), .Y(B[85]) );
  OA222X1_LVT U580 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n712), .A5(n680), 
        .A6(n713), .Y(B[84]) );
  OA222X1_LVT U581 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n714), .A5(n680), 
        .A6(n715), .Y(B[83]) );
  OA222X1_LVT U582 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n716), .A5(n680), 
        .A6(n717), .Y(B[82]) );
  OA222X1_LVT U583 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n718), .A5(n680), 
        .A6(n719), .Y(B[81]) );
  OA222X1_LVT U584 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n720), .A5(n680), 
        .A6(n721), .Y(B[80]) );
  AND2X1_LVT U585 ( .A1(n722), .A2(n680), .Y(B[7]) );
  OA222X1_LVT U586 ( .A1(SH[5]), .A2(SH[4]), .A3(SH[5]), .A4(n723), .A5(n680), 
        .A6(n724), .Y(B[79]) );
  AO22X1_LVT U587 ( .A1(SH[5]), .A2(n725), .A3(n680), .A4(n726), .Y(B[78]) );
  AO22X1_LVT U588 ( .A1(SH[5]), .A2(n727), .A3(n680), .A4(n728), .Y(B[77]) );
  AO22X1_LVT U589 ( .A1(SH[5]), .A2(n729), .A3(n680), .A4(n730), .Y(B[76]) );
  AO22X1_LVT U590 ( .A1(SH[5]), .A2(n731), .A3(n680), .A4(n732), .Y(B[75]) );
  AO22X1_LVT U591 ( .A1(SH[5]), .A2(n733), .A3(n680), .A4(n734), .Y(B[74]) );
  AO22X1_LVT U592 ( .A1(SH[5]), .A2(n735), .A3(n680), .A4(n736), .Y(B[73]) );
  AO22X1_LVT U593 ( .A1(SH[5]), .A2(n737), .A3(n680), .A4(n738), .Y(B[72]) );
  AO22X1_LVT U594 ( .A1(SH[5]), .A2(n739), .A3(n680), .A4(n740), .Y(B[71]) );
  AO22X1_LVT U595 ( .A1(SH[5]), .A2(n741), .A3(n680), .A4(n742), .Y(B[70]) );
  AND2X1_LVT U596 ( .A1(n743), .A2(n680), .Y(B[6]) );
  AO22X1_LVT U597 ( .A1(SH[5]), .A2(n744), .A3(n680), .A4(n745), .Y(B[69]) );
  AO22X1_LVT U598 ( .A1(SH[5]), .A2(n746), .A3(n680), .A4(n747), .Y(B[68]) );
  AO22X1_LVT U599 ( .A1(SH[5]), .A2(n748), .A3(n680), .A4(n686), .Y(B[67]) );
  AO22X1_LVT U600 ( .A1(SH[4]), .A2(n749), .A3(n681), .A4(n714), .Y(n686) );
  AO22X1_LVT U601 ( .A1(SH[5]), .A2(n750), .A3(n680), .A4(n687), .Y(B[66]) );
  AO22X1_LVT U602 ( .A1(SH[4]), .A2(n751), .A3(n681), .A4(n716), .Y(n687) );
  AO22X1_LVT U603 ( .A1(SH[5]), .A2(n752), .A3(n680), .A4(n688), .Y(B[65]) );
  AO22X1_LVT U604 ( .A1(SH[4]), .A2(n753), .A3(n681), .A4(n718), .Y(n688) );
  AO22X1_LVT U605 ( .A1(SH[4]), .A2(n755), .A3(n681), .A4(n720), .Y(n689) );
  AO22X1_LVT U606 ( .A1(SH[5]), .A2(n756), .A3(n680), .A4(n690), .Y(B[63]) );
  AO22X1_LVT U607 ( .A1(SH[4]), .A2(n757), .A3(n681), .A4(n723), .Y(n690) );
  AO22X1_LVT U608 ( .A1(SH[5]), .A2(n758), .A3(n680), .A4(n692), .Y(B[62]) );
  AO22X1_LVT U609 ( .A1(SH[4]), .A2(n759), .A3(n681), .A4(n760), .Y(n692) );
  AO22X1_LVT U610 ( .A1(SH[5]), .A2(n761), .A3(n680), .A4(n693), .Y(B[61]) );
  AO22X1_LVT U611 ( .A1(SH[4]), .A2(n762), .A3(n681), .A4(n763), .Y(n693) );
  AO22X1_LVT U612 ( .A1(SH[5]), .A2(n764), .A3(n680), .A4(n696), .Y(B[60]) );
  AO22X1_LVT U613 ( .A1(SH[4]), .A2(n765), .A3(n681), .A4(n766), .Y(n696) );
  AND2X1_LVT U614 ( .A1(n767), .A2(n680), .Y(B[5]) );
  AO22X1_LVT U615 ( .A1(SH[5]), .A2(n768), .A3(n680), .A4(n698), .Y(B[59]) );
  AO22X1_LVT U616 ( .A1(SH[4]), .A2(n769), .A3(n681), .A4(n770), .Y(n698) );
  AO22X1_LVT U617 ( .A1(SH[5]), .A2(n771), .A3(n680), .A4(n699), .Y(B[58]) );
  AO22X1_LVT U618 ( .A1(SH[4]), .A2(n772), .A3(n681), .A4(n773), .Y(n699) );
  AO22X1_LVT U619 ( .A1(SH[5]), .A2(n774), .A3(n680), .A4(n702), .Y(B[57]) );
  AO22X1_LVT U620 ( .A1(SH[4]), .A2(n775), .A3(n681), .A4(n776), .Y(n702) );
  AO22X1_LVT U621 ( .A1(SH[4]), .A2(n778), .A3(n681), .A4(n779), .Y(n704) );
  AO22X1_LVT U622 ( .A1(SH[5]), .A2(n780), .A3(n680), .A4(n706), .Y(B[55]) );
  AO22X1_LVT U623 ( .A1(SH[4]), .A2(n781), .A3(n681), .A4(n782), .Y(n706) );
  AO22X1_LVT U624 ( .A1(SH[5]), .A2(n783), .A3(n680), .A4(n709), .Y(B[54]) );
  AO22X1_LVT U625 ( .A1(SH[4]), .A2(n784), .A3(n681), .A4(n785), .Y(n709) );
  AO22X1_LVT U626 ( .A1(SH[5]), .A2(n786), .A3(n680), .A4(n711), .Y(B[53]) );
  AO22X1_LVT U627 ( .A1(SH[4]), .A2(n787), .A3(n681), .A4(n788), .Y(n711) );
  AO22X1_LVT U628 ( .A1(SH[4]), .A2(n790), .A3(n681), .A4(n791), .Y(n713) );
  AO22X1_LVT U629 ( .A1(SH[5]), .A2(n792), .A3(n680), .A4(n715), .Y(B[51]) );
  AO22X1_LVT U630 ( .A1(SH[4]), .A2(n793), .A3(n681), .A4(n749), .Y(n715) );
  AO22X1_LVT U631 ( .A1(SH[3]), .A2(n794), .A3(n682), .A4(n795), .Y(n749) );
  AO22X1_LVT U632 ( .A1(SH[5]), .A2(n796), .A3(n680), .A4(n717), .Y(B[50]) );
  AO22X1_LVT U633 ( .A1(SH[4]), .A2(n797), .A3(n681), .A4(n751), .Y(n717) );
  AO22X1_LVT U634 ( .A1(SH[3]), .A2(n798), .A3(n682), .A4(n799), .Y(n751) );
  AO22X1_LVT U635 ( .A1(SH[5]), .A2(n801), .A3(n680), .A4(n719), .Y(B[49]) );
  AO22X1_LVT U636 ( .A1(SH[4]), .A2(n802), .A3(n681), .A4(n753), .Y(n719) );
  AO22X1_LVT U637 ( .A1(SH[3]), .A2(n803), .A3(n682), .A4(n804), .Y(n753) );
  AO22X1_LVT U638 ( .A1(SH[4]), .A2(n806), .A3(n681), .A4(n755), .Y(n721) );
  AO22X1_LVT U639 ( .A1(SH[3]), .A2(n807), .A3(n682), .A4(n808), .Y(n755) );
  AO22X1_LVT U640 ( .A1(SH[5]), .A2(n809), .A3(n680), .A4(n724), .Y(B[47]) );
  AO22X1_LVT U641 ( .A1(SH[4]), .A2(n810), .A3(n681), .A4(n757), .Y(n724) );
  AO22X1_LVT U642 ( .A1(SH[3]), .A2(n811), .A3(n682), .A4(n812), .Y(n757) );
  AO22X1_LVT U643 ( .A1(SH[5]), .A2(n813), .A3(n680), .A4(n725), .Y(B[46]) );
  AO22X1_LVT U644 ( .A1(SH[4]), .A2(n814), .A3(n681), .A4(n759), .Y(n725) );
  AO22X1_LVT U645 ( .A1(SH[3]), .A2(n815), .A3(n682), .A4(n816), .Y(n759) );
  AO22X1_LVT U646 ( .A1(SH[5]), .A2(n817), .A3(n680), .A4(n727), .Y(B[45]) );
  AO22X1_LVT U647 ( .A1(SH[4]), .A2(n818), .A3(n681), .A4(n762), .Y(n727) );
  AO22X1_LVT U648 ( .A1(SH[3]), .A2(n819), .A3(n682), .A4(n820), .Y(n762) );
  AO22X1_LVT U649 ( .A1(SH[5]), .A2(n821), .A3(n680), .A4(n729), .Y(B[44]) );
  AO22X1_LVT U650 ( .A1(SH[4]), .A2(n822), .A3(n681), .A4(n765), .Y(n729) );
  AO22X1_LVT U651 ( .A1(SH[3]), .A2(n823), .A3(n682), .A4(n824), .Y(n765) );
  AO22X1_LVT U652 ( .A1(SH[5]), .A2(n825), .A3(n680), .A4(n731), .Y(B[43]) );
  AO22X1_LVT U653 ( .A1(SH[4]), .A2(n826), .A3(n681), .A4(n769), .Y(n731) );
  AO22X1_LVT U654 ( .A1(SH[3]), .A2(n827), .A3(n682), .A4(n794), .Y(n769) );
  AO22X1_LVT U655 ( .A1(SH[2]), .A2(n828), .A3(n683), .A4(n829), .Y(n794) );
  AO22X1_LVT U656 ( .A1(SH[5]), .A2(n830), .A3(n680), .A4(n733), .Y(B[42]) );
  AO22X1_LVT U657 ( .A1(SH[4]), .A2(n831), .A3(n681), .A4(n772), .Y(n733) );
  AO22X1_LVT U658 ( .A1(SH[3]), .A2(n832), .A3(n682), .A4(n798), .Y(n772) );
  AO22X1_LVT U659 ( .A1(SH[2]), .A2(n833), .A3(n683), .A4(n834), .Y(n798) );
  AO22X1_LVT U660 ( .A1(SH[5]), .A2(n685), .A3(n680), .A4(n735), .Y(B[41]) );
  AO22X1_LVT U661 ( .A1(SH[4]), .A2(n835), .A3(n681), .A4(n775), .Y(n735) );
  AO22X1_LVT U662 ( .A1(SH[3]), .A2(n836), .A3(n682), .A4(n803), .Y(n775) );
  AO22X1_LVT U663 ( .A1(SH[2]), .A2(n837), .A3(n683), .A4(n838), .Y(n803) );
  OA221X1_LVT U664 ( .A1(SH[3]), .A2(n839), .A3(n682), .A4(n840), .A5(n681), 
        .Y(n685) );
  AO22X1_LVT U665 ( .A1(SH[4]), .A2(n841), .A3(n681), .A4(n778), .Y(n737) );
  AO22X1_LVT U666 ( .A1(SH[3]), .A2(n842), .A3(n682), .A4(n807), .Y(n778) );
  AO22X1_LVT U667 ( .A1(SH[2]), .A2(n843), .A3(n683), .A4(n844), .Y(n807) );
  OA221X1_LVT U668 ( .A1(SH[3]), .A2(n845), .A3(n682), .A4(n846), .A5(n681), 
        .Y(n701) );
  AND2X1_LVT U669 ( .A1(n847), .A2(n680), .Y(B[3]) );
  AO22X1_LVT U670 ( .A1(SH[5]), .A2(n722), .A3(n680), .A4(n739), .Y(B[39]) );
  AO22X1_LVT U671 ( .A1(SH[4]), .A2(n848), .A3(n681), .A4(n781), .Y(n739) );
  AO22X1_LVT U672 ( .A1(SH[3]), .A2(n849), .A3(n682), .A4(n811), .Y(n781) );
  AO22X1_LVT U673 ( .A1(SH[2]), .A2(n850), .A3(n683), .A4(n828), .Y(n811) );
  AO22X1_LVT U674 ( .A1(SH[1]), .A2(n851), .A3(n684), .A4(n852), .Y(n828) );
  AND2X1_LVT U675 ( .A1(n853), .A2(n681), .Y(n722) );
  AO22X1_LVT U676 ( .A1(SH[5]), .A2(n743), .A3(n680), .A4(n741), .Y(B[38]) );
  AO22X1_LVT U677 ( .A1(SH[4]), .A2(n854), .A3(n681), .A4(n784), .Y(n741) );
  AO22X1_LVT U678 ( .A1(SH[3]), .A2(n855), .A3(n682), .A4(n815), .Y(n784) );
  AO22X1_LVT U679 ( .A1(SH[2]), .A2(n856), .A3(n683), .A4(n833), .Y(n815) );
  AO22X1_LVT U680 ( .A1(SH[1]), .A2(n857), .A3(n684), .A4(n858), .Y(n833) );
  AND2X1_LVT U681 ( .A1(n859), .A2(n681), .Y(n743) );
  AO22X1_LVT U682 ( .A1(SH[5]), .A2(n767), .A3(n680), .A4(n744), .Y(B[37]) );
  AO22X1_LVT U683 ( .A1(SH[4]), .A2(n860), .A3(n681), .A4(n787), .Y(n744) );
  AO22X1_LVT U684 ( .A1(SH[3]), .A2(n861), .A3(n682), .A4(n819), .Y(n787) );
  AO22X1_LVT U685 ( .A1(SH[2]), .A2(n862), .A3(n683), .A4(n837), .Y(n819) );
  AO22X1_LVT U686 ( .A1(SH[1]), .A2(n863), .A3(n684), .A4(n851), .Y(n837) );
  AO22X1_LVT U687 ( .A1(SH[0]), .A2(A[36]), .A3(n679), .A4(A[37]), .Y(n851) );
  AND2X1_LVT U688 ( .A1(n864), .A2(n681), .Y(n767) );
  AO22X1_LVT U689 ( .A1(SH[5]), .A2(n800), .A3(n680), .A4(n746), .Y(B[36]) );
  AO22X1_LVT U690 ( .A1(SH[4]), .A2(n865), .A3(n681), .A4(n790), .Y(n746) );
  AO22X1_LVT U691 ( .A1(SH[3]), .A2(n866), .A3(n682), .A4(n823), .Y(n790) );
  AO22X1_LVT U692 ( .A1(SH[2]), .A2(n867), .A3(n683), .A4(n843), .Y(n823) );
  AO22X1_LVT U693 ( .A1(SH[1]), .A2(n868), .A3(n684), .A4(n857), .Y(n843) );
  AO22X1_LVT U694 ( .A1(SH[0]), .A2(A[35]), .A3(n679), .A4(A[36]), .Y(n857) );
  AND2X1_LVT U695 ( .A1(n869), .A2(n681), .Y(n800) );
  AO22X1_LVT U696 ( .A1(SH[5]), .A2(n847), .A3(n680), .A4(n748), .Y(B[35]) );
  AO22X1_LVT U697 ( .A1(SH[4]), .A2(n870), .A3(n681), .A4(n793), .Y(n748) );
  AO22X1_LVT U698 ( .A1(SH[3]), .A2(n871), .A3(n682), .A4(n827), .Y(n793) );
  AO22X1_LVT U699 ( .A1(SH[2]), .A2(n872), .A3(n683), .A4(n850), .Y(n827) );
  AO22X1_LVT U700 ( .A1(SH[1]), .A2(n873), .A3(n684), .A4(n863), .Y(n850) );
  AO22X1_LVT U701 ( .A1(SH[0]), .A2(A[34]), .A3(n679), .A4(A[35]), .Y(n863) );
  AND2X1_LVT U702 ( .A1(n874), .A2(n681), .Y(n847) );
  AO22X1_LVT U703 ( .A1(SH[5]), .A2(n875), .A3(n680), .A4(n750), .Y(B[34]) );
  AO22X1_LVT U704 ( .A1(SH[4]), .A2(n876), .A3(n681), .A4(n797), .Y(n750) );
  AO22X1_LVT U705 ( .A1(SH[3]), .A2(n877), .A3(n682), .A4(n832), .Y(n797) );
  AO22X1_LVT U706 ( .A1(SH[2]), .A2(n878), .A3(n683), .A4(n856), .Y(n832) );
  AO22X1_LVT U707 ( .A1(SH[1]), .A2(n879), .A3(n684), .A4(n868), .Y(n856) );
  AO22X1_LVT U708 ( .A1(SH[0]), .A2(A[33]), .A3(n679), .A4(A[34]), .Y(n868) );
  AO22X1_LVT U709 ( .A1(SH[5]), .A2(n880), .A3(n680), .A4(n752), .Y(B[33]) );
  AO22X1_LVT U710 ( .A1(SH[4]), .A2(n881), .A3(n681), .A4(n802), .Y(n752) );
  AO22X1_LVT U711 ( .A1(SH[3]), .A2(n882), .A3(n682), .A4(n836), .Y(n802) );
  AO22X1_LVT U712 ( .A1(SH[2]), .A2(n883), .A3(n683), .A4(n862), .Y(n836) );
  AO22X1_LVT U713 ( .A1(SH[1]), .A2(n884), .A3(n684), .A4(n873), .Y(n862) );
  AO22X1_LVT U714 ( .A1(SH[0]), .A2(A[32]), .A3(n679), .A4(A[33]), .Y(n873) );
  AO22X1_LVT U715 ( .A1(SH[4]), .A2(n886), .A3(n681), .A4(n806), .Y(n754) );
  AO22X1_LVT U716 ( .A1(SH[3]), .A2(n887), .A3(n682), .A4(n842), .Y(n806) );
  AO22X1_LVT U717 ( .A1(SH[2]), .A2(n888), .A3(n683), .A4(n867), .Y(n842) );
  AO22X1_LVT U718 ( .A1(SH[1]), .A2(n889), .A3(n684), .A4(n879), .Y(n867) );
  AO22X1_LVT U719 ( .A1(SH[0]), .A2(A[31]), .A3(n679), .A4(A[32]), .Y(n879) );
  AND2X1_LVT U720 ( .A1(n680), .A2(n756), .Y(B[31]) );
  AO22X1_LVT U721 ( .A1(SH[4]), .A2(n890), .A3(n681), .A4(n810), .Y(n756) );
  AO22X1_LVT U722 ( .A1(SH[3]), .A2(n891), .A3(n682), .A4(n849), .Y(n810) );
  AO22X1_LVT U723 ( .A1(SH[2]), .A2(n892), .A3(n683), .A4(n872), .Y(n849) );
  AO22X1_LVT U724 ( .A1(SH[1]), .A2(n893), .A3(n684), .A4(n884), .Y(n872) );
  AO22X1_LVT U725 ( .A1(SH[0]), .A2(A[30]), .A3(n679), .A4(A[31]), .Y(n884) );
  AND2X1_LVT U726 ( .A1(n680), .A2(n758), .Y(B[30]) );
  AO22X1_LVT U727 ( .A1(SH[4]), .A2(n894), .A3(n681), .A4(n814), .Y(n758) );
  AO22X1_LVT U728 ( .A1(SH[3]), .A2(n895), .A3(n682), .A4(n855), .Y(n814) );
  AO22X1_LVT U729 ( .A1(SH[2]), .A2(n896), .A3(n683), .A4(n878), .Y(n855) );
  AO22X1_LVT U730 ( .A1(SH[1]), .A2(n897), .A3(n684), .A4(n889), .Y(n878) );
  AO22X1_LVT U731 ( .A1(SH[0]), .A2(A[29]), .A3(n679), .A4(A[30]), .Y(n889) );
  AND2X1_LVT U732 ( .A1(n898), .A2(n681), .Y(n875) );
  AND2X1_LVT U733 ( .A1(n680), .A2(n761), .Y(B[29]) );
  AO22X1_LVT U734 ( .A1(SH[4]), .A2(n899), .A3(n681), .A4(n818), .Y(n761) );
  AO22X1_LVT U735 ( .A1(SH[3]), .A2(n900), .A3(n682), .A4(n861), .Y(n818) );
  AO22X1_LVT U736 ( .A1(SH[2]), .A2(n901), .A3(n683), .A4(n883), .Y(n861) );
  AO22X1_LVT U737 ( .A1(SH[1]), .A2(n902), .A3(n684), .A4(n893), .Y(n883) );
  AO22X1_LVT U738 ( .A1(SH[0]), .A2(A[28]), .A3(n679), .A4(A[29]), .Y(n893) );
  AND2X1_LVT U739 ( .A1(n680), .A2(n764), .Y(B[28]) );
  AO22X1_LVT U740 ( .A1(SH[4]), .A2(n903), .A3(n681), .A4(n822), .Y(n764) );
  AO22X1_LVT U741 ( .A1(SH[3]), .A2(n904), .A3(n682), .A4(n866), .Y(n822) );
  AO22X1_LVT U742 ( .A1(SH[2]), .A2(n905), .A3(n683), .A4(n888), .Y(n866) );
  AO22X1_LVT U743 ( .A1(SH[1]), .A2(n906), .A3(n684), .A4(n897), .Y(n888) );
  AO22X1_LVT U744 ( .A1(SH[0]), .A2(A[27]), .A3(n679), .A4(A[28]), .Y(n897) );
  AO22X1_LVT U745 ( .A1(SH[3]), .A2(n907), .A3(n682), .A4(n908), .Y(n903) );
  AND2X1_LVT U746 ( .A1(n680), .A2(n768), .Y(B[27]) );
  AO22X1_LVT U747 ( .A1(SH[4]), .A2(n909), .A3(n681), .A4(n826), .Y(n768) );
  AO22X1_LVT U748 ( .A1(SH[3]), .A2(n910), .A3(n682), .A4(n871), .Y(n826) );
  AO22X1_LVT U749 ( .A1(SH[2]), .A2(n911), .A3(n683), .A4(n892), .Y(n871) );
  AO22X1_LVT U750 ( .A1(SH[1]), .A2(n912), .A3(n684), .A4(n902), .Y(n892) );
  AO22X1_LVT U751 ( .A1(SH[0]), .A2(A[26]), .A3(n679), .A4(A[27]), .Y(n902) );
  AO22X1_LVT U752 ( .A1(SH[3]), .A2(n913), .A3(n682), .A4(n914), .Y(n909) );
  AND2X1_LVT U753 ( .A1(n680), .A2(n771), .Y(B[26]) );
  AO22X1_LVT U754 ( .A1(SH[4]), .A2(n915), .A3(n681), .A4(n831), .Y(n771) );
  AO22X1_LVT U755 ( .A1(SH[3]), .A2(n916), .A3(n682), .A4(n877), .Y(n831) );
  AO22X1_LVT U756 ( .A1(SH[2]), .A2(n917), .A3(n683), .A4(n896), .Y(n877) );
  AO22X1_LVT U757 ( .A1(SH[1]), .A2(n918), .A3(n684), .A4(n906), .Y(n896) );
  AO22X1_LVT U758 ( .A1(SH[0]), .A2(A[25]), .A3(n679), .A4(A[26]), .Y(n906) );
  AO22X1_LVT U759 ( .A1(SH[3]), .A2(n919), .A3(n682), .A4(n920), .Y(n915) );
  AND2X1_LVT U760 ( .A1(n680), .A2(n774), .Y(B[25]) );
  AO22X1_LVT U761 ( .A1(SH[4]), .A2(n921), .A3(n681), .A4(n835), .Y(n774) );
  AO22X1_LVT U762 ( .A1(SH[3]), .A2(n922), .A3(n682), .A4(n882), .Y(n835) );
  AO22X1_LVT U763 ( .A1(SH[2]), .A2(n923), .A3(n683), .A4(n901), .Y(n882) );
  AO22X1_LVT U764 ( .A1(SH[1]), .A2(n924), .A3(n684), .A4(n912), .Y(n901) );
  AO22X1_LVT U765 ( .A1(SH[0]), .A2(A[24]), .A3(n679), .A4(A[25]), .Y(n912) );
  AO22X1_LVT U766 ( .A1(SH[3]), .A2(n840), .A3(n682), .A4(n839), .Y(n921) );
  AO22X1_LVT U767 ( .A1(SH[4]), .A2(n925), .A3(n681), .A4(n841), .Y(n777) );
  AO22X1_LVT U768 ( .A1(SH[3]), .A2(n926), .A3(n682), .A4(n887), .Y(n841) );
  AO22X1_LVT U769 ( .A1(SH[2]), .A2(n927), .A3(n683), .A4(n905), .Y(n887) );
  AO22X1_LVT U770 ( .A1(SH[1]), .A2(n928), .A3(n684), .A4(n918), .Y(n905) );
  AO22X1_LVT U771 ( .A1(SH[0]), .A2(A[23]), .A3(n679), .A4(A[24]), .Y(n918) );
  AO22X1_LVT U772 ( .A1(SH[3]), .A2(n846), .A3(n682), .A4(n845), .Y(n925) );
  AND2X1_LVT U773 ( .A1(n680), .A2(n780), .Y(B[23]) );
  AO22X1_LVT U774 ( .A1(SH[4]), .A2(n853), .A3(n681), .A4(n848), .Y(n780) );
  AO22X1_LVT U775 ( .A1(SH[3]), .A2(n929), .A3(n682), .A4(n891), .Y(n848) );
  AO22X1_LVT U776 ( .A1(SH[2]), .A2(n930), .A3(n683), .A4(n911), .Y(n891) );
  AO22X1_LVT U777 ( .A1(SH[1]), .A2(n931), .A3(n684), .A4(n924), .Y(n911) );
  AO22X1_LVT U778 ( .A1(SH[0]), .A2(A[22]), .A3(n679), .A4(A[23]), .Y(n924) );
  OA221X1_LVT U779 ( .A1(SH[2]), .A2(n932), .A3(n683), .A4(n933), .A5(n682), 
        .Y(n853) );
  AND2X1_LVT U780 ( .A1(n680), .A2(n783), .Y(B[22]) );
  AO22X1_LVT U781 ( .A1(SH[4]), .A2(n859), .A3(n681), .A4(n854), .Y(n783) );
  AO22X1_LVT U782 ( .A1(SH[3]), .A2(n934), .A3(n682), .A4(n895), .Y(n854) );
  AO22X1_LVT U783 ( .A1(SH[2]), .A2(n935), .A3(n683), .A4(n917), .Y(n895) );
  AO22X1_LVT U784 ( .A1(SH[1]), .A2(n936), .A3(n684), .A4(n928), .Y(n917) );
  AO22X1_LVT U785 ( .A1(SH[0]), .A2(A[21]), .A3(n679), .A4(A[22]), .Y(n928) );
  OA221X1_LVT U786 ( .A1(SH[2]), .A2(n937), .A3(n683), .A4(n938), .A5(n682), 
        .Y(n859) );
  AND2X1_LVT U787 ( .A1(n680), .A2(n786), .Y(B[21]) );
  AO22X1_LVT U788 ( .A1(SH[4]), .A2(n864), .A3(n681), .A4(n860), .Y(n786) );
  AO22X1_LVT U789 ( .A1(SH[3]), .A2(n939), .A3(n682), .A4(n900), .Y(n860) );
  AO22X1_LVT U790 ( .A1(SH[2]), .A2(n940), .A3(n683), .A4(n923), .Y(n900) );
  AO22X1_LVT U791 ( .A1(SH[1]), .A2(n941), .A3(n684), .A4(n931), .Y(n923) );
  AO22X1_LVT U792 ( .A1(SH[0]), .A2(A[20]), .A3(n679), .A4(A[21]), .Y(n931) );
  OA221X1_LVT U793 ( .A1(SH[2]), .A2(n942), .A3(n683), .A4(n943), .A5(n682), 
        .Y(n864) );
  AND2X1_LVT U794 ( .A1(n680), .A2(n789), .Y(B[20]) );
  AO22X1_LVT U795 ( .A1(SH[4]), .A2(n869), .A3(n681), .A4(n865), .Y(n789) );
  AO22X1_LVT U796 ( .A1(SH[3]), .A2(n908), .A3(n682), .A4(n904), .Y(n865) );
  AO22X1_LVT U797 ( .A1(SH[2]), .A2(n944), .A3(n683), .A4(n927), .Y(n904) );
  AO22X1_LVT U798 ( .A1(SH[1]), .A2(n945), .A3(n684), .A4(n936), .Y(n927) );
  AO22X1_LVT U799 ( .A1(SH[0]), .A2(A[19]), .A3(n679), .A4(A[20]), .Y(n936) );
  AND2X1_LVT U800 ( .A1(n682), .A2(n907), .Y(n869) );
  AND2X1_LVT U801 ( .A1(n946), .A2(n681), .Y(n880) );
  AND2X1_LVT U802 ( .A1(n680), .A2(n792), .Y(B[19]) );
  AO22X1_LVT U803 ( .A1(SH[4]), .A2(n874), .A3(n681), .A4(n870), .Y(n792) );
  AO22X1_LVT U804 ( .A1(SH[3]), .A2(n914), .A3(n682), .A4(n910), .Y(n870) );
  AO22X1_LVT U805 ( .A1(SH[2]), .A2(n947), .A3(n683), .A4(n930), .Y(n910) );
  AO22X1_LVT U806 ( .A1(SH[1]), .A2(n948), .A3(n684), .A4(n941), .Y(n930) );
  AO22X1_LVT U807 ( .A1(SH[0]), .A2(A[18]), .A3(n679), .A4(A[19]), .Y(n941) );
  AND2X1_LVT U808 ( .A1(n913), .A2(n682), .Y(n874) );
  AND2X1_LVT U809 ( .A1(n680), .A2(n796), .Y(B[18]) );
  AO22X1_LVT U810 ( .A1(SH[4]), .A2(n898), .A3(n681), .A4(n876), .Y(n796) );
  AO22X1_LVT U811 ( .A1(SH[3]), .A2(n920), .A3(n682), .A4(n916), .Y(n876) );
  AO22X1_LVT U812 ( .A1(SH[2]), .A2(n949), .A3(n683), .A4(n935), .Y(n916) );
  AO22X1_LVT U813 ( .A1(SH[1]), .A2(n950), .A3(n684), .A4(n945), .Y(n935) );
  AO22X1_LVT U814 ( .A1(SH[0]), .A2(A[17]), .A3(n679), .A4(A[18]), .Y(n945) );
  AND2X1_LVT U815 ( .A1(n919), .A2(n682), .Y(n898) );
  AND2X1_LVT U816 ( .A1(n680), .A2(n801), .Y(B[17]) );
  AO22X1_LVT U817 ( .A1(SH[4]), .A2(n946), .A3(n681), .A4(n881), .Y(n801) );
  AO22X1_LVT U818 ( .A1(SH[3]), .A2(n839), .A3(n682), .A4(n922), .Y(n881) );
  AO22X1_LVT U819 ( .A1(SH[2]), .A2(n951), .A3(n683), .A4(n940), .Y(n922) );
  AO22X1_LVT U820 ( .A1(SH[1]), .A2(n952), .A3(n684), .A4(n948), .Y(n940) );
  AO22X1_LVT U821 ( .A1(SH[0]), .A2(A[16]), .A3(n679), .A4(A[17]), .Y(n948) );
  AO22X1_LVT U822 ( .A1(SH[2]), .A2(n942), .A3(n683), .A4(n953), .Y(n839) );
  AND2X1_LVT U823 ( .A1(n840), .A2(n682), .Y(n946) );
  AND2X1_LVT U824 ( .A1(n943), .A2(n683), .Y(n840) );
  OA222X1_LVT U825 ( .A1(n681), .A2(n846), .A3(n681), .A4(n682), .A5(SH[4]), 
        .A6(n886), .Y(n805) );
  AO22X1_LVT U826 ( .A1(SH[3]), .A2(n845), .A3(n682), .A4(n926), .Y(n886) );
  AO22X1_LVT U827 ( .A1(SH[2]), .A2(n954), .A3(n683), .A4(n944), .Y(n926) );
  AO22X1_LVT U828 ( .A1(SH[1]), .A2(n955), .A3(n684), .A4(n950), .Y(n944) );
  AO22X1_LVT U829 ( .A1(SH[0]), .A2(A[15]), .A3(n679), .A4(A[16]), .Y(n950) );
  AO22X1_LVT U830 ( .A1(SH[2]), .A2(n956), .A3(n683), .A4(n957), .Y(n845) );
  AND2X1_LVT U831 ( .A1(n809), .A2(n680), .Y(B[15]) );
  AND2X1_LVT U832 ( .A1(n681), .A2(n890), .Y(n809) );
  AO22X1_LVT U833 ( .A1(SH[3]), .A2(n958), .A3(n682), .A4(n929), .Y(n890) );
  AO22X1_LVT U834 ( .A1(SH[2]), .A2(n959), .A3(n683), .A4(n947), .Y(n929) );
  AO22X1_LVT U835 ( .A1(SH[1]), .A2(n960), .A3(n684), .A4(n952), .Y(n947) );
  AO22X1_LVT U836 ( .A1(SH[0]), .A2(A[14]), .A3(n679), .A4(A[15]), .Y(n952) );
  AO22X1_LVT U837 ( .A1(SH[2]), .A2(n933), .A3(n683), .A4(n932), .Y(n958) );
  AND2X1_LVT U838 ( .A1(n813), .A2(n680), .Y(B[14]) );
  AND2X1_LVT U839 ( .A1(n681), .A2(n894), .Y(n813) );
  AO22X1_LVT U840 ( .A1(SH[3]), .A2(n961), .A3(n682), .A4(n934), .Y(n894) );
  AO22X1_LVT U841 ( .A1(SH[2]), .A2(n962), .A3(n683), .A4(n949), .Y(n934) );
  AO22X1_LVT U842 ( .A1(SH[1]), .A2(n963), .A3(n684), .A4(n955), .Y(n949) );
  AO22X1_LVT U843 ( .A1(SH[0]), .A2(A[13]), .A3(n679), .A4(A[14]), .Y(n955) );
  AO22X1_LVT U844 ( .A1(SH[2]), .A2(n938), .A3(n683), .A4(n937), .Y(n961) );
  AND2X1_LVT U845 ( .A1(n817), .A2(n680), .Y(B[13]) );
  AND2X1_LVT U846 ( .A1(n681), .A2(n899), .Y(n817) );
  AO22X1_LVT U847 ( .A1(SH[3]), .A2(n964), .A3(n682), .A4(n939), .Y(n899) );
  AO22X1_LVT U848 ( .A1(SH[2]), .A2(n953), .A3(n683), .A4(n951), .Y(n939) );
  AO22X1_LVT U849 ( .A1(SH[1]), .A2(n965), .A3(n684), .A4(n960), .Y(n951) );
  AO22X1_LVT U850 ( .A1(SH[0]), .A2(A[12]), .A3(n679), .A4(A[13]), .Y(n960) );
  AO22X1_LVT U851 ( .A1(SH[1]), .A2(n966), .A3(n684), .A4(n967), .Y(n953) );
  AO22X1_LVT U852 ( .A1(SH[2]), .A2(n943), .A3(n683), .A4(n942), .Y(n964) );
  AO22X1_LVT U853 ( .A1(SH[1]), .A2(n968), .A3(n684), .A4(n969), .Y(n942) );
  OA221X1_LVT U854 ( .A1(SH[0]), .A2(A[1]), .A3(n679), .A4(A[0]), .A5(n684), 
        .Y(n943) );
  OA221X1_LVT U855 ( .A1(SH[3]), .A2(n908), .A3(n682), .A4(n907), .A5(n681), 
        .Y(n821) );
  AO22X1_LVT U856 ( .A1(SH[2]), .A2(n970), .A3(n683), .A4(n956), .Y(n907) );
  AO22X1_LVT U857 ( .A1(SH[1]), .A2(n971), .A3(n684), .A4(n972), .Y(n956) );
  AND3X1_LVT U858 ( .A1(A[0]), .A2(n684), .A3(n679), .Y(n970) );
  AO22X1_LVT U859 ( .A1(SH[2]), .A2(n957), .A3(n683), .A4(n954), .Y(n908) );
  AO22X1_LVT U860 ( .A1(SH[1]), .A2(n973), .A3(n684), .A4(n963), .Y(n954) );
  AO22X1_LVT U861 ( .A1(SH[0]), .A2(A[11]), .A3(n679), .A4(A[12]), .Y(n963) );
  AO22X1_LVT U862 ( .A1(SH[1]), .A2(n974), .A3(n684), .A4(n975), .Y(n957) );
  AND3X1_LVT U863 ( .A1(SH[5]), .A2(SH[4]), .A3(n691), .Y(B[126]) );
  AND2X1_LVT U864 ( .A1(SH[5]), .A2(n694), .Y(B[125]) );
  AND3X1_LVT U865 ( .A1(SH[4]), .A2(SH[3]), .A3(n976), .Y(n694) );
  AND3X1_LVT U866 ( .A1(SH[5]), .A2(SH[4]), .A3(n695), .Y(B[124]) );
  AND3X1_LVT U867 ( .A1(SH[5]), .A2(SH[4]), .A3(n697), .Y(B[123]) );
  AND2X1_LVT U868 ( .A1(SH[5]), .A2(n700), .Y(B[122]) );
  AND3X1_LVT U869 ( .A1(SH[3]), .A2(SH[4]), .A3(n977), .Y(n700) );
  AND2X1_LVT U870 ( .A1(SH[5]), .A2(n703), .Y(B[121]) );
  AND3X1_LVT U871 ( .A1(SH[3]), .A2(SH[4]), .A3(n978), .Y(n703) );
  AND2X1_LVT U872 ( .A1(SH[5]), .A2(n705), .Y(B[120]) );
  AND3X1_LVT U873 ( .A1(SH[3]), .A2(SH[4]), .A3(n979), .Y(n705) );
  AND2X1_LVT U874 ( .A1(n825), .A2(n680), .Y(B[11]) );
  OA221X1_LVT U875 ( .A1(SH[3]), .A2(n914), .A3(n682), .A4(n913), .A5(n681), 
        .Y(n825) );
  AND2X1_LVT U876 ( .A1(n683), .A2(n933), .Y(n913) );
  AO22X1_LVT U877 ( .A1(SH[1]), .A2(n980), .A3(n684), .A4(n968), .Y(n933) );
  AO22X1_LVT U878 ( .A1(SH[0]), .A2(A[2]), .A3(n679), .A4(A[3]), .Y(n968) );
  AO22X1_LVT U879 ( .A1(SH[0]), .A2(A[0]), .A3(n679), .A4(A[1]), .Y(n980) );
  AO22X1_LVT U880 ( .A1(SH[2]), .A2(n932), .A3(n683), .A4(n959), .Y(n914) );
  AO22X1_LVT U881 ( .A1(SH[1]), .A2(n967), .A3(n684), .A4(n965), .Y(n959) );
  AO22X1_LVT U882 ( .A1(SH[0]), .A2(A[10]), .A3(n679), .A4(A[11]), .Y(n965) );
  AO22X1_LVT U883 ( .A1(SH[0]), .A2(A[8]), .A3(n679), .A4(A[9]), .Y(n967) );
  AO22X1_LVT U884 ( .A1(SH[1]), .A2(n969), .A3(n684), .A4(n966), .Y(n932) );
  AO22X1_LVT U885 ( .A1(SH[0]), .A2(A[6]), .A3(n679), .A4(A[7]), .Y(n966) );
  AO22X1_LVT U886 ( .A1(SH[0]), .A2(A[4]), .A3(n679), .A4(A[5]), .Y(n969) );
  AND2X1_LVT U887 ( .A1(SH[5]), .A2(n707), .Y(B[119]) );
  AND3X1_LVT U888 ( .A1(SH[3]), .A2(SH[4]), .A3(n981), .Y(n707) );
  AND3X1_LVT U889 ( .A1(SH[4]), .A2(SH[5]), .A3(n708), .Y(B[118]) );
  AND3X1_LVT U890 ( .A1(SH[4]), .A2(SH[5]), .A3(n710), .Y(B[117]) );
  AND3X1_LVT U891 ( .A1(SH[4]), .A2(SH[5]), .A3(n712), .Y(B[116]) );
  AND3X1_LVT U892 ( .A1(SH[4]), .A2(SH[5]), .A3(n714), .Y(B[115]) );
  OA222X1_LVT U893 ( .A1(SH[3]), .A2(SH[2]), .A3(SH[3]), .A4(n982), .A5(n682), 
        .A6(n983), .Y(n714) );
  AND3X1_LVT U894 ( .A1(SH[4]), .A2(SH[5]), .A3(n716), .Y(B[114]) );
  AO22X1_LVT U895 ( .A1(SH[3]), .A2(n984), .A3(n682), .A4(n977), .Y(n716) );
  AND3X1_LVT U896 ( .A1(SH[4]), .A2(SH[5]), .A3(n718), .Y(B[113]) );
  AO22X1_LVT U897 ( .A1(SH[3]), .A2(n985), .A3(n682), .A4(n978), .Y(n718) );
  AND3X1_LVT U898 ( .A1(SH[4]), .A2(SH[5]), .A3(n720), .Y(B[112]) );
  AO22X1_LVT U899 ( .A1(SH[3]), .A2(n986), .A3(n682), .A4(n979), .Y(n720) );
  AND3X1_LVT U900 ( .A1(SH[4]), .A2(SH[5]), .A3(n723), .Y(B[111]) );
  AO22X1_LVT U901 ( .A1(SH[3]), .A2(n987), .A3(n682), .A4(n981), .Y(n723) );
  AND2X1_LVT U902 ( .A1(SH[5]), .A2(n726), .Y(B[110]) );
  AO22X1_LVT U903 ( .A1(SH[4]), .A2(n760), .A3(n681), .A4(n691), .Y(n726) );
  AND3X1_LVT U904 ( .A1(SH[3]), .A2(SH[2]), .A3(n988), .Y(n691) );
  AO22X1_LVT U905 ( .A1(SH[3]), .A2(n989), .A3(n682), .A4(n990), .Y(n760) );
  AND2X1_LVT U906 ( .A1(n830), .A2(n680), .Y(B[10]) );
  OA221X1_LVT U907 ( .A1(SH[3]), .A2(n920), .A3(n682), .A4(n919), .A5(n681), 
        .Y(n830) );
  AND2X1_LVT U908 ( .A1(n683), .A2(n938), .Y(n919) );
  OA222X1_LVT U909 ( .A1(n684), .A2(A[0]), .A3(n684), .A4(n679), .A5(SH[1]), 
        .A6(n971), .Y(n938) );
  AO22X1_LVT U910 ( .A1(SH[0]), .A2(A[1]), .A3(n679), .A4(A[2]), .Y(n971) );
  AO22X1_LVT U911 ( .A1(SH[2]), .A2(n937), .A3(n683), .A4(n962), .Y(n920) );
  AO22X1_LVT U912 ( .A1(SH[1]), .A2(n975), .A3(n684), .A4(n973), .Y(n962) );
  AO22X1_LVT U913 ( .A1(SH[0]), .A2(A[9]), .A3(n679), .A4(A[10]), .Y(n973) );
  AO22X1_LVT U914 ( .A1(SH[0]), .A2(A[7]), .A3(n679), .A4(A[8]), .Y(n975) );
  AO22X1_LVT U915 ( .A1(SH[1]), .A2(n972), .A3(n684), .A4(n974), .Y(n937) );
  AO22X1_LVT U916 ( .A1(SH[0]), .A2(A[5]), .A3(n679), .A4(A[6]), .Y(n974) );
  AO22X1_LVT U917 ( .A1(SH[0]), .A2(A[3]), .A3(n679), .A4(A[4]), .Y(n972) );
  AND2X1_LVT U918 ( .A1(SH[5]), .A2(n728), .Y(B[109]) );
  OA222X1_LVT U919 ( .A1(SH[4]), .A2(SH[3]), .A3(SH[4]), .A4(n976), .A5(n681), 
        .A6(n763), .Y(n728) );
  AO22X1_LVT U920 ( .A1(SH[3]), .A2(n991), .A3(n682), .A4(n992), .Y(n763) );
  AND2X1_LVT U921 ( .A1(SH[5]), .A2(n730), .Y(B[108]) );
  AO22X1_LVT U922 ( .A1(SH[4]), .A2(n766), .A3(n681), .A4(n695), .Y(n730) );
  AND3X1_LVT U923 ( .A1(SH[2]), .A2(SH[3]), .A3(n993), .Y(n695) );
  AO22X1_LVT U924 ( .A1(SH[3]), .A2(n994), .A3(n682), .A4(n995), .Y(n766) );
  AND2X1_LVT U925 ( .A1(SH[5]), .A2(n732), .Y(B[107]) );
  AO22X1_LVT U926 ( .A1(SH[4]), .A2(n770), .A3(n681), .A4(n697), .Y(n732) );
  AND3X1_LVT U927 ( .A1(SH[2]), .A2(SH[3]), .A3(n982), .Y(n697) );
  AO22X1_LVT U928 ( .A1(SH[3]), .A2(n795), .A3(n682), .A4(n983), .Y(n770) );
  AO22X1_LVT U929 ( .A1(SH[2]), .A2(n996), .A3(n683), .A4(n997), .Y(n983) );
  AO22X1_LVT U930 ( .A1(SH[2]), .A2(n998), .A3(n683), .A4(n999), .Y(n795) );
  AND2X1_LVT U931 ( .A1(SH[5]), .A2(n734), .Y(B[106]) );
  OA222X1_LVT U932 ( .A1(SH[4]), .A2(SH[3]), .A3(SH[4]), .A4(n977), .A5(n681), 
        .A6(n773), .Y(n734) );
  AO22X1_LVT U933 ( .A1(SH[3]), .A2(n799), .A3(n682), .A4(n984), .Y(n773) );
  AO22X1_LVT U934 ( .A1(SH[2]), .A2(n1000), .A3(n683), .A4(n1001), .Y(n984) );
  AO22X1_LVT U935 ( .A1(SH[2]), .A2(n1002), .A3(n683), .A4(n1003), .Y(n799) );
  AO22X1_LVT U936 ( .A1(SH[2]), .A2(n1004), .A3(n683), .A4(n988), .Y(n977) );
  AND2X1_LVT U937 ( .A1(SH[5]), .A2(n736), .Y(B[105]) );
  OA222X1_LVT U938 ( .A1(SH[4]), .A2(SH[3]), .A3(SH[4]), .A4(n978), .A5(n681), 
        .A6(n776), .Y(n736) );
  AO22X1_LVT U939 ( .A1(SH[3]), .A2(n804), .A3(n682), .A4(n985), .Y(n776) );
  AO22X1_LVT U940 ( .A1(SH[2]), .A2(n1005), .A3(n683), .A4(n1006), .Y(n985) );
  AO22X1_LVT U941 ( .A1(SH[2]), .A2(n1007), .A3(n683), .A4(n1008), .Y(n804) );
  OA222X1_LVT U942 ( .A1(SH[2]), .A2(SH[1]), .A3(SH[2]), .A4(n1009), .A5(n683), 
        .A6(n1010), .Y(n978) );
  AND2X1_LVT U943 ( .A1(SH[5]), .A2(n738), .Y(B[104]) );
  OA222X1_LVT U944 ( .A1(SH[4]), .A2(SH[3]), .A3(SH[4]), .A4(n979), .A5(n681), 
        .A6(n779), .Y(n738) );
  AO22X1_LVT U945 ( .A1(SH[3]), .A2(n808), .A3(n682), .A4(n986), .Y(n779) );
  AO22X1_LVT U946 ( .A1(SH[2]), .A2(n1011), .A3(n683), .A4(n1012), .Y(n986) );
  AO22X1_LVT U947 ( .A1(SH[2]), .A2(n1013), .A3(n683), .A4(n1014), .Y(n808) );
  AO22X1_LVT U948 ( .A1(SH[2]), .A2(n1015), .A3(n683), .A4(n993), .Y(n979) );
  AND2X1_LVT U949 ( .A1(SH[5]), .A2(n740), .Y(B[103]) );
  OA222X1_LVT U950 ( .A1(SH[4]), .A2(SH[3]), .A3(SH[4]), .A4(n981), .A5(n681), 
        .A6(n782), .Y(n740) );
  AO22X1_LVT U951 ( .A1(SH[3]), .A2(n812), .A3(n682), .A4(n987), .Y(n782) );
  AO22X1_LVT U952 ( .A1(SH[2]), .A2(n999), .A3(n683), .A4(n996), .Y(n987) );
  AO22X1_LVT U953 ( .A1(SH[1]), .A2(n1016), .A3(n684), .A4(n1017), .Y(n996) );
  AO22X1_LVT U954 ( .A1(SH[1]), .A2(n1018), .A3(n684), .A4(n1019), .Y(n999) );
  AO22X1_LVT U955 ( .A1(SH[2]), .A2(n829), .A3(n683), .A4(n998), .Y(n812) );
  AO22X1_LVT U956 ( .A1(SH[1]), .A2(n1020), .A3(n684), .A4(n1021), .Y(n998) );
  AO22X1_LVT U957 ( .A1(SH[1]), .A2(n1022), .A3(n684), .A4(n1023), .Y(n829) );
  AO22X1_LVT U958 ( .A1(SH[2]), .A2(n997), .A3(n683), .A4(n982), .Y(n981) );
  AO22X1_LVT U959 ( .A1(SH[1]), .A2(n1024), .A3(n684), .A4(n1009), .Y(n982) );
  AO22X1_LVT U960 ( .A1(SH[1]), .A2(n1025), .A3(n684), .A4(n1026), .Y(n997) );
  AND2X1_LVT U961 ( .A1(SH[5]), .A2(n742), .Y(B[102]) );
  AO22X1_LVT U962 ( .A1(SH[4]), .A2(n785), .A3(n681), .A4(n708), .Y(n742) );
  OA222X1_LVT U963 ( .A1(SH[3]), .A2(SH[2]), .A3(SH[3]), .A4(n988), .A5(n682), 
        .A6(n990), .Y(n708) );
  AO22X1_LVT U964 ( .A1(SH[2]), .A2(n1001), .A3(n683), .A4(n1004), .Y(n990) );
  AO22X1_LVT U965 ( .A1(SH[1]), .A2(n1027), .A3(n684), .A4(n1028), .Y(n1004)
         );
  AO22X1_LVT U966 ( .A1(SH[1]), .A2(n1029), .A3(n684), .A4(n1030), .Y(n1001)
         );
  AND3X1_LVT U967 ( .A1(SH[1]), .A2(SH[0]), .A3(A[63]), .Y(n988) );
  AO22X1_LVT U968 ( .A1(SH[3]), .A2(n816), .A3(n682), .A4(n989), .Y(n785) );
  AO22X1_LVT U969 ( .A1(SH[2]), .A2(n1003), .A3(n683), .A4(n1000), .Y(n989) );
  AO22X1_LVT U970 ( .A1(SH[1]), .A2(n1031), .A3(n684), .A4(n1032), .Y(n1000)
         );
  AO22X1_LVT U971 ( .A1(SH[1]), .A2(n1033), .A3(n684), .A4(n1034), .Y(n1003)
         );
  AO22X1_LVT U972 ( .A1(SH[2]), .A2(n834), .A3(n683), .A4(n1002), .Y(n816) );
  AO22X1_LVT U973 ( .A1(SH[1]), .A2(n1035), .A3(n684), .A4(n1036), .Y(n1002)
         );
  AO22X1_LVT U974 ( .A1(SH[1]), .A2(n1037), .A3(n684), .A4(n1038), .Y(n834) );
  AND2X1_LVT U975 ( .A1(SH[5]), .A2(n745), .Y(B[101]) );
  AO22X1_LVT U976 ( .A1(SH[4]), .A2(n788), .A3(n681), .A4(n710), .Y(n745) );
  AO22X1_LVT U977 ( .A1(SH[3]), .A2(n992), .A3(n682), .A4(n976), .Y(n710) );
  AND3X1_LVT U978 ( .A1(SH[1]), .A2(SH[2]), .A3(n1009), .Y(n976) );
  AO22X1_LVT U979 ( .A1(SH[0]), .A2(A[62]), .A3(n679), .A4(A[63]), .Y(n1009)
         );
  AO22X1_LVT U980 ( .A1(SH[2]), .A2(n1006), .A3(n683), .A4(n1010), .Y(n992) );
  AO22X1_LVT U981 ( .A1(SH[1]), .A2(n1026), .A3(n684), .A4(n1024), .Y(n1010)
         );
  AO22X1_LVT U982 ( .A1(SH[0]), .A2(A[60]), .A3(n679), .A4(A[61]), .Y(n1024)
         );
  AO22X1_LVT U983 ( .A1(SH[0]), .A2(A[58]), .A3(n679), .A4(A[59]), .Y(n1026)
         );
  AO22X1_LVT U984 ( .A1(SH[1]), .A2(n1017), .A3(n684), .A4(n1025), .Y(n1006)
         );
  AO22X1_LVT U985 ( .A1(SH[0]), .A2(A[56]), .A3(n679), .A4(A[57]), .Y(n1025)
         );
  AO22X1_LVT U986 ( .A1(SH[0]), .A2(A[54]), .A3(n679), .A4(A[55]), .Y(n1017)
         );
  AO22X1_LVT U987 ( .A1(SH[3]), .A2(n820), .A3(n682), .A4(n991), .Y(n788) );
  AO22X1_LVT U988 ( .A1(SH[2]), .A2(n1008), .A3(n683), .A4(n1005), .Y(n991) );
  AO22X1_LVT U989 ( .A1(SH[1]), .A2(n1019), .A3(n684), .A4(n1016), .Y(n1005)
         );
  AO22X1_LVT U990 ( .A1(SH[0]), .A2(A[52]), .A3(n679), .A4(A[53]), .Y(n1016)
         );
  AO22X1_LVT U991 ( .A1(SH[0]), .A2(A[50]), .A3(n679), .A4(A[51]), .Y(n1019)
         );
  AO22X1_LVT U992 ( .A1(SH[1]), .A2(n1021), .A3(n684), .A4(n1018), .Y(n1008)
         );
  AO22X1_LVT U993 ( .A1(SH[0]), .A2(A[48]), .A3(n679), .A4(A[49]), .Y(n1018)
         );
  AO22X1_LVT U994 ( .A1(SH[0]), .A2(A[46]), .A3(n679), .A4(A[47]), .Y(n1021)
         );
  AO22X1_LVT U995 ( .A1(SH[2]), .A2(n838), .A3(n683), .A4(n1007), .Y(n820) );
  AO22X1_LVT U996 ( .A1(SH[1]), .A2(n1023), .A3(n684), .A4(n1020), .Y(n1007)
         );
  AO22X1_LVT U997 ( .A1(SH[0]), .A2(A[44]), .A3(n679), .A4(A[45]), .Y(n1020)
         );
  AO22X1_LVT U998 ( .A1(SH[0]), .A2(A[42]), .A3(n679), .A4(A[43]), .Y(n1023)
         );
  AO22X1_LVT U999 ( .A1(SH[1]), .A2(n852), .A3(n684), .A4(n1022), .Y(n838) );
  AO22X1_LVT U1000 ( .A1(SH[0]), .A2(A[40]), .A3(n679), .A4(A[41]), .Y(n1022)
         );
  AO22X1_LVT U1001 ( .A1(SH[0]), .A2(A[38]), .A3(n679), .A4(A[39]), .Y(n852)
         );
  AND2X1_LVT U1002 ( .A1(SH[5]), .A2(n747), .Y(B[100]) );
  AO22X1_LVT U1003 ( .A1(SH[4]), .A2(n791), .A3(n681), .A4(n712), .Y(n747) );
  OA222X1_LVT U1004 ( .A1(SH[3]), .A2(SH[2]), .A3(SH[3]), .A4(n993), .A5(n682), 
        .A6(n995), .Y(n712) );
  AO22X1_LVT U1005 ( .A1(SH[2]), .A2(n1012), .A3(n683), .A4(n1015), .Y(n995)
         );
  AO22X1_LVT U1006 ( .A1(SH[1]), .A2(n1030), .A3(n684), .A4(n1027), .Y(n1015)
         );
  AO22X1_LVT U1007 ( .A1(SH[0]), .A2(A[59]), .A3(n679), .A4(A[60]), .Y(n1027)
         );
  AO22X1_LVT U1008 ( .A1(SH[0]), .A2(A[57]), .A3(n679), .A4(A[58]), .Y(n1030)
         );
  AO22X1_LVT U1009 ( .A1(SH[1]), .A2(n1032), .A3(n684), .A4(n1029), .Y(n1012)
         );
  AO22X1_LVT U1010 ( .A1(SH[0]), .A2(A[55]), .A3(n679), .A4(A[56]), .Y(n1029)
         );
  AO22X1_LVT U1011 ( .A1(SH[0]), .A2(A[53]), .A3(n679), .A4(A[54]), .Y(n1032)
         );
  OA222X1_LVT U1012 ( .A1(SH[1]), .A2(SH[0]), .A3(SH[1]), .A4(A[63]), .A5(n684), .A6(n1028), .Y(n993) );
  AO22X1_LVT U1013 ( .A1(SH[0]), .A2(A[61]), .A3(n679), .A4(A[62]), .Y(n1028)
         );
  AO22X1_LVT U1014 ( .A1(SH[3]), .A2(n824), .A3(n682), .A4(n994), .Y(n791) );
  AO22X1_LVT U1015 ( .A1(SH[2]), .A2(n1014), .A3(n683), .A4(n1011), .Y(n994)
         );
  AO22X1_LVT U1016 ( .A1(SH[1]), .A2(n1034), .A3(n684), .A4(n1031), .Y(n1011)
         );
  AO22X1_LVT U1017 ( .A1(SH[0]), .A2(A[51]), .A3(n679), .A4(A[52]), .Y(n1031)
         );
  AO22X1_LVT U1018 ( .A1(SH[0]), .A2(A[49]), .A3(n679), .A4(A[50]), .Y(n1034)
         );
  AO22X1_LVT U1019 ( .A1(SH[1]), .A2(n1036), .A3(n684), .A4(n1033), .Y(n1014)
         );
  AO22X1_LVT U1020 ( .A1(SH[0]), .A2(A[47]), .A3(n679), .A4(A[48]), .Y(n1033)
         );
  AO22X1_LVT U1021 ( .A1(SH[0]), .A2(A[45]), .A3(n679), .A4(A[46]), .Y(n1036)
         );
  AO22X1_LVT U1022 ( .A1(SH[2]), .A2(n844), .A3(n683), .A4(n1013), .Y(n824) );
  AO22X1_LVT U1023 ( .A1(SH[1]), .A2(n1038), .A3(n684), .A4(n1035), .Y(n1013)
         );
  AO22X1_LVT U1024 ( .A1(SH[0]), .A2(A[43]), .A3(n679), .A4(A[44]), .Y(n1035)
         );
  AO22X1_LVT U1025 ( .A1(SH[0]), .A2(A[41]), .A3(n679), .A4(A[42]), .Y(n1038)
         );
  AO22X1_LVT U1026 ( .A1(SH[1]), .A2(n858), .A3(n684), .A4(n1037), .Y(n844) );
  AO22X1_LVT U1027 ( .A1(SH[0]), .A2(A[39]), .A3(n679), .A4(A[40]), .Y(n1037)
         );
  AO22X1_LVT U1028 ( .A1(SH[0]), .A2(A[37]), .A3(n679), .A4(A[38]), .Y(n858)
         );
  AND3X1_LVT U1029 ( .A1(n846), .A2(n681), .A3(n682), .Y(n885) );
  AND4X1_LVT U1030 ( .A1(A[0]), .A2(n683), .A3(n684), .A4(n679), .Y(n846) );
endmodule


module MulDiv_DW01_sub_J39_0 ( A, B, CI, DIFF, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] DIFF;
  input CI;
  output CO;
  wire   n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85;

  INVX0_LVT U49 ( .A(A[2]), .Y(n69) );
  INVX0_LVT U50 ( .A(A[1]), .Y(n67) );
  INVX0_LVT U51 ( .A(A[0]), .Y(n66) );
  INVX0_LVT U52 ( .A(A[3]), .Y(n68) );
  OR2X1_LVT U53 ( .A1(n68), .A2(B[3]), .Y(n77) );
  FADDX1_LVT U54 ( .A(B[5]), .B(A[5]), .CI(n71), .S(DIFF[5]) );
  INVX1_LVT U55 ( .A(B[0]), .Y(n64) );
  INVX1_LVT U56 ( .A(B[1]), .Y(n65) );
  INVX1_LVT U57 ( .A(A[4]), .Y(n70) );
  NAND3X0_LVT U58 ( .A1(n72), .A2(n73), .A3(n74), .Y(n71) );
  NAND3X0_LVT U59 ( .A1(B[3]), .A2(n68), .A3(n75), .Y(n74) );
  NAND2X0_LVT U60 ( .A1(n75), .A2(n76), .Y(n73) );
  NAND3X0_LVT U61 ( .A1(B[4]), .A2(n70), .A3(n75), .Y(n72) );
  AO222X1_LVT U62 ( .A1(B[4]), .A2(n77), .A3(B[4]), .A4(n70), .A5(n77), .A6(
        n70), .Y(n75) );
  FADDX1_LVT U63 ( .A(A[4]), .B(B[4]), .CI(n78), .S(DIFF[4]) );
  AO22X1_LVT U64 ( .A1(B[3]), .A2(n68), .A3(n77), .A4(n76), .Y(n78) );
  FADDX1_LVT U65 ( .A(A[3]), .B(B[3]), .CI(n76), .S(DIFF[3]) );
  AND2X1_LVT U66 ( .A1(n79), .A2(n80), .Y(n76) );
  NAND3X0_LVT U67 ( .A1(n81), .A2(n82), .A3(n83), .Y(n80) );
  NAND2X0_LVT U68 ( .A1(B[2]), .A2(n69), .Y(n82) );
  AO222X1_LVT U69 ( .A1(B[2]), .A2(n69), .A3(B[2]), .A4(n84), .A5(n69), .A6(
        n84), .Y(n79) );
  NAND2X0_LVT U70 ( .A1(A[1]), .A2(n65), .Y(n84) );
  FADDX1_LVT U71 ( .A(B[2]), .B(n69), .CI(n85), .S(DIFF[2]) );
  AO22X1_LVT U72 ( .A1(A[1]), .A2(n65), .A3(n83), .A4(n81), .Y(n85) );
  NAND2X0_LVT U73 ( .A1(B[1]), .A2(n67), .Y(n81) );
  FADDX1_LVT U74 ( .A(B[1]), .B(n67), .CI(n83), .S(DIFF[1]) );
  NAND2X0_LVT U75 ( .A1(B[0]), .A2(n66), .Y(n83) );
  AO22X1_LVT U76 ( .A1(A[0]), .A2(n64), .A3(n66), .A4(B[0]), .Y(DIFF[0]) );
endmodule


module MulDiv_DW_rightsh_J39_0 ( A, DATA_TC, SH, B );
  input [126:0] A;
  input [5:0] SH;
  output [126:0] B;
  input DATA_TC;
  wire   n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043;

  AO22X1_LVT U696 ( .A1(n852), .A2(A[104]), .A3(n853), .A4(A[112]), .Y(n832)
         );
  AO22X1_LVT U697 ( .A1(SH[4]), .A2(n832), .A3(n854), .A4(n905), .Y(n833) );
  AO22X1_LVT U698 ( .A1(SH[5]), .A2(n833), .A3(n904), .A4(n855), .Y(B[56]) );
  AO22X1_LVT U699 ( .A1(n852), .A2(A[96]), .A3(n853), .A4(A[104]), .Y(n834) );
  AO22X1_LVT U700 ( .A1(SH[4]), .A2(n834), .A3(n854), .A4(n935), .Y(n835) );
  AO22X1_LVT U701 ( .A1(SH[5]), .A2(n835), .A3(n934), .A4(n855), .Y(B[48]) );
  AO22X1_LVT U702 ( .A1(A[12]), .A2(n852), .A3(A[20]), .A4(n853), .Y(n836) );
  AO22X1_LVT U703 ( .A1(SH[4]), .A2(n1010), .A3(n854), .A4(n836), .Y(n837) );
  AO22X1_LVT U704 ( .A1(SH[5]), .A2(n946), .A3(n855), .A4(n837), .Y(B[12]) );
  AO22X1_LVT U705 ( .A1(SH[4]), .A2(n905), .A3(n854), .A4(n960), .Y(n838) );
  AO22X1_LVT U706 ( .A1(SH[5]), .A2(n838), .A3(n860), .A4(n855), .Y(B[40]) );
  AO22X1_LVT U707 ( .A1(SH[4]), .A2(n959), .A3(n854), .A4(n862), .Y(n839) );
  AO22X1_LVT U708 ( .A1(SH[5]), .A2(n904), .A3(n855), .A4(n839), .Y(B[24]) );
  AO22X1_LVT U709 ( .A1(n852), .A2(A[2]), .A3(n853), .A4(A[10]), .Y(n840) );
  AO22X1_LVT U710 ( .A1(SH[4]), .A2(n1001), .A3(n854), .A4(n840), .Y(n841) );
  AO22X1_LVT U711 ( .A1(SH[5]), .A2(n986), .A3(n855), .A4(n841), .Y(B[2]) );
  AO22X1_LVT U712 ( .A1(SH[4]), .A2(n1031), .A3(n854), .A4(n1032), .Y(n842) );
  AO22X1_LVT U713 ( .A1(SH[5]), .A2(n934), .A3(n855), .A4(n842), .Y(B[16]) );
  AO22X1_LVT U714 ( .A1(n852), .A2(A[4]), .A3(A[12]), .A4(n853), .Y(n843) );
  AO22X1_LVT U715 ( .A1(SH[4]), .A2(n929), .A3(n854), .A4(n843), .Y(n844) );
  AO22X1_LVT U716 ( .A1(SH[5]), .A2(n928), .A3(n855), .A4(n844), .Y(B[4]) );
  AO22X1_LVT U717 ( .A1(n852), .A2(A[0]), .A3(n853), .A4(A[8]), .Y(n845) );
  AO22X1_LVT U718 ( .A1(SH[4]), .A2(n1032), .A3(n854), .A4(n845), .Y(n846) );
  AO22X1_LVT U719 ( .A1(SH[5]), .A2(n991), .A3(n855), .A4(n846), .Y(B[0]) );
  AO22X1_LVT U720 ( .A1(SH[3]), .A2(A[9]), .A3(n852), .A4(A[1]), .Y(n847) );
  AO22X1_LVT U721 ( .A1(SH[4]), .A2(n1025), .A3(n854), .A4(n847), .Y(n848) );
  AO22X1_LVT U722 ( .A1(SH[5]), .A2(n989), .A3(n855), .A4(n848), .Y(B[1]) );
  AO22X1_LVT U723 ( .A1(SH[4]), .A2(n935), .A3(n854), .A4(n992), .Y(n849) );
  AO22X1_LVT U724 ( .A1(SH[5]), .A2(n849), .A3(n991), .A4(n855), .Y(B[32]) );
  AO22X1_LVT U725 ( .A1(n852), .A2(A[100]), .A3(n853), .A4(A[108]), .Y(n850)
         );
  AO22X1_LVT U726 ( .A1(SH[4]), .A2(n850), .A3(n854), .A4(n919), .Y(n851) );
  AO22X1_LVT U727 ( .A1(SH[5]), .A2(n851), .A3(n918), .A4(n855), .Y(B[52]) );
  INVX1_LVT U728 ( .A(SH[3]), .Y(n852) );
  INVX1_LVT U729 ( .A(n852), .Y(n853) );
  INVX1_LVT U730 ( .A(SH[5]), .Y(n855) );
  INVX1_LVT U731 ( .A(SH[4]), .Y(n854) );
  AO22X1_LVT U732 ( .A1(SH[5]), .A2(n856), .A3(n855), .A4(n857), .Y(B[9]) );
  AO22X1_LVT U733 ( .A1(SH[4]), .A2(n858), .A3(n854), .A4(n859), .Y(n857) );
  AO22X1_LVT U734 ( .A1(n853), .A2(A[17]), .A3(n852), .A4(A[9]), .Y(n859) );
  AO22X1_LVT U735 ( .A1(SH[5]), .A2(n860), .A3(n855), .A4(n861), .Y(B[8]) );
  AO22X1_LVT U736 ( .A1(SH[4]), .A2(n862), .A3(n854), .A4(n863), .Y(n861) );
  AO22X1_LVT U737 ( .A1(SH[3]), .A2(A[16]), .A3(n852), .A4(A[8]), .Y(n863) );
  AO22X1_LVT U738 ( .A1(SH[5]), .A2(n864), .A3(n855), .A4(n865), .Y(B[7]) );
  AO22X1_LVT U739 ( .A1(SH[4]), .A2(n866), .A3(n854), .A4(n867), .Y(n865) );
  AO22X1_LVT U740 ( .A1(n853), .A2(A[15]), .A3(n852), .A4(A[7]), .Y(n867) );
  AO22X1_LVT U741 ( .A1(SH[5]), .A2(n868), .A3(n855), .A4(n869), .Y(B[6]) );
  AO22X1_LVT U742 ( .A1(SH[4]), .A2(n870), .A3(n854), .A4(n871), .Y(n869) );
  AO22X1_LVT U743 ( .A1(SH[3]), .A2(A[14]), .A3(n852), .A4(A[6]), .Y(n871) );
  AO22X1_LVT U744 ( .A1(SH[5]), .A2(n872), .A3(n855), .A4(n873), .Y(B[63]) );
  AO22X1_LVT U745 ( .A1(SH[4]), .A2(n874), .A3(n854), .A4(n875), .Y(n872) );
  AO22X1_LVT U746 ( .A1(n853), .A2(A[119]), .A3(n852), .A4(A[111]), .Y(n874)
         );
  AO22X1_LVT U747 ( .A1(SH[5]), .A2(n876), .A3(n855), .A4(n877), .Y(B[62]) );
  AO22X1_LVT U748 ( .A1(SH[4]), .A2(n878), .A3(n854), .A4(n879), .Y(n876) );
  AO22X1_LVT U749 ( .A1(n853), .A2(A[118]), .A3(n852), .A4(A[110]), .Y(n878)
         );
  AO22X1_LVT U750 ( .A1(SH[5]), .A2(n880), .A3(n855), .A4(n881), .Y(B[61]) );
  AO22X1_LVT U751 ( .A1(SH[4]), .A2(n882), .A3(n854), .A4(n883), .Y(n880) );
  AO22X1_LVT U752 ( .A1(n853), .A2(A[117]), .A3(n852), .A4(A[109]), .Y(n882)
         );
  AO22X1_LVT U753 ( .A1(SH[5]), .A2(n884), .A3(n855), .A4(n885), .Y(B[60]) );
  AO22X1_LVT U754 ( .A1(SH[4]), .A2(n886), .A3(n854), .A4(n887), .Y(n884) );
  AO22X1_LVT U755 ( .A1(SH[3]), .A2(A[116]), .A3(n852), .A4(A[108]), .Y(n886)
         );
  AO22X1_LVT U756 ( .A1(SH[5]), .A2(n888), .A3(n855), .A4(n889), .Y(B[5]) );
  AO22X1_LVT U757 ( .A1(SH[4]), .A2(n890), .A3(n854), .A4(n891), .Y(n889) );
  AO22X1_LVT U758 ( .A1(n853), .A2(A[13]), .A3(n852), .A4(A[5]), .Y(n891) );
  AO22X1_LVT U759 ( .A1(SH[5]), .A2(n892), .A3(n855), .A4(n893), .Y(B[59]) );
  AO22X1_LVT U760 ( .A1(SH[4]), .A2(n894), .A3(n854), .A4(n895), .Y(n892) );
  AO22X1_LVT U761 ( .A1(n853), .A2(A[115]), .A3(n852), .A4(A[107]), .Y(n894)
         );
  AO22X1_LVT U762 ( .A1(SH[5]), .A2(n896), .A3(n855), .A4(n897), .Y(B[58]) );
  AO22X1_LVT U763 ( .A1(SH[4]), .A2(n898), .A3(n854), .A4(n899), .Y(n896) );
  AO22X1_LVT U764 ( .A1(n853), .A2(A[114]), .A3(n852), .A4(A[106]), .Y(n898)
         );
  AO22X1_LVT U765 ( .A1(SH[5]), .A2(n900), .A3(n855), .A4(n901), .Y(B[57]) );
  AO22X1_LVT U766 ( .A1(SH[4]), .A2(n902), .A3(n854), .A4(n903), .Y(n900) );
  AO22X1_LVT U767 ( .A1(SH[3]), .A2(A[113]), .A3(n852), .A4(A[105]), .Y(n902)
         );
  AO22X1_LVT U768 ( .A1(SH[5]), .A2(n906), .A3(n855), .A4(n907), .Y(B[55]) );
  AO22X1_LVT U769 ( .A1(SH[4]), .A2(n908), .A3(n854), .A4(n909), .Y(n906) );
  AO22X1_LVT U770 ( .A1(n853), .A2(A[111]), .A3(n852), .A4(A[103]), .Y(n908)
         );
  AO22X1_LVT U771 ( .A1(SH[5]), .A2(n910), .A3(n855), .A4(n911), .Y(B[54]) );
  AO22X1_LVT U772 ( .A1(SH[4]), .A2(n912), .A3(n854), .A4(n913), .Y(n910) );
  AO22X1_LVT U773 ( .A1(n853), .A2(A[110]), .A3(n852), .A4(A[102]), .Y(n912)
         );
  AO22X1_LVT U774 ( .A1(SH[5]), .A2(n914), .A3(n855), .A4(n915), .Y(B[53]) );
  AO22X1_LVT U775 ( .A1(SH[4]), .A2(n916), .A3(n854), .A4(n917), .Y(n914) );
  AO22X1_LVT U776 ( .A1(SH[3]), .A2(A[109]), .A3(n852), .A4(A[101]), .Y(n916)
         );
  AO22X1_LVT U777 ( .A1(SH[5]), .A2(n920), .A3(n855), .A4(n921), .Y(B[51]) );
  AO22X1_LVT U778 ( .A1(SH[4]), .A2(n922), .A3(n854), .A4(n923), .Y(n920) );
  AO22X1_LVT U779 ( .A1(n853), .A2(A[107]), .A3(n852), .A4(A[99]), .Y(n922) );
  AO22X1_LVT U780 ( .A1(SH[5]), .A2(n924), .A3(n855), .A4(n925), .Y(B[50]) );
  AO22X1_LVT U781 ( .A1(SH[4]), .A2(n926), .A3(n854), .A4(n927), .Y(n924) );
  AO22X1_LVT U782 ( .A1(n853), .A2(A[106]), .A3(n852), .A4(A[98]), .Y(n926) );
  AO22X1_LVT U783 ( .A1(SH[5]), .A2(n930), .A3(n855), .A4(n931), .Y(B[49]) );
  AO22X1_LVT U784 ( .A1(SH[4]), .A2(n932), .A3(n854), .A4(n933), .Y(n930) );
  AO22X1_LVT U785 ( .A1(SH[3]), .A2(A[105]), .A3(n852), .A4(A[97]), .Y(n932)
         );
  AO22X1_LVT U786 ( .A1(SH[5]), .A2(n936), .A3(n855), .A4(n937), .Y(B[47]) );
  AO22X1_LVT U787 ( .A1(SH[4]), .A2(n875), .A3(n854), .A4(n938), .Y(n936) );
  AO22X1_LVT U788 ( .A1(n853), .A2(A[103]), .A3(n852), .A4(A[95]), .Y(n875) );
  AO22X1_LVT U789 ( .A1(SH[5]), .A2(n939), .A3(n855), .A4(n940), .Y(B[46]) );
  AO22X1_LVT U790 ( .A1(SH[4]), .A2(n879), .A3(n854), .A4(n941), .Y(n939) );
  AO22X1_LVT U791 ( .A1(n853), .A2(A[102]), .A3(n852), .A4(A[94]), .Y(n879) );
  AO22X1_LVT U792 ( .A1(SH[5]), .A2(n942), .A3(n855), .A4(n943), .Y(B[45]) );
  AO22X1_LVT U793 ( .A1(SH[4]), .A2(n883), .A3(n854), .A4(n944), .Y(n942) );
  AO22X1_LVT U794 ( .A1(SH[3]), .A2(A[101]), .A3(n852), .A4(A[93]), .Y(n883)
         );
  AO22X1_LVT U795 ( .A1(SH[5]), .A2(n945), .A3(n855), .A4(n946), .Y(B[44]) );
  AO22X1_LVT U796 ( .A1(SH[4]), .A2(n887), .A3(n854), .A4(n947), .Y(n945) );
  AO22X1_LVT U797 ( .A1(n853), .A2(A[100]), .A3(n852), .A4(A[92]), .Y(n887) );
  AO22X1_LVT U798 ( .A1(SH[5]), .A2(n948), .A3(n855), .A4(n949), .Y(B[43]) );
  AO22X1_LVT U799 ( .A1(SH[4]), .A2(n895), .A3(n854), .A4(n950), .Y(n948) );
  AO22X1_LVT U800 ( .A1(n853), .A2(A[99]), .A3(n852), .A4(A[91]), .Y(n895) );
  AO22X1_LVT U801 ( .A1(SH[5]), .A2(n951), .A3(n855), .A4(n952), .Y(B[42]) );
  AO22X1_LVT U802 ( .A1(SH[4]), .A2(n899), .A3(n854), .A4(n953), .Y(n951) );
  AO22X1_LVT U803 ( .A1(n853), .A2(A[98]), .A3(n852), .A4(A[90]), .Y(n899) );
  AO22X1_LVT U804 ( .A1(SH[5]), .A2(n954), .A3(n855), .A4(n856), .Y(B[41]) );
  AO22X1_LVT U805 ( .A1(SH[4]), .A2(n955), .A3(n854), .A4(n956), .Y(n856) );
  AO22X1_LVT U806 ( .A1(SH[4]), .A2(n903), .A3(n854), .A4(n957), .Y(n954) );
  AO22X1_LVT U807 ( .A1(SH[3]), .A2(A[97]), .A3(n852), .A4(A[89]), .Y(n903) );
  AO22X1_LVT U808 ( .A1(SH[4]), .A2(n958), .A3(n854), .A4(n959), .Y(n860) );
  AO22X1_LVT U809 ( .A1(n853), .A2(A[96]), .A3(n852), .A4(A[88]), .Y(n905) );
  AO22X1_LVT U810 ( .A1(SH[5]), .A2(n961), .A3(n855), .A4(n962), .Y(B[3]) );
  AO22X1_LVT U811 ( .A1(SH[4]), .A2(n963), .A3(n854), .A4(n964), .Y(n962) );
  AO22X1_LVT U812 ( .A1(n853), .A2(A[11]), .A3(n852), .A4(A[3]), .Y(n964) );
  AO22X1_LVT U813 ( .A1(SH[5]), .A2(n965), .A3(n855), .A4(n864), .Y(B[39]) );
  AO22X1_LVT U814 ( .A1(SH[4]), .A2(n966), .A3(n854), .A4(n967), .Y(n864) );
  AO22X1_LVT U815 ( .A1(SH[4]), .A2(n909), .A3(n854), .A4(n968), .Y(n965) );
  AO22X1_LVT U816 ( .A1(n853), .A2(A[95]), .A3(n852), .A4(A[87]), .Y(n909) );
  AO22X1_LVT U817 ( .A1(SH[5]), .A2(n969), .A3(n855), .A4(n868), .Y(B[38]) );
  AO22X1_LVT U818 ( .A1(SH[4]), .A2(n970), .A3(n854), .A4(n971), .Y(n868) );
  AO22X1_LVT U819 ( .A1(SH[4]), .A2(n913), .A3(n854), .A4(n972), .Y(n969) );
  AO22X1_LVT U820 ( .A1(n853), .A2(A[94]), .A3(n852), .A4(A[86]), .Y(n913) );
  AO22X1_LVT U821 ( .A1(SH[5]), .A2(n973), .A3(n855), .A4(n888), .Y(B[37]) );
  AO22X1_LVT U822 ( .A1(SH[4]), .A2(n974), .A3(n854), .A4(n975), .Y(n888) );
  AO22X1_LVT U823 ( .A1(SH[4]), .A2(n917), .A3(n854), .A4(n976), .Y(n973) );
  AO22X1_LVT U824 ( .A1(n853), .A2(A[93]), .A3(n852), .A4(A[85]), .Y(n917) );
  AO22X1_LVT U825 ( .A1(SH[5]), .A2(n977), .A3(n855), .A4(n928), .Y(B[36]) );
  AO22X1_LVT U826 ( .A1(SH[4]), .A2(n978), .A3(n854), .A4(n979), .Y(n928) );
  AO22X1_LVT U827 ( .A1(SH[4]), .A2(n919), .A3(n854), .A4(n980), .Y(n977) );
  AO22X1_LVT U828 ( .A1(n853), .A2(A[92]), .A3(n852), .A4(A[84]), .Y(n919) );
  AO22X1_LVT U829 ( .A1(SH[5]), .A2(n981), .A3(n855), .A4(n961), .Y(B[35]) );
  AO22X1_LVT U830 ( .A1(SH[4]), .A2(n982), .A3(n854), .A4(n983), .Y(n961) );
  AO22X1_LVT U831 ( .A1(SH[4]), .A2(n923), .A3(n854), .A4(n984), .Y(n981) );
  AO22X1_LVT U832 ( .A1(n853), .A2(A[91]), .A3(n852), .A4(A[83]), .Y(n923) );
  AO22X1_LVT U833 ( .A1(SH[5]), .A2(n985), .A3(n855), .A4(n986), .Y(B[34]) );
  AO22X1_LVT U834 ( .A1(SH[4]), .A2(n927), .A3(n854), .A4(n987), .Y(n985) );
  AO22X1_LVT U835 ( .A1(n853), .A2(A[90]), .A3(n852), .A4(A[82]), .Y(n927) );
  AO22X1_LVT U836 ( .A1(SH[5]), .A2(n988), .A3(n855), .A4(n989), .Y(B[33]) );
  AO22X1_LVT U837 ( .A1(SH[4]), .A2(n933), .A3(n854), .A4(n990), .Y(n988) );
  AO22X1_LVT U838 ( .A1(n853), .A2(A[89]), .A3(n852), .A4(A[81]), .Y(n933) );
  AO22X1_LVT U839 ( .A1(n853), .A2(A[88]), .A3(n852), .A4(A[80]), .Y(n935) );
  AO22X1_LVT U840 ( .A1(SH[5]), .A2(n873), .A3(n855), .A4(n993), .Y(B[31]) );
  AO22X1_LVT U841 ( .A1(SH[4]), .A2(n994), .A3(n854), .A4(n995), .Y(n993) );
  AO22X1_LVT U842 ( .A1(SH[4]), .A2(n938), .A3(n854), .A4(n996), .Y(n873) );
  AO22X1_LVT U843 ( .A1(n853), .A2(A[87]), .A3(n852), .A4(A[79]), .Y(n938) );
  AO22X1_LVT U844 ( .A1(SH[5]), .A2(n877), .A3(n855), .A4(n997), .Y(B[30]) );
  AO22X1_LVT U845 ( .A1(SH[4]), .A2(n998), .A3(n854), .A4(n999), .Y(n997) );
  AO22X1_LVT U846 ( .A1(SH[4]), .A2(n941), .A3(n854), .A4(n1000), .Y(n877) );
  AO22X1_LVT U847 ( .A1(n853), .A2(A[86]), .A3(n852), .A4(A[78]), .Y(n941) );
  AO22X1_LVT U848 ( .A1(SH[4]), .A2(n1002), .A3(n854), .A4(n1003), .Y(n986) );
  AO22X1_LVT U849 ( .A1(SH[5]), .A2(n881), .A3(n855), .A4(n1004), .Y(B[29]) );
  AO22X1_LVT U850 ( .A1(SH[4]), .A2(n1005), .A3(n854), .A4(n1006), .Y(n1004)
         );
  AO22X1_LVT U851 ( .A1(SH[4]), .A2(n944), .A3(n854), .A4(n1007), .Y(n881) );
  AO22X1_LVT U852 ( .A1(n853), .A2(A[85]), .A3(n852), .A4(A[77]), .Y(n944) );
  AO22X1_LVT U853 ( .A1(SH[5]), .A2(n885), .A3(n855), .A4(n1008), .Y(B[28]) );
  AO22X1_LVT U854 ( .A1(SH[4]), .A2(n1009), .A3(n854), .A4(n1010), .Y(n1008)
         );
  AO22X1_LVT U855 ( .A1(SH[4]), .A2(n947), .A3(n854), .A4(n1011), .Y(n885) );
  AO22X1_LVT U856 ( .A1(n853), .A2(A[84]), .A3(n852), .A4(A[76]), .Y(n947) );
  AO22X1_LVT U857 ( .A1(SH[5]), .A2(n893), .A3(n855), .A4(n1012), .Y(B[27]) );
  AO22X1_LVT U858 ( .A1(SH[4]), .A2(n1013), .A3(n854), .A4(n1014), .Y(n1012)
         );
  AO22X1_LVT U859 ( .A1(SH[4]), .A2(n950), .A3(n854), .A4(n1015), .Y(n893) );
  AO22X1_LVT U860 ( .A1(n853), .A2(A[83]), .A3(n852), .A4(A[75]), .Y(n950) );
  AO22X1_LVT U861 ( .A1(SH[5]), .A2(n897), .A3(n855), .A4(n1016), .Y(B[26]) );
  AO22X1_LVT U862 ( .A1(SH[4]), .A2(n1017), .A3(n854), .A4(n1018), .Y(n1016)
         );
  AO22X1_LVT U863 ( .A1(SH[4]), .A2(n953), .A3(n854), .A4(n1019), .Y(n897) );
  AO22X1_LVT U864 ( .A1(n853), .A2(A[82]), .A3(n852), .A4(A[74]), .Y(n953) );
  AO22X1_LVT U865 ( .A1(SH[5]), .A2(n901), .A3(n855), .A4(n1020), .Y(B[25]) );
  AO22X1_LVT U866 ( .A1(SH[4]), .A2(n956), .A3(n854), .A4(n858), .Y(n1020) );
  AO22X1_LVT U867 ( .A1(n853), .A2(A[33]), .A3(n852), .A4(A[25]), .Y(n858) );
  AO22X1_LVT U868 ( .A1(n853), .A2(A[49]), .A3(n852), .A4(A[41]), .Y(n956) );
  AO22X1_LVT U869 ( .A1(SH[4]), .A2(n957), .A3(n854), .A4(n955), .Y(n901) );
  AO22X1_LVT U870 ( .A1(n853), .A2(A[65]), .A3(n852), .A4(A[57]), .Y(n955) );
  AO22X1_LVT U871 ( .A1(n853), .A2(A[81]), .A3(n852), .A4(A[73]), .Y(n957) );
  AO22X1_LVT U872 ( .A1(n853), .A2(A[32]), .A3(n852), .A4(A[24]), .Y(n862) );
  AO22X1_LVT U873 ( .A1(n853), .A2(A[48]), .A3(n852), .A4(A[40]), .Y(n959) );
  AO22X1_LVT U874 ( .A1(SH[4]), .A2(n960), .A3(n854), .A4(n958), .Y(n904) );
  AO22X1_LVT U875 ( .A1(n853), .A2(A[64]), .A3(n852), .A4(A[56]), .Y(n958) );
  AO22X1_LVT U876 ( .A1(n853), .A2(A[80]), .A3(n852), .A4(A[72]), .Y(n960) );
  AO22X1_LVT U877 ( .A1(SH[5]), .A2(n907), .A3(n855), .A4(n1021), .Y(B[23]) );
  AO22X1_LVT U878 ( .A1(SH[4]), .A2(n967), .A3(n854), .A4(n866), .Y(n1021) );
  AO22X1_LVT U879 ( .A1(n853), .A2(A[31]), .A3(n852), .A4(A[23]), .Y(n866) );
  AO22X1_LVT U880 ( .A1(n853), .A2(A[47]), .A3(n852), .A4(A[39]), .Y(n967) );
  AO22X1_LVT U881 ( .A1(SH[4]), .A2(n968), .A3(n854), .A4(n966), .Y(n907) );
  AO22X1_LVT U882 ( .A1(n853), .A2(A[63]), .A3(n852), .A4(A[55]), .Y(n966) );
  AO22X1_LVT U883 ( .A1(n853), .A2(A[79]), .A3(n852), .A4(A[71]), .Y(n968) );
  AO22X1_LVT U884 ( .A1(SH[5]), .A2(n911), .A3(n855), .A4(n1022), .Y(B[22]) );
  AO22X1_LVT U885 ( .A1(SH[4]), .A2(n971), .A3(n854), .A4(n870), .Y(n1022) );
  AO22X1_LVT U886 ( .A1(n853), .A2(A[30]), .A3(n852), .A4(A[22]), .Y(n870) );
  AO22X1_LVT U887 ( .A1(n853), .A2(A[46]), .A3(n852), .A4(A[38]), .Y(n971) );
  AO22X1_LVT U888 ( .A1(SH[4]), .A2(n972), .A3(n854), .A4(n970), .Y(n911) );
  AO22X1_LVT U889 ( .A1(n853), .A2(A[62]), .A3(n852), .A4(A[54]), .Y(n970) );
  AO22X1_LVT U890 ( .A1(n853), .A2(A[78]), .A3(n852), .A4(A[70]), .Y(n972) );
  AO22X1_LVT U891 ( .A1(SH[5]), .A2(n915), .A3(n855), .A4(n1023), .Y(B[21]) );
  AO22X1_LVT U892 ( .A1(SH[4]), .A2(n975), .A3(n854), .A4(n890), .Y(n1023) );
  AO22X1_LVT U893 ( .A1(n853), .A2(A[29]), .A3(n852), .A4(A[21]), .Y(n890) );
  AO22X1_LVT U894 ( .A1(n853), .A2(A[45]), .A3(n852), .A4(A[37]), .Y(n975) );
  AO22X1_LVT U895 ( .A1(SH[4]), .A2(n976), .A3(n854), .A4(n974), .Y(n915) );
  AO22X1_LVT U896 ( .A1(n853), .A2(A[61]), .A3(n852), .A4(A[53]), .Y(n974) );
  AO22X1_LVT U897 ( .A1(n853), .A2(A[77]), .A3(n852), .A4(A[69]), .Y(n976) );
  AO22X1_LVT U898 ( .A1(SH[5]), .A2(n918), .A3(n855), .A4(n1024), .Y(B[20]) );
  AO22X1_LVT U899 ( .A1(SH[4]), .A2(n979), .A3(n854), .A4(n929), .Y(n1024) );
  AO22X1_LVT U900 ( .A1(SH[3]), .A2(A[28]), .A3(n852), .A4(A[20]), .Y(n929) );
  AO22X1_LVT U901 ( .A1(n853), .A2(A[44]), .A3(n852), .A4(A[36]), .Y(n979) );
  AO22X1_LVT U902 ( .A1(SH[4]), .A2(n980), .A3(n854), .A4(n978), .Y(n918) );
  AO22X1_LVT U903 ( .A1(n853), .A2(A[60]), .A3(n852), .A4(A[52]), .Y(n978) );
  AO22X1_LVT U904 ( .A1(n853), .A2(A[76]), .A3(n852), .A4(A[68]), .Y(n980) );
  AO22X1_LVT U905 ( .A1(SH[4]), .A2(n1026), .A3(n854), .A4(n1027), .Y(n989) );
  AO22X1_LVT U906 ( .A1(SH[5]), .A2(n921), .A3(n855), .A4(n1028), .Y(B[19]) );
  AO22X1_LVT U907 ( .A1(SH[4]), .A2(n983), .A3(n854), .A4(n963), .Y(n1028) );
  AO22X1_LVT U908 ( .A1(n853), .A2(A[27]), .A3(n852), .A4(A[19]), .Y(n963) );
  AO22X1_LVT U909 ( .A1(n853), .A2(A[43]), .A3(n852), .A4(A[35]), .Y(n983) );
  AO22X1_LVT U910 ( .A1(SH[4]), .A2(n984), .A3(n854), .A4(n982), .Y(n921) );
  AO22X1_LVT U911 ( .A1(n853), .A2(A[59]), .A3(n852), .A4(A[51]), .Y(n982) );
  AO22X1_LVT U912 ( .A1(SH[3]), .A2(A[75]), .A3(n852), .A4(A[67]), .Y(n984) );
  AO22X1_LVT U913 ( .A1(SH[5]), .A2(n925), .A3(n855), .A4(n1029), .Y(B[18]) );
  AO22X1_LVT U914 ( .A1(SH[4]), .A2(n1003), .A3(n854), .A4(n1001), .Y(n1029)
         );
  AO22X1_LVT U915 ( .A1(n853), .A2(A[26]), .A3(n852), .A4(A[18]), .Y(n1001) );
  AO22X1_LVT U916 ( .A1(n853), .A2(A[42]), .A3(n852), .A4(A[34]), .Y(n1003) );
  AO22X1_LVT U917 ( .A1(SH[4]), .A2(n987), .A3(n854), .A4(n1002), .Y(n925) );
  AO22X1_LVT U918 ( .A1(n853), .A2(A[58]), .A3(n852), .A4(A[50]), .Y(n1002) );
  AO22X1_LVT U919 ( .A1(n853), .A2(A[74]), .A3(n852), .A4(A[66]), .Y(n987) );
  AO22X1_LVT U920 ( .A1(SH[5]), .A2(n931), .A3(n855), .A4(n1030), .Y(B[17]) );
  AO22X1_LVT U921 ( .A1(SH[4]), .A2(n1027), .A3(n854), .A4(n1025), .Y(n1030)
         );
  AO22X1_LVT U922 ( .A1(n853), .A2(A[25]), .A3(n852), .A4(A[17]), .Y(n1025) );
  AO22X1_LVT U923 ( .A1(n853), .A2(A[41]), .A3(n852), .A4(A[33]), .Y(n1027) );
  AO22X1_LVT U924 ( .A1(SH[4]), .A2(n990), .A3(n854), .A4(n1026), .Y(n931) );
  AO22X1_LVT U925 ( .A1(n853), .A2(A[57]), .A3(n852), .A4(A[49]), .Y(n1026) );
  AO22X1_LVT U926 ( .A1(n853), .A2(A[73]), .A3(n852), .A4(A[65]), .Y(n990) );
  AO22X1_LVT U927 ( .A1(SH[4]), .A2(n992), .A3(n854), .A4(n1033), .Y(n934) );
  AO22X1_LVT U928 ( .A1(n853), .A2(A[72]), .A3(n852), .A4(A[64]), .Y(n992) );
  AO22X1_LVT U929 ( .A1(SH[5]), .A2(n937), .A3(n855), .A4(n1034), .Y(B[15]) );
  AO22X1_LVT U930 ( .A1(SH[4]), .A2(n995), .A3(n854), .A4(n1035), .Y(n1034) );
  AO22X1_LVT U931 ( .A1(n853), .A2(A[23]), .A3(n852), .A4(A[15]), .Y(n1035) );
  AO22X1_LVT U932 ( .A1(n853), .A2(A[39]), .A3(n852), .A4(A[31]), .Y(n995) );
  AO22X1_LVT U933 ( .A1(SH[4]), .A2(n996), .A3(n854), .A4(n994), .Y(n937) );
  AO22X1_LVT U934 ( .A1(n853), .A2(A[55]), .A3(n852), .A4(A[47]), .Y(n994) );
  AO22X1_LVT U935 ( .A1(n853), .A2(A[71]), .A3(n852), .A4(A[63]), .Y(n996) );
  AO22X1_LVT U936 ( .A1(SH[5]), .A2(n940), .A3(n855), .A4(n1036), .Y(B[14]) );
  AO22X1_LVT U937 ( .A1(SH[4]), .A2(n999), .A3(n854), .A4(n1037), .Y(n1036) );
  AO22X1_LVT U938 ( .A1(n853), .A2(A[22]), .A3(n852), .A4(A[14]), .Y(n1037) );
  AO22X1_LVT U939 ( .A1(n853), .A2(A[38]), .A3(n852), .A4(A[30]), .Y(n999) );
  AO22X1_LVT U940 ( .A1(SH[4]), .A2(n1000), .A3(n854), .A4(n998), .Y(n940) );
  AO22X1_LVT U941 ( .A1(n853), .A2(A[54]), .A3(n852), .A4(A[46]), .Y(n998) );
  AO22X1_LVT U942 ( .A1(n853), .A2(A[70]), .A3(n852), .A4(A[62]), .Y(n1000) );
  AO22X1_LVT U943 ( .A1(SH[5]), .A2(n943), .A3(n855), .A4(n1038), .Y(B[13]) );
  AO22X1_LVT U944 ( .A1(SH[4]), .A2(n1006), .A3(n854), .A4(n1039), .Y(n1038)
         );
  AO22X1_LVT U945 ( .A1(n853), .A2(A[21]), .A3(n852), .A4(A[13]), .Y(n1039) );
  AO22X1_LVT U946 ( .A1(n853), .A2(A[37]), .A3(n852), .A4(A[29]), .Y(n1006) );
  AO22X1_LVT U947 ( .A1(SH[4]), .A2(n1007), .A3(n854), .A4(n1005), .Y(n943) );
  AO22X1_LVT U948 ( .A1(n853), .A2(A[53]), .A3(n852), .A4(A[45]), .Y(n1005) );
  AO22X1_LVT U949 ( .A1(n853), .A2(A[69]), .A3(n852), .A4(A[61]), .Y(n1007) );
  AO22X1_LVT U950 ( .A1(n853), .A2(A[36]), .A3(n852), .A4(A[28]), .Y(n1010) );
  AO22X1_LVT U951 ( .A1(SH[4]), .A2(n1011), .A3(n854), .A4(n1009), .Y(n946) );
  AO22X1_LVT U952 ( .A1(n853), .A2(A[52]), .A3(n852), .A4(A[44]), .Y(n1009) );
  AO22X1_LVT U953 ( .A1(n853), .A2(A[68]), .A3(n852), .A4(A[60]), .Y(n1011) );
  AO22X1_LVT U954 ( .A1(SH[5]), .A2(n949), .A3(n855), .A4(n1040), .Y(B[11]) );
  AO22X1_LVT U955 ( .A1(SH[4]), .A2(n1014), .A3(n854), .A4(n1041), .Y(n1040)
         );
  AO22X1_LVT U956 ( .A1(n853), .A2(A[19]), .A3(n852), .A4(A[11]), .Y(n1041) );
  AO22X1_LVT U957 ( .A1(n853), .A2(A[35]), .A3(n852), .A4(A[27]), .Y(n1014) );
  AO22X1_LVT U958 ( .A1(SH[4]), .A2(n1015), .A3(n854), .A4(n1013), .Y(n949) );
  AO22X1_LVT U959 ( .A1(n853), .A2(A[51]), .A3(n852), .A4(A[43]), .Y(n1013) );
  AO22X1_LVT U960 ( .A1(n853), .A2(A[67]), .A3(n852), .A4(A[59]), .Y(n1015) );
  AO22X1_LVT U961 ( .A1(SH[5]), .A2(n952), .A3(n855), .A4(n1042), .Y(B[10]) );
  AO22X1_LVT U962 ( .A1(SH[4]), .A2(n1018), .A3(n854), .A4(n1043), .Y(n1042)
         );
  AO22X1_LVT U963 ( .A1(n853), .A2(A[18]), .A3(n852), .A4(A[10]), .Y(n1043) );
  AO22X1_LVT U964 ( .A1(n853), .A2(A[34]), .A3(n852), .A4(A[26]), .Y(n1018) );
  AO22X1_LVT U965 ( .A1(SH[4]), .A2(n1019), .A3(n854), .A4(n1017), .Y(n952) );
  AO22X1_LVT U966 ( .A1(n853), .A2(A[50]), .A3(n852), .A4(A[42]), .Y(n1017) );
  AO22X1_LVT U967 ( .A1(n853), .A2(A[66]), .A3(n852), .A4(A[58]), .Y(n1019) );
  AO22X1_LVT U968 ( .A1(n853), .A2(A[24]), .A3(n852), .A4(A[16]), .Y(n1032) );
  AO22X1_LVT U969 ( .A1(SH[4]), .A2(n1033), .A3(n854), .A4(n1031), .Y(n991) );
  AO22X1_LVT U970 ( .A1(n853), .A2(A[40]), .A3(n852), .A4(A[32]), .Y(n1031) );
  AO22X1_LVT U971 ( .A1(n853), .A2(A[56]), .A3(n852), .A4(A[48]), .Y(n1033) );
endmodule


module MulDiv_DW01_sub_J39_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   n161, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465;

  HADDX1_LVT U223 ( .A0(n389), .B0(n390), .C1(n161), .SO(DIFF[1]) );
  AO22X1_LVT U229 ( .A1(B[56]), .A2(n362), .A3(n402), .A4(n361), .Y(DIFF[56])
         );
  AO22X1_LVT U230 ( .A1(B[48]), .A2(n408), .A3(n365), .A4(n366), .Y(DIFF[48])
         );
  AO22X1_LVT U231 ( .A1(n461), .A2(n381), .A3(n382), .A4(B[12]), .Y(DIFF[12])
         );
  AO22X1_LVT U232 ( .A1(B[40]), .A2(n371), .A3(n422), .A4(n370), .Y(DIFF[40])
         );
  AO22X1_LVT U233 ( .A1(B[24]), .A2(n378), .A3(n445), .A4(n377), .Y(DIFF[24])
         );
  AO22X1_LVT U234 ( .A1(B[2]), .A2(n161), .A3(n387), .A4(n388), .Y(DIFF[2]) );
  AO22X1_LVT U235 ( .A1(B[16]), .A2(n380), .A3(n453), .A4(n379), .Y(DIFF[16])
         );
  AO22X1_LVT U236 ( .A1(B[4]), .A2(n386), .A3(n412), .A4(n385), .Y(DIFF[4]) );
  AO22X1_LVT U237 ( .A1(B[32]), .A2(n424), .A3(n372), .A4(n373), .Y(DIFF[32])
         );
  AO22X1_LVT U238 ( .A1(B[52]), .A2(n364), .A3(n406), .A4(n363), .Y(DIFF[52])
         );
  NOR4X1_LVT U239 ( .A1(B[9]), .A2(B[8]), .A3(B[11]), .A4(B[10]), .Y(n463) );
  INVX0_LVT U240 ( .A(n406), .Y(n364) );
  INVX0_LVT U241 ( .A(n461), .Y(n382) );
  INVX0_LVT U242 ( .A(B[2]), .Y(n387) );
  INVX0_LVT U243 ( .A(B[0]), .Y(n390) );
  INVX0_LVT U244 ( .A(B[1]), .Y(n389) );
  INVX0_LVT U245 ( .A(B[16]), .Y(n379) );
  INVX0_LVT U246 ( .A(B[40]), .Y(n370) );
  INVX0_LVT U247 ( .A(B[8]), .Y(n383) );
  INVX0_LVT U248 ( .A(B[56]), .Y(n361) );
  INVX0_LVT U249 ( .A(B[52]), .Y(n363) );
  INVX0_LVT U250 ( .A(B[12]), .Y(n381) );
  INVX0_LVT U251 ( .A(B[44]), .Y(n369) );
  INVX0_LVT U252 ( .A(B[46]), .Y(n367) );
  INVX0_LVT U253 ( .A(B[48]), .Y(n365) );
  INVX0_LVT U254 ( .A(B[4]), .Y(n385) );
  INVX0_LVT U255 ( .A(B[28]), .Y(n376) );
  INVX0_LVT U256 ( .A(B[24]), .Y(n377) );
  INVX0_LVT U257 ( .A(B[32]), .Y(n372) );
  INVX0_LVT U258 ( .A(B[30]), .Y(n374) );
  NOR4X1_LVT U259 ( .A1(B[49]), .A2(B[48]), .A3(B[51]), .A4(B[50]), .Y(n409)
         );
  NOR4X1_LVT U260 ( .A1(B[46]), .A2(B[47]), .A3(n414), .A4(n415), .Y(n408) );
  NOR4X1_LVT U261 ( .A1(B[38]), .A2(B[39]), .A3(n426), .A4(n427), .Y(n425) );
  NOR4X1_LVT U262 ( .A1(B[30]), .A2(B[31]), .A3(n437), .A4(n438), .Y(n424) );
  NOR4X1_LVT U263 ( .A1(B[22]), .A2(B[23]), .A3(n448), .A4(n449), .Y(n447) );
  NOR4X1_LVT U264 ( .A1(B[25]), .A2(B[24]), .A3(B[27]), .A4(B[26]), .Y(n440)
         );
  NOR4X1_LVT U265 ( .A1(B[41]), .A2(B[40]), .A3(B[43]), .A4(B[42]), .Y(n417)
         );
  INVX1_LVT U266 ( .A(n402), .Y(n362) );
  INVX1_LVT U267 ( .A(n408), .Y(n366) );
  INVX1_LVT U268 ( .A(n414), .Y(n368) );
  INVX1_LVT U269 ( .A(n422), .Y(n371) );
  INVX1_LVT U270 ( .A(n424), .Y(n373) );
  INVX1_LVT U271 ( .A(n437), .Y(n375) );
  INVX1_LVT U272 ( .A(n445), .Y(n378) );
  INVX1_LVT U273 ( .A(n453), .Y(n380) );
  INVX1_LVT U274 ( .A(n392), .Y(n384) );
  INVX1_LVT U275 ( .A(n412), .Y(n386) );
  INVX1_LVT U276 ( .A(n161), .Y(n388) );
  HADDX1_LVT U277 ( .A0(B[9]), .B0(n391), .SO(DIFF[9]) );
  NAND2X0_LVT U278 ( .A1(n384), .A2(n383), .Y(n391) );
  AO22X1_LVT U279 ( .A1(n384), .A2(B[8]), .A3(n392), .A4(n383), .Y(DIFF[8]) );
  HADDX1_LVT U280 ( .A0(B[7]), .B0(n393), .SO(DIFF[7]) );
  OR2X1_LVT U281 ( .A1(B[6]), .A2(n394), .Y(n393) );
  HADDX1_LVT U282 ( .A0(B[6]), .B0(n394), .SO(DIFF[6]) );
  HADDX1_LVT U283 ( .A0(n395), .B0(B[63]), .SO(DIFF[63]) );
  OR2X1_LVT U284 ( .A1(B[62]), .A2(n396), .Y(n395) );
  HADDX1_LVT U285 ( .A0(B[62]), .B0(n396), .SO(DIFF[62]) );
  OR3X1_LVT U286 ( .A1(B[61]), .A2(B[60]), .A3(n397), .Y(n396) );
  HADDX1_LVT U287 ( .A0(B[61]), .B0(n398), .SO(DIFF[61]) );
  OR2X1_LVT U288 ( .A1(B[60]), .A2(n397), .Y(n398) );
  HADDX1_LVT U289 ( .A0(B[60]), .B0(n397), .SO(DIFF[60]) );
  OR3X1_LVT U290 ( .A1(B[59]), .A2(B[58]), .A3(n399), .Y(n397) );
  HADDX1_LVT U291 ( .A0(n400), .B0(B[5]), .SO(DIFF[5]) );
  NAND2X0_LVT U292 ( .A1(n385), .A2(n386), .Y(n400) );
  HADDX1_LVT U293 ( .A0(B[59]), .B0(n401), .SO(DIFF[59]) );
  OR2X1_LVT U294 ( .A1(B[58]), .A2(n399), .Y(n401) );
  HADDX1_LVT U295 ( .A0(B[58]), .B0(n399), .SO(DIFF[58]) );
  OR3X1_LVT U296 ( .A1(B[57]), .A2(B[56]), .A3(n402), .Y(n399) );
  HADDX1_LVT U297 ( .A0(n403), .B0(B[57]), .SO(DIFF[57]) );
  NAND2X0_LVT U298 ( .A1(n361), .A2(n362), .Y(n403) );
  OR3X1_LVT U299 ( .A1(B[55]), .A2(B[54]), .A3(n404), .Y(n402) );
  HADDX1_LVT U300 ( .A0(n405), .B0(B[55]), .SO(DIFF[55]) );
  OR2X1_LVT U301 ( .A1(B[54]), .A2(n404), .Y(n405) );
  HADDX1_LVT U302 ( .A0(B[54]), .B0(n404), .SO(DIFF[54]) );
  OR3X1_LVT U303 ( .A1(B[53]), .A2(B[52]), .A3(n406), .Y(n404) );
  HADDX1_LVT U304 ( .A0(n407), .B0(B[53]), .SO(DIFF[53]) );
  NAND2X0_LVT U305 ( .A1(n363), .A2(n364), .Y(n407) );
  NAND2X0_LVT U306 ( .A1(n408), .A2(n409), .Y(n406) );
  HADDX1_LVT U307 ( .A0(n410), .B0(B[51]), .SO(DIFF[51]) );
  OR2X1_LVT U308 ( .A1(B[50]), .A2(n411), .Y(n410) );
  HADDX1_LVT U309 ( .A0(B[50]), .B0(n411), .SO(DIFF[50]) );
  OR3X1_LVT U310 ( .A1(B[49]), .A2(B[48]), .A3(n366), .Y(n411) );
  HADDX1_LVT U311 ( .A0(B[49]), .B0(n413), .SO(DIFF[49]) );
  NAND2X0_LVT U312 ( .A1(n408), .A2(n365), .Y(n413) );
  HADDX1_LVT U313 ( .A0(B[47]), .B0(n416), .SO(DIFF[47]) );
  NAND4X0_LVT U314 ( .A1(n368), .A2(n417), .A3(n371), .A4(n367), .Y(n416) );
  HADDX1_LVT U315 ( .A0(B[46]), .B0(n418), .SO(DIFF[46]) );
  NAND3X0_LVT U316 ( .A1(n417), .A2(n368), .A3(n371), .Y(n418) );
  OR2X1_LVT U317 ( .A1(B[45]), .A2(B[44]), .Y(n414) );
  HADDX1_LVT U318 ( .A0(B[45]), .B0(n419), .SO(DIFF[45]) );
  NAND3X0_LVT U319 ( .A1(n417), .A2(n371), .A3(n369), .Y(n419) );
  HADDX1_LVT U320 ( .A0(B[44]), .B0(n415), .SO(DIFF[44]) );
  NAND2X0_LVT U321 ( .A1(n417), .A2(n371), .Y(n415) );
  HADDX1_LVT U322 ( .A0(n420), .B0(B[43]), .SO(DIFF[43]) );
  OR2X1_LVT U323 ( .A1(B[42]), .A2(n421), .Y(n420) );
  HADDX1_LVT U324 ( .A0(B[42]), .B0(n421), .SO(DIFF[42]) );
  OR3X1_LVT U325 ( .A1(B[41]), .A2(B[40]), .A3(n422), .Y(n421) );
  HADDX1_LVT U326 ( .A0(B[41]), .B0(n423), .SO(DIFF[41]) );
  NAND2X0_LVT U327 ( .A1(n371), .A2(n370), .Y(n423) );
  NAND2X0_LVT U328 ( .A1(n424), .A2(n425), .Y(n422) );
  HADDX1_LVT U329 ( .A0(B[3]), .B0(n428), .SO(DIFF[3]) );
  NAND2X0_LVT U330 ( .A1(n161), .A2(n387), .Y(n428) );
  HADDX1_LVT U331 ( .A0(B[39]), .B0(n429), .SO(DIFF[39]) );
  OR3X1_LVT U332 ( .A1(B[38]), .A2(n427), .A3(n430), .Y(n429) );
  HADDX1_LVT U333 ( .A0(B[38]), .B0(n431), .SO(DIFF[38]) );
  OR3X1_LVT U334 ( .A1(n373), .A2(n426), .A3(n427), .Y(n431) );
  OR2X1_LVT U335 ( .A1(B[37]), .A2(B[36]), .Y(n427) );
  HADDX1_LVT U336 ( .A0(n432), .B0(B[37]), .SO(DIFF[37]) );
  OR2X1_LVT U337 ( .A1(B[36]), .A2(n430), .Y(n432) );
  HADDX1_LVT U338 ( .A0(B[36]), .B0(n430), .SO(DIFF[36]) );
  OR2X1_LVT U339 ( .A1(n373), .A2(n426), .Y(n430) );
  OR3X1_LVT U340 ( .A1(B[35]), .A2(B[34]), .A3(n433), .Y(n426) );
  HADDX1_LVT U341 ( .A0(B[35]), .B0(n434), .SO(DIFF[35]) );
  OR3X1_LVT U342 ( .A1(B[34]), .A2(n433), .A3(n373), .Y(n434) );
  HADDX1_LVT U343 ( .A0(B[34]), .B0(n435), .SO(DIFF[34]) );
  OR2X1_LVT U344 ( .A1(n373), .A2(n433), .Y(n435) );
  OR2X1_LVT U345 ( .A1(B[33]), .A2(B[32]), .Y(n433) );
  HADDX1_LVT U346 ( .A0(B[33]), .B0(n436), .SO(DIFF[33]) );
  NAND2X0_LVT U347 ( .A1(n424), .A2(n372), .Y(n436) );
  HADDX1_LVT U348 ( .A0(B[31]), .B0(n439), .SO(DIFF[31]) );
  NAND4X0_LVT U349 ( .A1(n375), .A2(n440), .A3(n378), .A4(n374), .Y(n439) );
  HADDX1_LVT U350 ( .A0(B[30]), .B0(n441), .SO(DIFF[30]) );
  NAND3X0_LVT U351 ( .A1(n440), .A2(n375), .A3(n378), .Y(n441) );
  OR2X1_LVT U352 ( .A1(B[29]), .A2(B[28]), .Y(n437) );
  HADDX1_LVT U353 ( .A0(B[29]), .B0(n442), .SO(DIFF[29]) );
  NAND3X0_LVT U354 ( .A1(n440), .A2(n378), .A3(n376), .Y(n442) );
  HADDX1_LVT U355 ( .A0(B[28]), .B0(n438), .SO(DIFF[28]) );
  NAND2X0_LVT U356 ( .A1(n440), .A2(n378), .Y(n438) );
  HADDX1_LVT U357 ( .A0(n443), .B0(B[27]), .SO(DIFF[27]) );
  OR2X1_LVT U358 ( .A1(B[26]), .A2(n444), .Y(n443) );
  HADDX1_LVT U359 ( .A0(B[26]), .B0(n444), .SO(DIFF[26]) );
  OR3X1_LVT U360 ( .A1(B[25]), .A2(B[24]), .A3(n445), .Y(n444) );
  HADDX1_LVT U361 ( .A0(B[25]), .B0(n446), .SO(DIFF[25]) );
  NAND2X0_LVT U362 ( .A1(n378), .A2(n377), .Y(n446) );
  NAND2X0_LVT U363 ( .A1(n380), .A2(n447), .Y(n445) );
  HADDX1_LVT U364 ( .A0(B[23]), .B0(n450), .SO(DIFF[23]) );
  OR3X1_LVT U365 ( .A1(B[22]), .A2(n449), .A3(n451), .Y(n450) );
  HADDX1_LVT U366 ( .A0(B[22]), .B0(n452), .SO(DIFF[22]) );
  OR3X1_LVT U367 ( .A1(n453), .A2(n448), .A3(n449), .Y(n452) );
  OR2X1_LVT U368 ( .A1(B[21]), .A2(B[20]), .Y(n449) );
  HADDX1_LVT U369 ( .A0(n454), .B0(B[21]), .SO(DIFF[21]) );
  OR2X1_LVT U370 ( .A1(B[20]), .A2(n451), .Y(n454) );
  HADDX1_LVT U371 ( .A0(B[20]), .B0(n451), .SO(DIFF[20]) );
  OR2X1_LVT U372 ( .A1(n453), .A2(n448), .Y(n451) );
  OR3X1_LVT U373 ( .A1(B[19]), .A2(B[18]), .A3(n455), .Y(n448) );
  HADDX1_LVT U374 ( .A0(B[19]), .B0(n456), .SO(DIFF[19]) );
  OR3X1_LVT U375 ( .A1(B[18]), .A2(n455), .A3(n453), .Y(n456) );
  HADDX1_LVT U376 ( .A0(B[18]), .B0(n457), .SO(DIFF[18]) );
  OR2X1_LVT U377 ( .A1(n453), .A2(n455), .Y(n457) );
  OR2X1_LVT U378 ( .A1(B[17]), .A2(B[16]), .Y(n455) );
  HADDX1_LVT U379 ( .A0(B[17]), .B0(n458), .SO(DIFF[17]) );
  NAND2X0_LVT U380 ( .A1(n380), .A2(n379), .Y(n458) );
  OR3X1_LVT U381 ( .A1(B[15]), .A2(B[14]), .A3(n459), .Y(n453) );
  HADDX1_LVT U382 ( .A0(n460), .B0(B[15]), .SO(DIFF[15]) );
  OR2X1_LVT U383 ( .A1(B[14]), .A2(n459), .Y(n460) );
  HADDX1_LVT U384 ( .A0(B[14]), .B0(n459), .SO(DIFF[14]) );
  OR3X1_LVT U385 ( .A1(B[13]), .A2(B[12]), .A3(n461), .Y(n459) );
  HADDX1_LVT U386 ( .A0(n462), .B0(B[13]), .SO(DIFF[13]) );
  NAND2X0_LVT U387 ( .A1(n381), .A2(n382), .Y(n462) );
  NAND2X0_LVT U388 ( .A1(n384), .A2(n463), .Y(n461) );
  HADDX1_LVT U389 ( .A0(n464), .B0(B[11]), .SO(DIFF[11]) );
  OR2X1_LVT U390 ( .A1(B[10]), .A2(n465), .Y(n464) );
  HADDX1_LVT U391 ( .A0(B[10]), .B0(n465), .SO(DIFF[10]) );
  OR3X1_LVT U392 ( .A1(B[9]), .A2(B[8]), .A3(n392), .Y(n465) );
  OR3X1_LVT U393 ( .A1(B[7]), .A2(B[6]), .A3(n394), .Y(n392) );
  OR3X1_LVT U394 ( .A1(B[5]), .A2(B[4]), .A3(n412), .Y(n394) );
  OR3X1_LVT U395 ( .A1(B[3]), .A2(B[2]), .A3(n388), .Y(n412) );
endmodule


module MulDiv_DW01_sub_J39_3 ( A, B, CI, DIFF, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] DIFF;
  input CI;
  output CO;
  wire   n782, n783, n784, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n810, n811, n812, n813, n815, n816, n817, n818,
         n819, n820, n822, n823, n824, n825, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;

  AO222X1_LVT U649 ( .A1(n815), .A2(n817), .A3(n818), .A4(n819), .A5(n820), 
        .A6(1'b1), .Y(n1041) );
  OA221X1_LVT U650 ( .A1(1'b0), .A2(n823), .A3(n1067), .A4(n824), .A5(n825), 
        .Y(n1037) );
  OA221X1_LVT U651 ( .A1(1'b0), .A2(n811), .A3(n1013), .A4(n812), .A5(n813), 
        .Y(n980) );
  OA221X1_LVT U652 ( .A1(1'b0), .A2(n805), .A3(n1038), .A4(n806), .A5(n808), 
        .Y(n810) );
  OA221X1_LVT U653 ( .A1(1'b0), .A2(n793), .A3(n921), .A4(n794), .A5(n796), 
        .Y(n798) );
  OA221X1_LVT U654 ( .A1(1'b0), .A2(n798), .A3(n920), .A4(n799), .A5(n800), 
        .Y(n917) );
  OA221X1_LVT U655 ( .A1(1'b0), .A2(n786), .A3(n951), .A4(n787), .A5(n788), 
        .Y(n921) );
  INVX0_LVT U656 ( .A(n906), .Y(n782) );
  INVX0_LVT U657 ( .A(B[2]), .Y(n783) );
  AO222X1_LVT U658 ( .A1(n783), .A2(n782), .A3(n1050), .A4(n1049), .A5(A[1]), 
        .A6(n876), .Y(n784) );
  OA21X1_LVT U659 ( .A1(n782), .A2(n783), .A3(n784), .Y(n977) );
  AO222X1_LVT U661 ( .A1(B[54]), .A2(n885), .A3(B[54]), .A4(n956), .A5(n885), 
        .A6(n956), .Y(n786) );
  NAND2X0_LVT U662 ( .A1(n954), .A2(n955), .Y(n787) );
  NAND2X0_LVT U663 ( .A1(n953), .A2(n952), .Y(n788) );
  INVX0_LVT U664 ( .A(A[62]), .Y(n789) );
  AO22X1_LVT U665 ( .A1(B[61]), .A2(n879), .A3(B[62]), .A4(n789), .Y(n790) );
  INVX0_LVT U666 ( .A(n790), .Y(n791) );
  NAND3X0_LVT U667 ( .A1(n927), .A2(n926), .A3(n791), .Y(n792) );
  OA22X1_LVT U668 ( .A1(n923), .A2(n790), .A3(n922), .A4(n792), .Y(n793) );
  OR2X1_LVT U669 ( .A1(n925), .A2(n792), .Y(n794) );
  OR2X1_LVT U670 ( .A1(B[61]), .A2(n879), .Y(n795) );
  AO222X1_LVT U671 ( .A1(B[62]), .A2(n789), .A3(B[62]), .A4(n795), .A5(n789), 
        .A6(n795), .Y(n796) );
  OR2X1_LVT U673 ( .A1(n924), .A2(n794), .Y(n799) );
  OR3X1_LVT U674 ( .A1(n918), .A2(n919), .A3(n799), .Y(n800) );
  NAND2X0_LVT U675 ( .A1(B[30]), .A2(n895), .Y(n801) );
  AND4X1_LVT U676 ( .A1(n1045), .A2(n1044), .A3(n1040), .A4(n801), .Y(n802) );
  NAND2X0_LVT U677 ( .A1(n802), .A2(n1043), .Y(n803) );
  NAND2X0_LVT U678 ( .A1(n1041), .A2(n1042), .Y(n804) );
  NAND2X0_LVT U679 ( .A1(n802), .A2(n1039), .Y(n805) );
  NAND2X0_LVT U680 ( .A1(n1040), .A2(n801), .Y(n806) );
  NAND2X0_LVT U681 ( .A1(n856), .A2(A[29]), .Y(n807) );
  AO222X1_LVT U682 ( .A1(B[30]), .A2(n895), .A3(B[30]), .A4(n807), .A5(n895), 
        .A6(n807), .Y(n808) );
  OA221X1_LVT U684 ( .A1(n803), .A2(n1037), .A3(n803), .A4(n804), .A5(n810), 
        .Y(n918) );
  AO222X1_LVT U685 ( .A1(B[38]), .A2(n891), .A3(B[38]), .A4(n1019), .A5(n891), 
        .A6(n1019), .Y(n811) );
  NAND2X0_LVT U686 ( .A1(n1015), .A2(n1016), .Y(n812) );
  NAND2X0_LVT U687 ( .A1(n1014), .A2(n1011), .Y(n813) );
  INVX0_LVT U689 ( .A(n1093), .Y(n815) );
  INVX0_LVT U690 ( .A(A[14]), .Y(n816) );
  AOI22X1_LVT U691 ( .A1(n899), .A2(B[13]), .A3(B[14]), .A4(n816), .Y(n817) );
  AO21X1_LVT U692 ( .A1(n872), .A2(n1092), .A3(n1094), .Y(n818) );
  AND3X1_LVT U693 ( .A1(n1096), .A2(n817), .A3(n1095), .Y(n819) );
  OAI222X1_LVT U694 ( .A1(n816), .A2(B[14]), .A3(n816), .A4(n1097), .A5(B[14]), 
        .A6(n1097), .Y(n820) );
  NAND2X0_LVT U696 ( .A1(n862), .A2(A[21]), .Y(n822) );
  AO222X1_LVT U697 ( .A1(B[22]), .A2(n897), .A3(B[22]), .A4(n822), .A5(n897), 
        .A6(n822), .Y(n823) );
  NAND2X0_LVT U698 ( .A1(n1070), .A2(n1071), .Y(n824) );
  NAND2X0_LVT U699 ( .A1(n1069), .A2(n1068), .Y(n825) );
  OR2X1_LVT U701 ( .A1(n981), .A2(n980), .Y(n827) );
  INVX0_LVT U702 ( .A(n982), .Y(n828) );
  NAND3X0_LVT U703 ( .A1(n986), .A2(n985), .A3(n828), .Y(n829) );
  NAND2X0_LVT U704 ( .A1(n983), .A2(n984), .Y(n830) );
  AO222X1_LVT U705 ( .A1(B[46]), .A2(n888), .A3(B[46]), .A4(n987), .A5(n888), 
        .A6(n987), .Y(n831) );
  AND4X1_LVT U706 ( .A1(n827), .A2(n829), .A3(n830), .A4(n831), .Y(n920) );
  NAND2X0_LVT U707 ( .A1(n1041), .A2(n1042), .Y(n832) );
  NAND2X0_LVT U708 ( .A1(n1037), .A2(n832), .Y(n1055) );
  INVX0_LVT U709 ( .A(n950), .Y(n835) );
  INVX0_LVT U710 ( .A(n918), .Y(n834) );
  INVX0_LVT U711 ( .A(n912), .Y(n872) );
  INVX0_LVT U712 ( .A(n977), .Y(n875) );
  INVX0_LVT U713 ( .A(n981), .Y(n844) );
  INVX0_LVT U714 ( .A(n964), .Y(n838) );
  INVX0_LVT U715 ( .A(n996), .Y(n845) );
  INVX0_LVT U716 ( .A(n1102), .Y(n868) );
  INVX0_LVT U717 ( .A(n1024), .Y(n851) );
  NOR2X1_LVT U718 ( .A1(n894), .A2(B[31]), .Y(n1035) );
  NOR2X1_LVT U719 ( .A1(n902), .A2(B[7]), .Y(n911) );
  INVX0_LVT U720 ( .A(A[20]), .Y(n898) );
  INVX0_LVT U721 ( .A(A[28]), .Y(n896) );
  INVX0_LVT U722 ( .A(A[30]), .Y(n895) );
  INVX0_LVT U723 ( .A(A[31]), .Y(n894) );
  INVX0_LVT U724 ( .A(A[13]), .Y(n899) );
  INVX0_LVT U725 ( .A(A[12]), .Y(n900) );
  INVX0_LVT U726 ( .A(B[0]), .Y(n877) );
  INVX0_LVT U727 ( .A(A[4]), .Y(n904) );
  INVX0_LVT U728 ( .A(B[1]), .Y(n876) );
  INVX0_LVT U729 ( .A(A[2]), .Y(n906) );
  INVX0_LVT U730 ( .A(A[1]), .Y(n907) );
  INVX0_LVT U731 ( .A(A[3]), .Y(n905) );
  INVX0_LVT U732 ( .A(A[6]), .Y(n903) );
  INVX0_LVT U733 ( .A(A[7]), .Y(n902) );
  INVX0_LVT U734 ( .A(A[9]), .Y(n901) );
  INVX0_LVT U735 ( .A(A[63]), .Y(n878) );
  INVX0_LVT U736 ( .A(A[22]), .Y(n897) );
  INVX0_LVT U737 ( .A(A[54]), .Y(n885) );
  INVX0_LVT U738 ( .A(A[53]), .Y(n886) );
  INVX0_LVT U739 ( .A(A[52]), .Y(n887) );
  INVX0_LVT U740 ( .A(B[47]), .Y(n843) );
  INVX0_LVT U741 ( .A(A[58]), .Y(n881) );
  INVX0_LVT U742 ( .A(A[57]), .Y(n882) );
  INVX0_LVT U743 ( .A(A[56]), .Y(n883) );
  INVX0_LVT U744 ( .A(A[55]), .Y(n884) );
  INVX0_LVT U745 ( .A(A[61]), .Y(n879) );
  INVX0_LVT U746 ( .A(A[60]), .Y(n880) );
  INVX0_LVT U747 ( .A(B[59]), .Y(n837) );
  INVX0_LVT U748 ( .A(A[36]), .Y(n893) );
  INVX0_LVT U749 ( .A(A[38]), .Y(n891) );
  INVX0_LVT U750 ( .A(A[37]), .Y(n892) );
  INVX0_LVT U751 ( .A(A[44]), .Y(n890) );
  INVX0_LVT U752 ( .A(A[46]), .Y(n888) );
  INVX0_LVT U753 ( .A(A[45]), .Y(n889) );
  INVX1_LVT U754 ( .A(B[5]), .Y(n873) );
  INVX1_LVT U755 ( .A(B[8]), .Y(n871) );
  INVX1_LVT U756 ( .A(B[10]), .Y(n870) );
  INVX1_LVT U757 ( .A(B[11]), .Y(n869) );
  INVX1_LVT U758 ( .A(B[15]), .Y(n867) );
  INVX1_LVT U759 ( .A(B[21]), .Y(n862) );
  INVX1_LVT U760 ( .A(B[27]), .Y(n857) );
  INVX1_LVT U761 ( .A(B[29]), .Y(n856) );
  INVX1_LVT U762 ( .A(B[24]), .Y(n860) );
  INVX1_LVT U763 ( .A(B[26]), .Y(n858) );
  INVX1_LVT U764 ( .A(A[0]), .Y(n833) );
  INVX1_LVT U765 ( .A(n927), .Y(n836) );
  INVX1_LVT U766 ( .A(B[51]), .Y(n839) );
  INVX1_LVT U767 ( .A(B[50]), .Y(n840) );
  INVX1_LVT U768 ( .A(B[49]), .Y(n841) );
  INVX1_LVT U769 ( .A(B[48]), .Y(n842) );
  INVX1_LVT U770 ( .A(B[43]), .Y(n846) );
  INVX1_LVT U771 ( .A(B[42]), .Y(n847) );
  INVX1_LVT U772 ( .A(B[41]), .Y(n848) );
  INVX1_LVT U773 ( .A(B[40]), .Y(n849) );
  INVX1_LVT U774 ( .A(B[39]), .Y(n850) );
  INVX1_LVT U775 ( .A(B[35]), .Y(n852) );
  INVX1_LVT U776 ( .A(B[34]), .Y(n853) );
  INVX1_LVT U777 ( .A(B[33]), .Y(n854) );
  INVX1_LVT U778 ( .A(B[32]), .Y(n855) );
  INVX1_LVT U779 ( .A(B[25]), .Y(n859) );
  INVX1_LVT U780 ( .A(B[23]), .Y(n861) );
  INVX1_LVT U781 ( .A(B[19]), .Y(n863) );
  INVX1_LVT U782 ( .A(B[18]), .Y(n864) );
  INVX1_LVT U783 ( .A(B[17]), .Y(n865) );
  INVX1_LVT U784 ( .A(B[16]), .Y(n866) );
  INVX1_LVT U785 ( .A(B[3]), .Y(n874) );
  FADDX1_LVT U786 ( .A(B[9]), .B(n901), .CI(n908), .S(DIFF[9]) );
  FADDX1_LVT U787 ( .A(A[8]), .B(n871), .CI(n909), .S(DIFF[8]) );
  AO21X1_LVT U788 ( .A1(n910), .A2(n872), .A3(n911), .Y(n909) );
  FADDX1_LVT U789 ( .A(A[7]), .B(B[7]), .CI(n912), .S(DIFF[7]) );
  FADDX1_LVT U790 ( .A(B[6]), .B(n903), .CI(n913), .S(DIFF[6]) );
  AO22X1_LVT U791 ( .A1(A[5]), .A2(n873), .A3(n914), .A4(n915), .Y(n913) );
  FADDX1_LVT U792 ( .A(B[64]), .B(A[64]), .CI(n916), .S(DIFF[64]) );
  AO222X1_LVT U793 ( .A1(B[63]), .A2(n878), .A3(B[63]), .A4(n917), .A5(n878), 
        .A6(n917), .Y(n916) );
  FADDX1_LVT U794 ( .A(A[63]), .B(B[63]), .CI(n917), .S(DIFF[63]) );
  FADDX1_LVT U795 ( .A(n928), .B(A[62]), .CI(B[62]), .S(DIFF[62]) );
  AO222X1_LVT U796 ( .A1(B[61]), .A2(n879), .A3(B[61]), .A4(n929), .A5(n879), 
        .A6(n929), .Y(n928) );
  FADDX1_LVT U797 ( .A(A[61]), .B(B[61]), .CI(n929), .S(DIFF[61]) );
  OA21X1_LVT U798 ( .A1(n930), .A2(n931), .A3(n923), .Y(n929) );
  AO222X1_LVT U799 ( .A1(B[60]), .A2(n880), .A3(B[60]), .A4(n932), .A5(n880), 
        .A6(n932), .Y(n923) );
  NAND2X0_LVT U800 ( .A1(n926), .A2(n927), .Y(n931) );
  NAND2X0_LVT U801 ( .A1(B[60]), .A2(n880), .Y(n926) );
  FADDX1_LVT U802 ( .A(A[60]), .B(B[60]), .CI(n933), .S(DIFF[60]) );
  OA21X1_LVT U803 ( .A1(n836), .A2(n930), .A3(n932), .Y(n933) );
  NAND2X0_LVT U804 ( .A1(A[59]), .A2(n837), .Y(n932) );
  OR2X1_LVT U805 ( .A1(n837), .A2(A[59]), .Y(n927) );
  FADDX1_LVT U806 ( .A(A[5]), .B(n914), .CI(n873), .S(DIFF[5]) );
  NAND2X0_LVT U807 ( .A1(n934), .A2(n935), .Y(n914) );
  FADDX1_LVT U808 ( .A(A[59]), .B(B[59]), .CI(n930), .S(DIFF[59]) );
  OA21X1_LVT U809 ( .A1(n936), .A2(n925), .A3(n922), .Y(n930) );
  OA21X1_LVT U810 ( .A1(n937), .A2(n938), .A3(n939), .Y(n922) );
  AO222X1_LVT U811 ( .A1(B[58]), .A2(n881), .A3(B[58]), .A4(n940), .A5(n881), 
        .A6(n940), .Y(n939) );
  NAND2X0_LVT U812 ( .A1(n941), .A2(n942), .Y(n938) );
  NAND4X0_LVT U813 ( .A1(n941), .A2(n942), .A3(n943), .A4(n944), .Y(n925) );
  NAND2X0_LVT U814 ( .A1(B[57]), .A2(n882), .Y(n942) );
  NAND2X0_LVT U815 ( .A1(B[58]), .A2(n881), .Y(n941) );
  FADDX1_LVT U816 ( .A(A[58]), .B(B[58]), .CI(n945), .S(DIFF[58]) );
  AO22X1_LVT U817 ( .A1(n946), .A2(n940), .A3(B[57]), .A4(n882), .Y(n945) );
  OR2X1_LVT U818 ( .A1(n882), .A2(B[57]), .Y(n940) );
  FADDX1_LVT U819 ( .A(A[57]), .B(B[57]), .CI(n946), .S(DIFF[57]) );
  OA21X1_LVT U820 ( .A1(n936), .A2(n947), .A3(n937), .Y(n946) );
  AO222X1_LVT U821 ( .A1(B[56]), .A2(n883), .A3(B[56]), .A4(n948), .A5(n883), 
        .A6(n948), .Y(n937) );
  NAND2X0_LVT U822 ( .A1(n943), .A2(n944), .Y(n947) );
  NAND2X0_LVT U823 ( .A1(B[55]), .A2(n884), .Y(n944) );
  NAND2X0_LVT U824 ( .A1(B[56]), .A2(n883), .Y(n943) );
  FADDX1_LVT U825 ( .A(A[56]), .B(B[56]), .CI(n949), .S(DIFF[56]) );
  AO22X1_LVT U826 ( .A1(n936), .A2(n948), .A3(B[55]), .A4(n884), .Y(n949) );
  OR2X1_LVT U827 ( .A1(n884), .A2(B[55]), .Y(n948) );
  FADDX1_LVT U828 ( .A(A[55]), .B(B[55]), .CI(n936), .S(DIFF[55]) );
  OA21X1_LVT U829 ( .A1(n950), .A2(n924), .A3(n921), .Y(n936) );
  NAND2X0_LVT U830 ( .A1(n952), .A2(n957), .Y(n924) );
  AND4X1_LVT U831 ( .A1(n954), .A2(n955), .A3(n958), .A4(n959), .Y(n952) );
  NAND2X0_LVT U832 ( .A1(B[53]), .A2(n886), .Y(n955) );
  NAND2X0_LVT U833 ( .A1(B[54]), .A2(n885), .Y(n954) );
  FADDX1_LVT U834 ( .A(A[54]), .B(B[54]), .CI(n960), .S(DIFF[54]) );
  AO22X1_LVT U835 ( .A1(n961), .A2(n956), .A3(B[53]), .A4(n886), .Y(n960) );
  OR2X1_LVT U836 ( .A1(n886), .A2(B[53]), .Y(n956) );
  FADDX1_LVT U837 ( .A(A[53]), .B(B[53]), .CI(n961), .S(DIFF[53]) );
  AND2X1_LVT U838 ( .A1(n951), .A2(n962), .Y(n961) );
  NAND3X0_LVT U839 ( .A1(n963), .A2(n958), .A3(n959), .Y(n962) );
  NAND2X0_LVT U840 ( .A1(B[52]), .A2(n887), .Y(n958) );
  AO222X1_LVT U841 ( .A1(B[52]), .A2(n887), .A3(B[52]), .A4(n964), .A5(n887), 
        .A6(n964), .Y(n951) );
  FADDX1_LVT U842 ( .A(B[52]), .B(n965), .CI(n887), .S(DIFF[52]) );
  OA21X1_LVT U843 ( .A1(n838), .A2(n963), .A3(n959), .Y(n965) );
  OR2X1_LVT U844 ( .A1(n839), .A2(A[51]), .Y(n959) );
  NAND2X0_LVT U845 ( .A1(A[51]), .A2(n839), .Y(n964) );
  FADDX1_LVT U846 ( .A(A[51]), .B(n839), .CI(n963), .S(DIFF[51]) );
  AO21X1_LVT U847 ( .A1(n957), .A2(n835), .A3(n953), .Y(n963) );
  AO222X1_LVT U848 ( .A1(A[50]), .A2(n840), .A3(n966), .A4(n967), .A5(n968), 
        .A6(n969), .Y(n953) );
  AND2X1_LVT U849 ( .A1(n967), .A2(n970), .Y(n968) );
  AND4X1_LVT U850 ( .A1(n967), .A2(n970), .A3(n971), .A4(n972), .Y(n957) );
  OR2X1_LVT U851 ( .A1(n840), .A2(A[50]), .Y(n967) );
  FADDX1_LVT U852 ( .A(A[50]), .B(n973), .CI(n840), .S(DIFF[50]) );
  OA21X1_LVT U853 ( .A1(n966), .A2(n974), .A3(n970), .Y(n973) );
  OR2X1_LVT U854 ( .A1(n841), .A2(A[49]), .Y(n970) );
  AND2X1_LVT U855 ( .A1(A[49]), .A2(n841), .Y(n966) );
  FADDX1_LVT U856 ( .A(A[4]), .B(B[4]), .CI(n975), .S(DIFF[4]) );
  AO22X1_LVT U857 ( .A1(B[3]), .A2(n905), .A3(n875), .A4(n976), .Y(n975) );
  FADDX1_LVT U858 ( .A(A[49]), .B(n841), .CI(n974), .S(DIFF[49]) );
  OA222X1_LVT U859 ( .A1(n969), .A2(n971), .A3(n969), .A4(n972), .A5(n969), 
        .A6(n835), .Y(n974) );
  AO22X1_LVT U860 ( .A1(A[48]), .A2(n842), .A3(n978), .A4(n971), .Y(n969) );
  OR2X1_LVT U861 ( .A1(n842), .A2(A[48]), .Y(n971) );
  FADDX1_LVT U862 ( .A(A[48]), .B(n979), .CI(n842), .S(DIFF[48]) );
  OA21X1_LVT U863 ( .A1(n978), .A2(n835), .A3(n972), .Y(n979) );
  OR2X1_LVT U864 ( .A1(n843), .A2(A[47]), .Y(n972) );
  AND2X1_LVT U865 ( .A1(A[47]), .A2(n843), .Y(n978) );
  FADDX1_LVT U866 ( .A(A[47]), .B(B[47]), .CI(n950), .S(DIFF[47]) );
  OA21X1_LVT U867 ( .A1(n918), .A2(n919), .A3(n920), .Y(n950) );
  NAND2X0_LVT U868 ( .A1(n844), .A2(n988), .Y(n919) );
  NAND2X0_LVT U869 ( .A1(n989), .A2(n983), .Y(n981) );
  AND4X1_LVT U870 ( .A1(n985), .A2(n986), .A3(n990), .A4(n991), .Y(n983) );
  NAND2X0_LVT U871 ( .A1(B[45]), .A2(n889), .Y(n986) );
  NAND2X0_LVT U872 ( .A1(B[46]), .A2(n888), .Y(n985) );
  FADDX1_LVT U873 ( .A(A[46]), .B(B[46]), .CI(n992), .S(DIFF[46]) );
  AO22X1_LVT U874 ( .A1(n993), .A2(n987), .A3(B[45]), .A4(n889), .Y(n992) );
  OR2X1_LVT U875 ( .A1(n889), .A2(B[45]), .Y(n987) );
  FADDX1_LVT U876 ( .A(A[45]), .B(B[45]), .CI(n993), .S(DIFF[45]) );
  AND2X1_LVT U877 ( .A1(n982), .A2(n994), .Y(n993) );
  NAND3X0_LVT U878 ( .A1(n995), .A2(n990), .A3(n991), .Y(n994) );
  NAND2X0_LVT U879 ( .A1(B[44]), .A2(n890), .Y(n990) );
  AO222X1_LVT U880 ( .A1(B[44]), .A2(n890), .A3(B[44]), .A4(n996), .A5(n890), 
        .A6(n996), .Y(n982) );
  FADDX1_LVT U881 ( .A(B[44]), .B(n997), .CI(n890), .S(DIFF[44]) );
  OA21X1_LVT U882 ( .A1(n845), .A2(n995), .A3(n991), .Y(n997) );
  OR2X1_LVT U883 ( .A1(n846), .A2(A[43]), .Y(n991) );
  NAND2X0_LVT U884 ( .A1(A[43]), .A2(n846), .Y(n996) );
  FADDX1_LVT U885 ( .A(A[43]), .B(n846), .CI(n995), .S(DIFF[43]) );
  AO21X1_LVT U886 ( .A1(n989), .A2(n998), .A3(n984), .Y(n995) );
  AO222X1_LVT U887 ( .A1(A[42]), .A2(n847), .A3(n999), .A4(n1000), .A5(n1001), 
        .A6(n1002), .Y(n984) );
  AND2X1_LVT U888 ( .A1(n1000), .A2(n1003), .Y(n1001) );
  AND4X1_LVT U889 ( .A1(n1000), .A2(n1003), .A3(n1004), .A4(n1005), .Y(n989)
         );
  OR2X1_LVT U890 ( .A1(n847), .A2(A[42]), .Y(n1000) );
  FADDX1_LVT U891 ( .A(A[42]), .B(n1006), .CI(n847), .S(DIFF[42]) );
  OA21X1_LVT U892 ( .A1(n999), .A2(n1007), .A3(n1003), .Y(n1006) );
  OR2X1_LVT U893 ( .A1(n848), .A2(A[41]), .Y(n1003) );
  AND2X1_LVT U894 ( .A1(A[41]), .A2(n848), .Y(n999) );
  FADDX1_LVT U895 ( .A(A[41]), .B(n848), .CI(n1007), .S(DIFF[41]) );
  OA222X1_LVT U896 ( .A1(n1002), .A2(n1004), .A3(n1002), .A4(n1005), .A5(n1002), .A6(n998), .Y(n1007) );
  AO22X1_LVT U897 ( .A1(A[40]), .A2(n849), .A3(n1008), .A4(n1004), .Y(n1002)
         );
  OR2X1_LVT U898 ( .A1(n849), .A2(A[40]), .Y(n1004) );
  FADDX1_LVT U899 ( .A(A[40]), .B(n1009), .CI(n849), .S(DIFF[40]) );
  OA21X1_LVT U900 ( .A1(n1008), .A2(n998), .A3(n1005), .Y(n1009) );
  OR2X1_LVT U901 ( .A1(n850), .A2(A[39]), .Y(n1005) );
  AND2X1_LVT U902 ( .A1(A[39]), .A2(n850), .Y(n1008) );
  FADDX1_LVT U903 ( .A(n977), .B(A[3]), .CI(n874), .S(DIFF[3]) );
  FADDX1_LVT U904 ( .A(A[39]), .B(n850), .CI(n998), .S(DIFF[39]) );
  NAND2X0_LVT U905 ( .A1(n980), .A2(n1010), .Y(n998) );
  NAND2X0_LVT U906 ( .A1(n988), .A2(n834), .Y(n1010) );
  AND2X1_LVT U907 ( .A1(n1011), .A2(n1012), .Y(n988) );
  AND4X1_LVT U908 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .Y(n1011)
         );
  NAND2X0_LVT U909 ( .A1(B[37]), .A2(n892), .Y(n1016) );
  NAND2X0_LVT U910 ( .A1(B[38]), .A2(n891), .Y(n1015) );
  FADDX1_LVT U911 ( .A(A[38]), .B(B[38]), .CI(n1020), .S(DIFF[38]) );
  AO22X1_LVT U912 ( .A1(n1021), .A2(n1019), .A3(B[37]), .A4(n892), .Y(n1020)
         );
  OR2X1_LVT U913 ( .A1(n892), .A2(B[37]), .Y(n1019) );
  FADDX1_LVT U914 ( .A(A[37]), .B(B[37]), .CI(n1021), .S(DIFF[37]) );
  AND2X1_LVT U915 ( .A1(n1013), .A2(n1022), .Y(n1021) );
  NAND3X0_LVT U916 ( .A1(n1023), .A2(n1017), .A3(n1018), .Y(n1022) );
  NAND2X0_LVT U917 ( .A1(B[36]), .A2(n893), .Y(n1017) );
  AO222X1_LVT U918 ( .A1(B[36]), .A2(n893), .A3(B[36]), .A4(n1024), .A5(n893), 
        .A6(n1024), .Y(n1013) );
  FADDX1_LVT U919 ( .A(B[36]), .B(n1025), .CI(n893), .S(DIFF[36]) );
  OA21X1_LVT U920 ( .A1(n851), .A2(n1023), .A3(n1018), .Y(n1025) );
  OR2X1_LVT U921 ( .A1(n852), .A2(A[35]), .Y(n1018) );
  NAND2X0_LVT U922 ( .A1(A[35]), .A2(n852), .Y(n1024) );
  FADDX1_LVT U923 ( .A(A[35]), .B(n852), .CI(n1023), .S(DIFF[35]) );
  AO21X1_LVT U924 ( .A1(n1012), .A2(n834), .A3(n1014), .Y(n1023) );
  AO222X1_LVT U925 ( .A1(A[34]), .A2(n853), .A3(n1026), .A4(n1027), .A5(n1028), 
        .A6(n1029), .Y(n1014) );
  AND2X1_LVT U926 ( .A1(n1027), .A2(n1030), .Y(n1028) );
  AND4X1_LVT U927 ( .A1(n1027), .A2(n1030), .A3(n1031), .A4(n1032), .Y(n1012)
         );
  OR2X1_LVT U928 ( .A1(n853), .A2(A[34]), .Y(n1027) );
  FADDX1_LVT U929 ( .A(A[34]), .B(n1033), .CI(n853), .S(DIFF[34]) );
  OA21X1_LVT U930 ( .A1(n1026), .A2(n1034), .A3(n1030), .Y(n1033) );
  OR2X1_LVT U931 ( .A1(n854), .A2(A[33]), .Y(n1030) );
  AND2X1_LVT U932 ( .A1(A[33]), .A2(n854), .Y(n1026) );
  FADDX1_LVT U933 ( .A(A[33]), .B(n854), .CI(n1034), .S(DIFF[33]) );
  OA222X1_LVT U934 ( .A1(n1029), .A2(n1031), .A3(n1029), .A4(n1032), .A5(n1029), .A6(n834), .Y(n1034) );
  AO22X1_LVT U935 ( .A1(A[32]), .A2(n855), .A3(n1035), .A4(n1031), .Y(n1029)
         );
  OR2X1_LVT U936 ( .A1(n855), .A2(A[32]), .Y(n1031) );
  FADDX1_LVT U937 ( .A(A[32]), .B(n855), .CI(n1036), .S(DIFF[32]) );
  AO21X1_LVT U938 ( .A1(n1032), .A2(n834), .A3(n1035), .Y(n1036) );
  NAND2X0_LVT U939 ( .A1(B[31]), .A2(n894), .Y(n1032) );
  FADDX1_LVT U940 ( .A(A[31]), .B(B[31]), .CI(n918), .S(DIFF[31]) );
  FADDX1_LVT U941 ( .A(B[30]), .B(n895), .CI(n1046), .S(DIFF[30]) );
  AO22X1_LVT U942 ( .A1(A[29]), .A2(n856), .A3(n1047), .A4(n1040), .Y(n1046)
         );
  OR2X1_LVT U943 ( .A1(n856), .A2(A[29]), .Y(n1040) );
  FADDX1_LVT U944 ( .A(B[2]), .B(n906), .CI(n1048), .S(DIFF[2]) );
  AO22X1_LVT U945 ( .A1(A[1]), .A2(n876), .A3(n1049), .A4(n1050), .Y(n1048) );
  FADDX1_LVT U946 ( .A(A[29]), .B(n1047), .CI(n856), .S(DIFF[29]) );
  NAND2X0_LVT U947 ( .A1(n1038), .A2(n1051), .Y(n1047) );
  NAND3X0_LVT U948 ( .A1(n1044), .A2(n1052), .A3(n1045), .Y(n1051) );
  NAND2X0_LVT U949 ( .A1(B[28]), .A2(n896), .Y(n1044) );
  AO222X1_LVT U950 ( .A1(B[28]), .A2(n896), .A3(B[28]), .A4(n1053), .A5(n896), 
        .A6(n1053), .Y(n1038) );
  NAND2X0_LVT U951 ( .A1(A[27]), .A2(n857), .Y(n1053) );
  FADDX1_LVT U952 ( .A(B[28]), .B(n896), .CI(n1054), .S(DIFF[28]) );
  AO22X1_LVT U953 ( .A1(A[27]), .A2(n857), .A3(n1052), .A4(n1045), .Y(n1054)
         );
  OR2X1_LVT U954 ( .A1(n857), .A2(A[27]), .Y(n1045) );
  FADDX1_LVT U955 ( .A(A[27]), .B(n1052), .CI(n857), .S(DIFF[27]) );
  AO21X1_LVT U956 ( .A1(n1043), .A2(n1055), .A3(n1039), .Y(n1052) );
  AO222X1_LVT U957 ( .A1(A[26]), .A2(n858), .A3(n1056), .A4(n1057), .A5(n1058), 
        .A6(n1059), .Y(n1039) );
  AND2X1_LVT U958 ( .A1(n1057), .A2(n1060), .Y(n1058) );
  AND4X1_LVT U959 ( .A1(n1057), .A2(n1060), .A3(n1061), .A4(n1062), .Y(n1043)
         );
  OR2X1_LVT U960 ( .A1(n858), .A2(A[26]), .Y(n1057) );
  FADDX1_LVT U961 ( .A(A[26]), .B(n858), .CI(n1063), .S(DIFF[26]) );
  AO21X1_LVT U962 ( .A1(n1064), .A2(n1060), .A3(n1056), .Y(n1063) );
  AND2X1_LVT U963 ( .A1(A[25]), .A2(n859), .Y(n1056) );
  OR2X1_LVT U964 ( .A1(n859), .A2(A[25]), .Y(n1060) );
  FADDX1_LVT U965 ( .A(A[25]), .B(n1064), .CI(n859), .S(DIFF[25]) );
  OA222X1_LVT U966 ( .A1(n1059), .A2(n1055), .A3(n1059), .A4(n1061), .A5(n1059), .A6(n1062), .Y(n1064) );
  AO22X1_LVT U967 ( .A1(A[24]), .A2(n860), .A3(n1065), .A4(n1061), .Y(n1059)
         );
  OR2X1_LVT U968 ( .A1(n860), .A2(A[24]), .Y(n1061) );
  FADDX1_LVT U969 ( .A(A[24]), .B(n860), .CI(n1066), .S(DIFF[24]) );
  AO21X1_LVT U970 ( .A1(n1055), .A2(n1062), .A3(n1065), .Y(n1066) );
  AND2X1_LVT U971 ( .A1(A[23]), .A2(n861), .Y(n1065) );
  OR2X1_LVT U972 ( .A1(n861), .A2(A[23]), .Y(n1062) );
  FADDX1_LVT U973 ( .A(A[23]), .B(n1055), .CI(n861), .S(DIFF[23]) );
  AND2X1_LVT U974 ( .A1(n1072), .A2(n1068), .Y(n1042) );
  AND4X1_LVT U975 ( .A1(n1070), .A2(n1071), .A3(n1073), .A4(n1074), .Y(n1068)
         );
  NAND2X0_LVT U976 ( .A1(B[22]), .A2(n897), .Y(n1070) );
  FADDX1_LVT U977 ( .A(B[22]), .B(n897), .CI(n1075), .S(DIFF[22]) );
  AO22X1_LVT U978 ( .A1(A[21]), .A2(n862), .A3(n1076), .A4(n1071), .Y(n1075)
         );
  OR2X1_LVT U979 ( .A1(n862), .A2(A[21]), .Y(n1071) );
  FADDX1_LVT U980 ( .A(A[21]), .B(n1076), .CI(n862), .S(DIFF[21]) );
  NAND2X0_LVT U981 ( .A1(n1067), .A2(n1077), .Y(n1076) );
  NAND3X0_LVT U982 ( .A1(n1073), .A2(n1078), .A3(n1074), .Y(n1077) );
  NAND2X0_LVT U983 ( .A1(B[20]), .A2(n898), .Y(n1073) );
  AO222X1_LVT U984 ( .A1(B[20]), .A2(n898), .A3(B[20]), .A4(n1079), .A5(n898), 
        .A6(n1079), .Y(n1067) );
  NAND2X0_LVT U985 ( .A1(A[19]), .A2(n863), .Y(n1079) );
  FADDX1_LVT U986 ( .A(B[20]), .B(n898), .CI(n1080), .S(DIFF[20]) );
  AO22X1_LVT U987 ( .A1(A[19]), .A2(n863), .A3(n1078), .A4(n1074), .Y(n1080)
         );
  OR2X1_LVT U988 ( .A1(n863), .A2(A[19]), .Y(n1074) );
  FADDX1_LVT U989 ( .A(B[1]), .B(n907), .CI(n1049), .S(DIFF[1]) );
  FADDX1_LVT U990 ( .A(A[19]), .B(n1078), .CI(n863), .S(DIFF[19]) );
  AO21X1_LVT U991 ( .A1(n1041), .A2(n1072), .A3(n1069), .Y(n1078) );
  AO222X1_LVT U992 ( .A1(A[18]), .A2(n864), .A3(n1081), .A4(n1082), .A5(n1083), 
        .A6(n1084), .Y(n1069) );
  AND2X1_LVT U993 ( .A1(n1082), .A2(n1085), .Y(n1083) );
  AND4X1_LVT U994 ( .A1(n1082), .A2(n1085), .A3(n1086), .A4(n1087), .Y(n1072)
         );
  OR2X1_LVT U995 ( .A1(n864), .A2(A[18]), .Y(n1082) );
  FADDX1_LVT U996 ( .A(A[18]), .B(n864), .CI(n1088), .S(DIFF[18]) );
  AO21X1_LVT U997 ( .A1(n1089), .A2(n1085), .A3(n1081), .Y(n1088) );
  AND2X1_LVT U998 ( .A1(A[17]), .A2(n865), .Y(n1081) );
  OR2X1_LVT U999 ( .A1(n865), .A2(A[17]), .Y(n1085) );
  FADDX1_LVT U1000 ( .A(A[17]), .B(n1089), .CI(n865), .S(DIFF[17]) );
  OA222X1_LVT U1001 ( .A1(n1084), .A2(n1041), .A3(n1084), .A4(n1086), .A5(
        n1084), .A6(n1087), .Y(n1089) );
  AO22X1_LVT U1002 ( .A1(A[16]), .A2(n866), .A3(n1090), .A4(n1086), .Y(n1084)
         );
  OR2X1_LVT U1003 ( .A1(n866), .A2(A[16]), .Y(n1086) );
  FADDX1_LVT U1004 ( .A(A[16]), .B(n1091), .CI(n866), .S(DIFF[16]) );
  OA21X1_LVT U1005 ( .A1(n1041), .A2(n1090), .A3(n1087), .Y(n1091) );
  OR2X1_LVT U1006 ( .A1(n867), .A2(A[15]), .Y(n1087) );
  AND2X1_LVT U1007 ( .A1(A[15]), .A2(n867), .Y(n1090) );
  FADDX1_LVT U1008 ( .A(n1041), .B(A[15]), .CI(n867), .S(DIFF[15]) );
  FADDX1_LVT U1009 ( .A(A[14]), .B(B[14]), .CI(n1098), .S(DIFF[14]) );
  AO22X1_LVT U1010 ( .A1(n1099), .A2(n1097), .A3(B[13]), .A4(n899), .Y(n1098)
         );
  OR2X1_LVT U1011 ( .A1(n899), .A2(B[13]), .Y(n1097) );
  FADDX1_LVT U1012 ( .A(A[13]), .B(B[13]), .CI(n1099), .S(DIFF[13]) );
  AND2X1_LVT U1013 ( .A1(n1093), .A2(n1100), .Y(n1099) );
  NAND3X0_LVT U1014 ( .A1(n1101), .A2(n1095), .A3(n1096), .Y(n1100) );
  NAND2X0_LVT U1015 ( .A1(B[12]), .A2(n900), .Y(n1095) );
  AO222X1_LVT U1016 ( .A1(B[12]), .A2(n900), .A3(B[12]), .A4(n1102), .A5(n900), 
        .A6(n1102), .Y(n1093) );
  FADDX1_LVT U1017 ( .A(B[12]), .B(n1103), .CI(n900), .S(DIFF[12]) );
  OA21X1_LVT U1018 ( .A1(n868), .A2(n1101), .A3(n1096), .Y(n1103) );
  OR2X1_LVT U1019 ( .A1(n869), .A2(A[11]), .Y(n1096) );
  NAND2X0_LVT U1020 ( .A1(A[11]), .A2(n869), .Y(n1102) );
  FADDX1_LVT U1021 ( .A(A[11]), .B(n869), .CI(n1101), .S(DIFF[11]) );
  AO21X1_LVT U1022 ( .A1(n1092), .A2(n872), .A3(n1094), .Y(n1101) );
  AO222X1_LVT U1023 ( .A1(A[10]), .A2(n870), .A3(n1104), .A4(n1105), .A5(n1106), .A6(n1107), .Y(n1094) );
  AND2X1_LVT U1024 ( .A1(n1108), .A2(n1105), .Y(n1106) );
  AND4X1_LVT U1025 ( .A1(n1109), .A2(n910), .A3(n1108), .A4(n1105), .Y(n1092)
         );
  OR2X1_LVT U1026 ( .A1(n870), .A2(A[10]), .Y(n1105) );
  FADDX1_LVT U1027 ( .A(A[10]), .B(n1110), .CI(n870), .S(DIFF[10]) );
  OA21X1_LVT U1028 ( .A1(n1104), .A2(n908), .A3(n1108), .Y(n1110) );
  NAND2X0_LVT U1029 ( .A1(B[9]), .A2(n901), .Y(n1108) );
  OA222X1_LVT U1030 ( .A1(n1107), .A2(n1109), .A3(n1107), .A4(n910), .A5(n1107), .A6(n872), .Y(n908) );
  OA221X1_LVT U1031 ( .A1(n1111), .A2(n934), .A3(n1111), .A4(n935), .A5(n1112), 
        .Y(n912) );
  AO222X1_LVT U1032 ( .A1(B[6]), .A2(n903), .A3(B[6]), .A4(n1113), .A5(n903), 
        .A6(n1113), .Y(n1112) );
  NAND2X0_LVT U1033 ( .A1(A[5]), .A2(n873), .Y(n1113) );
  NAND3X0_LVT U1034 ( .A1(n1114), .A2(n977), .A3(n1115), .Y(n935) );
  NAND2X0_LVT U1035 ( .A1(B[3]), .A2(n905), .Y(n1115) );
  NAND2X0_LVT U1036 ( .A1(B[0]), .A2(n833), .Y(n1049) );
  NAND2X0_LVT U1037 ( .A1(B[1]), .A2(n907), .Y(n1050) );
  NAND2X0_LVT U1038 ( .A1(B[4]), .A2(n904), .Y(n1114) );
  AO222X1_LVT U1039 ( .A1(B[4]), .A2(n904), .A3(B[4]), .A4(n976), .A5(n904), 
        .A6(n976), .Y(n934) );
  NAND2X0_LVT U1040 ( .A1(A[3]), .A2(n874), .Y(n976) );
  NAND2X0_LVT U1041 ( .A1(n1116), .A2(n915), .Y(n1111) );
  OR2X1_LVT U1042 ( .A1(n873), .A2(A[5]), .Y(n915) );
  NAND2X0_LVT U1043 ( .A1(B[6]), .A2(n903), .Y(n1116) );
  NAND2X0_LVT U1044 ( .A1(B[7]), .A2(n902), .Y(n910) );
  AO22X1_LVT U1045 ( .A1(A[8]), .A2(n871), .A3(n911), .A4(n1109), .Y(n1107) );
  OR2X1_LVT U1046 ( .A1(n871), .A2(A[8]), .Y(n1109) );
  NOR2X0_LVT U1047 ( .A1(n901), .A2(B[9]), .Y(n1104) );
  AO22X1_LVT U1048 ( .A1(A[0]), .A2(n877), .A3(n833), .A4(B[0]), .Y(DIFF[0])
         );
endmodule


module MulDiv ( clock, reset, io_req_ready, io_req_valid, io_req_bits_fn, 
        io_req_bits_dw, io_req_bits_in1, io_req_bits_in2, io_req_bits_tag, 
        io_kill, io_resp_ready, io_resp_valid, io_resp_bits_data, 
        io_resp_bits_tag_4__BAR, io_resp_bits_tag_2_, io_resp_bits_tag_0_, 
        io_resp_bits_tag_3__BAR, io_resp_bits_tag_1__BAR );
  input [3:0] io_req_bits_fn;
  input [63:0] io_req_bits_in1;
  input [63:0] io_req_bits_in2;
  input [4:0] io_req_bits_tag;
  output [63:0] io_resp_bits_data;
  input clock, reset, io_req_valid, io_req_bits_dw, io_kill, io_resp_ready;
  output io_req_ready, io_resp_valid, io_resp_bits_tag_4__BAR,
         io_resp_bits_tag_2_, io_resp_bits_tag_0_, io_resp_bits_tag_3__BAR,
         io_resp_bits_tag_1__BAR;
  wire   resHi, n_T_59_8_, neg_out, n_T_71_39_, isHi, n_T_97_6_, n_T_273_5_,
         n_T_430_5_, N282, N283, N284, N285, N293, N294, N295, N296, N297,
         N298, N299, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424,
         N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435,
         N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479,
         N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490,
         N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523,
         net34684, net34690, net34695, net34700, net34705, n166, n167, n168,
         n169, n170, n171, n179, n185, n196, n202, n205, n217, n219, n220,
         n228, n229, n231, n232, n233, n234, n236, n237, n238, n239, n240,
         n241, n243, n246, n247, n248, n249, n250, n251, n252, n254, n255,
         n256, n257, n258, n259, n260, n261, n263, n264, n266, n267, n268,
         n269, n270, n272, n273, n274, n275, n277, n278, n281, n282, n283,
         n284, n286, n290, n291, n292, n293, n296, n793, n794, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n80, n81, n82, n83,
         n85, n86, n87, n88, n90, n91, n92, n93, n95, n96, n97, n98, n100,
         n101, n102, n103, n104, n105, n106, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n120, n121, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n135, n136, n137,
         n138, n139, n140, n141, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n172, n173, n174, n175, n176, n177, n178, n180,
         n181, n182, n183, n184, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n197, n198, n199, n200, n201, n203, n204, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n218,
         n221, n222, n223, n224, n225, n226, n227, n230, n235, n242, n244,
         n245, n253, n262, n265, n271, n276, n279, n280, n285, n287, n288,
         n289, n294, n295, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n795, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64;
  wire   [64:0] divisor;
  wire   [64:0] subtractor;
  wire   [63:0] result;
  wire   [63:1] negated_remainder;
  wire   [128:0] n_T_51;
  wire   [72:0] n_T_65;
  wire   [9:4] n_T_69;
  wire   [5:4] n_T_85;
  wire   [63:0] n_T_87;
  wire   [4:0] n_T_272;
  wire   [4:0] n_T_429;
  wire   [5:0] n_T_434;
  wire   [126:0] n_T_442;

  SNPS_CLOCK_GATE_HIGH_MulDiv_0 clk_gate_divisor_reg ( .CLK(clock), .EN(N322), 
        .ENCLK(net34684), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_4 clk_gate_req_dw_reg ( .CLK(clock), .EN(n235), 
        .ENCLK(net34690), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_3 clk_gate_count_reg ( .CLK(clock), .EN(N293), 
        .ENCLK(net34695), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_2 clk_gate_state_reg ( .CLK(clock), .EN(N282), 
        .ENCLK(net34700), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_MulDiv_1 clk_gate_remainder_reg ( .CLK(clock), .EN(N493), .ENCLK(net34705), .TE(1'b0) );
  MulDiv_DP_OP_279J39_124_314_J39_0 DP_OP_279J39_124_314 ( .I1({n301, 
        n_T_51[7], n307, n_T_51[5], n306, n305, n304, n303, n302}), .I2(
        divisor), .I3(n_T_51[128:64]), .O1(n_T_65) );
  MulDiv_DW_leftsh_J39_0 ash_111 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_T_51[63:7], 
        n307, n_T_51[5], n306, n305, n304, n303, n302}), .SH({n170, n169, n168, 
        n167, n166, n171}), .B(n_T_442) );
  MulDiv_DW01_sub_J39_0 sub_x_110 ( .A({n_T_430_5_, n_T_429}), .B({n_T_273_5_, 
        n_T_272}), .CI(1'b0), .DIFF(n_T_434) );
  MulDiv_DW_rightsh_J39_0 ashr_12 ( .A({n_T_51[126:7], n307, n_T_51[5], n306, 
        n305, n304, n303, n302}), .DATA_TC(1'b0), .SH({n_T_85, n300, 1'b0, 
        1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, n_T_87}) );
  MulDiv_DW01_sub_J39_2 sub_x_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(result), 
        .CI(1'b0), .DIFF({negated_remainder, SYNOPSYS_UNCONNECTED_64}) );
  MulDiv_DW01_sub_J39_3 sub_x_7 ( .A({n_T_51[127:64], n301}), .B(divisor), 
        .CI(1'b0), .DIFF(subtractor) );
  DFFX1_LVT remainder_reg_0_ ( .D(N394), .CLK(n288), .Q(n_T_51[0]) );
  DFFX1_LVT remainder_reg_1_ ( .D(N395), .CLK(n288), .Q(n_T_51[1]), .QN(n296)
         );
  DFFX1_LVT remainder_reg_2_ ( .D(N396), .CLK(n288), .QN(n208) );
  DFFX1_LVT remainder_reg_3_ ( .D(N397), .CLK(n288), .Q(n_T_51[3]) );
  DFFX1_LVT remainder_reg_4_ ( .D(N398), .CLK(n288), .Q(n_T_51[4]), .QN(n293)
         );
  DFFX1_LVT remainder_reg_5_ ( .D(N399), .CLK(n288), .Q(n_T_51[5]), .QN(n292)
         );
  DFFX1_LVT remainder_reg_6_ ( .D(N400), .CLK(n288), .Q(n_T_51[6]), .QN(n291)
         );
  DFFX1_LVT remainder_reg_7_ ( .D(N401), .CLK(n288), .Q(n_T_51[7]), .QN(n290)
         );
  DFFX1_LVT remainder_reg_8_ ( .D(N402), .CLK(n288), .Q(n_T_51[8]), .QN(n186)
         );
  DFFX1_LVT remainder_reg_9_ ( .D(N403), .CLK(n288), .Q(n_T_51[9]), .QN(n147)
         );
  DFFX1_LVT remainder_reg_10_ ( .D(N404), .CLK(n287), .Q(n_T_51[10]), .QN(n286) );
  DFFX1_LVT remainder_reg_11_ ( .D(N405), .CLK(n287), .Q(n_T_51[11]), .QN(n153) );
  DFFX1_LVT remainder_reg_12_ ( .D(N406), .CLK(n287), .Q(n_T_51[12]), .QN(n284) );
  DFFX1_LVT remainder_reg_13_ ( .D(N407), .CLK(n287), .Q(n_T_51[13]), .QN(n283) );
  DFFX1_LVT remainder_reg_14_ ( .D(N408), .CLK(n287), .Q(n_T_51[14]), .QN(n282) );
  DFFX1_LVT remainder_reg_15_ ( .D(N409), .CLK(n287), .Q(n_T_51[15]), .QN(n281) );
  DFFX1_LVT remainder_reg_16_ ( .D(N410), .CLK(n287), .Q(n_T_51[16]), .QN(n183) );
  DFFX1_LVT remainder_reg_17_ ( .D(N411), .CLK(n287), .Q(n_T_51[17]), .QN(n278) );
  DFFX1_LVT remainder_reg_18_ ( .D(N412), .CLK(n287), .Q(n_T_51[18]), .QN(n277) );
  DFFX1_LVT remainder_reg_19_ ( .D(N413), .CLK(n287), .Q(n_T_51[19]), .QN(n152) );
  DFFX1_LVT remainder_reg_20_ ( .D(N414), .CLK(n287), .Q(n_T_51[20]), .QN(n275) );
  DFFX1_LVT remainder_reg_21_ ( .D(N415), .CLK(n287), .Q(n_T_51[21]), .QN(n274) );
  DFFX1_LVT remainder_reg_22_ ( .D(N416), .CLK(n285), .Q(n_T_51[22]), .QN(n273) );
  DFFX1_LVT remainder_reg_23_ ( .D(N417), .CLK(n285), .Q(n_T_51[23]), .QN(n272) );
  DFFX1_LVT remainder_reg_24_ ( .D(N418), .CLK(n285), .Q(n_T_51[24]), .QN(n270) );
  DFFX1_LVT remainder_reg_25_ ( .D(N419), .CLK(n285), .Q(n_T_51[25]), .QN(n269) );
  DFFX1_LVT remainder_reg_26_ ( .D(N420), .CLK(n285), .Q(n_T_51[26]), .QN(n268) );
  DFFX1_LVT remainder_reg_27_ ( .D(N421), .CLK(n285), .Q(n_T_51[27]), .QN(n267) );
  DFFX1_LVT remainder_reg_28_ ( .D(N422), .CLK(n285), .Q(n_T_51[28]), .QN(n266) );
  DFFX1_LVT remainder_reg_29_ ( .D(N423), .CLK(n285), .Q(n_T_51[29]), .QN(n181) );
  DFFX1_LVT remainder_reg_30_ ( .D(N424), .CLK(n285), .Q(n_T_51[30]), .QN(n264) );
  DFFX1_LVT remainder_reg_31_ ( .D(N425), .CLK(n285), .Q(n_T_51[31]), .QN(n263) );
  DFFX1_LVT state_reg_0_ ( .D(N283), .CLK(net34700), .Q(n150), .QN(n220) );
  DFFX1_LVT state_reg_1_ ( .D(N284), .CLK(net34700), .Q(n184), .QN(n219) );
  DFFX1_LVT state_reg_2_ ( .D(N285), .CLK(net34700), .Q(n154), .QN(n217) );
  DFFX1_LVT req_dw_reg ( .D(io_req_bits_dw), .CLK(net34690), .Q(n206), .QN(
        n156) );
  DFFX1_LVT req_tag_reg_4_ ( .D(io_req_bits_tag[4]), .CLK(net34690), .QN(
        io_resp_bits_tag_4__BAR) );
  DFFX1_LVT req_tag_reg_3_ ( .D(io_req_bits_tag[3]), .CLK(net34690), .QN(
        io_resp_bits_tag_3__BAR) );
  DFFX1_LVT req_tag_reg_2_ ( .D(io_req_bits_tag[2]), .CLK(net34690), .Q(
        io_resp_bits_tag_2_) );
  DFFX1_LVT req_tag_reg_1_ ( .D(io_req_bits_tag[1]), .CLK(net34690), .QN(
        io_resp_bits_tag_1__BAR) );
  DFFX1_LVT req_tag_reg_0_ ( .D(io_req_bits_tag[0]), .CLK(net34690), .Q(
        io_resp_bits_tag_0_) );
  DFFSSRX1_LVT count_reg_6_ ( .D(n783), .SETB(n200), .RSTB(n_T_97_6_), .CLK(
        net34695), .Q(n_T_69[9]), .QN(n155) );
  DFFX1_LVT count_reg_5_ ( .D(N299), .CLK(net34695), .Q(n_T_69[8]), .QN(n197)
         );
  DFFX1_LVT count_reg_4_ ( .D(N298), .CLK(net34695), .Q(n_T_69[7]) );
  DFFX1_LVT count_reg_3_ ( .D(N297), .CLK(net34695), .Q(n_T_69[6]), .QN(n198)
         );
  DFFX1_LVT count_reg_2_ ( .D(N296), .CLK(net34695), .Q(n_T_71_39_), .QN(n210)
         );
  DFFX1_LVT count_reg_1_ ( .D(N295), .CLK(net34695), .Q(n_T_69[4]), .QN(n148)
         );
  DFFX1_LVT neg_out_reg ( .D(n793), .CLK(net34695), .Q(neg_out), .QN(n212) );
  DFFX1_LVT divisor_reg_64_ ( .D(N387), .CLK(n299), .Q(divisor[64]) );
  DFFX1_LVT divisor_reg_63_ ( .D(N386), .CLK(n299), .Q(divisor[63]), .QN(n175)
         );
  DFFX1_LVT divisor_reg_62_ ( .D(N385), .CLK(n299), .Q(divisor[62]), .QN(n177)
         );
  DFFX1_LVT divisor_reg_61_ ( .D(N384), .CLK(n299), .Q(divisor[61]) );
  DFFX1_LVT divisor_reg_60_ ( .D(N383), .CLK(n299), .Q(divisor[60]) );
  DFFX1_LVT divisor_reg_59_ ( .D(N382), .CLK(n298), .Q(divisor[59]), .QN(n180)
         );
  DFFX1_LVT divisor_reg_58_ ( .D(N381), .CLK(n298), .Q(divisor[58]), .QN(n179)
         );
  DFFX1_LVT divisor_reg_57_ ( .D(N380), .CLK(n298), .Q(divisor[57]) );
  DFFX1_LVT divisor_reg_56_ ( .D(N379), .CLK(n298), .Q(divisor[56]) );
  DFFX1_LVT divisor_reg_55_ ( .D(N378), .CLK(n298), .Q(divisor[55]) );
  DFFX1_LVT divisor_reg_54_ ( .D(N377), .CLK(n298), .Q(divisor[54]), .QN(n195)
         );
  DFFX1_LVT divisor_reg_53_ ( .D(N376), .CLK(n298), .Q(divisor[53]) );
  DFFX1_LVT divisor_reg_52_ ( .D(N375), .CLK(n298), .Q(divisor[52]) );
  DFFX1_LVT divisor_reg_51_ ( .D(N374), .CLK(n298), .Q(divisor[51]) );
  DFFX1_LVT divisor_reg_50_ ( .D(N373), .CLK(n298), .Q(divisor[50]), .QN(n159)
         );
  DFFX1_LVT divisor_reg_49_ ( .D(N372), .CLK(n298), .Q(divisor[49]) );
  DFFX1_LVT divisor_reg_48_ ( .D(N371), .CLK(n298), .Q(divisor[48]) );
  DFFX1_LVT divisor_reg_47_ ( .D(N370), .CLK(n297), .Q(divisor[47]), .QN(n178)
         );
  DFFX1_LVT divisor_reg_46_ ( .D(N369), .CLK(n297), .Q(divisor[46]), .QN(n194)
         );
  DFFX1_LVT divisor_reg_45_ ( .D(N368), .CLK(n297), .Q(divisor[45]), .QN(n173)
         );
  DFFX1_LVT divisor_reg_44_ ( .D(N367), .CLK(n297), .Q(divisor[44]) );
  DFFX1_LVT divisor_reg_43_ ( .D(N366), .CLK(n297), .Q(divisor[43]) );
  DFFX1_LVT divisor_reg_42_ ( .D(N365), .CLK(n297), .Q(divisor[42]), .QN(n185)
         );
  DFFX1_LVT divisor_reg_41_ ( .D(N364), .CLK(n297), .Q(divisor[41]) );
  DFFX1_LVT divisor_reg_40_ ( .D(N363), .CLK(n297), .Q(divisor[40]), .QN(n163)
         );
  DFFX1_LVT divisor_reg_39_ ( .D(N362), .CLK(n297), .Q(divisor[39]) );
  DFFX1_LVT divisor_reg_38_ ( .D(N361), .CLK(n297), .Q(divisor[38]), .QN(n192)
         );
  DFFX1_LVT divisor_reg_37_ ( .D(N360), .CLK(n297), .Q(divisor[37]) );
  DFFX1_LVT divisor_reg_36_ ( .D(N359), .CLK(n297), .Q(divisor[36]) );
  DFFX1_LVT divisor_reg_35_ ( .D(N358), .CLK(n295), .Q(divisor[35]) );
  DFFX1_LVT divisor_reg_34_ ( .D(N357), .CLK(n295), .Q(divisor[34]), .QN(n160)
         );
  DFFX1_LVT divisor_reg_33_ ( .D(N356), .CLK(n295), .Q(divisor[33]) );
  DFFX1_LVT divisor_reg_32_ ( .D(N355), .CLK(n295), .Q(divisor[32]) );
  DFFX1_LVT divisor_reg_31_ ( .D(N354), .CLK(n295), .Q(divisor[31]), .QN(n176)
         );
  DFFX1_LVT divisor_reg_30_ ( .D(N353), .CLK(n295), .Q(divisor[30]), .QN(n174)
         );
  DFFX1_LVT divisor_reg_29_ ( .D(N352), .CLK(n295), .Q(divisor[29]) );
  DFFX1_LVT divisor_reg_28_ ( .D(N351), .CLK(n295), .Q(divisor[28]) );
  DFFX1_LVT divisor_reg_27_ ( .D(N350), .CLK(n295), .Q(divisor[27]) );
  DFFX1_LVT divisor_reg_26_ ( .D(N349), .CLK(n295), .Q(divisor[26]), .QN(n196)
         );
  DFFX1_LVT divisor_reg_25_ ( .D(N348), .CLK(n295), .Q(divisor[25]) );
  DFFX1_LVT divisor_reg_24_ ( .D(N347), .CLK(n295), .Q(divisor[24]), .QN(n164)
         );
  DFFX1_LVT divisor_reg_23_ ( .D(N346), .CLK(n294), .Q(divisor[23]) );
  DFFX1_LVT divisor_reg_22_ ( .D(N345), .CLK(n294), .Q(divisor[22]), .QN(n190)
         );
  DFFX1_LVT divisor_reg_21_ ( .D(N344), .CLK(n294), .Q(divisor[21]) );
  DFFX1_LVT divisor_reg_20_ ( .D(N343), .CLK(n294), .Q(divisor[20]) );
  DFFX1_LVT divisor_reg_19_ ( .D(N342), .CLK(n294), .Q(divisor[19]) );
  DFFX1_LVT divisor_reg_18_ ( .D(N341), .CLK(n294), .Q(divisor[18]), .QN(n161)
         );
  DFFX1_LVT divisor_reg_17_ ( .D(N340), .CLK(n294), .Q(divisor[17]) );
  DFFX1_LVT divisor_reg_16_ ( .D(N339), .CLK(n294), .Q(divisor[16]) );
  DFFX1_LVT divisor_reg_15_ ( .D(N338), .CLK(n294), .Q(divisor[15]), .QN(n162)
         );
  DFFX1_LVT divisor_reg_14_ ( .D(N337), .CLK(n294), .Q(divisor[14]), .QN(n193)
         );
  DFFX1_LVT divisor_reg_13_ ( .D(N336), .CLK(n294), .Q(divisor[13]), .QN(n172)
         );
  DFFX1_LVT divisor_reg_12_ ( .D(N335), .CLK(n294), .Q(divisor[12]) );
  DFFX1_LVT divisor_reg_11_ ( .D(N334), .CLK(n289), .Q(divisor[11]) );
  DFFX1_LVT divisor_reg_10_ ( .D(N333), .CLK(n289), .Q(divisor[10]), .QN(n202)
         );
  DFFX1_LVT divisor_reg_9_ ( .D(N332), .CLK(n289), .Q(divisor[9]) );
  DFFX1_LVT divisor_reg_8_ ( .D(N331), .CLK(n289), .Q(divisor[8]), .QN(n165)
         );
  DFFX1_LVT divisor_reg_7_ ( .D(N330), .CLK(n289), .Q(divisor[7]) );
  DFFX1_LVT divisor_reg_6_ ( .D(N329), .CLK(n289), .Q(divisor[6]), .QN(n191)
         );
  DFFX1_LVT divisor_reg_5_ ( .D(N328), .CLK(n289), .Q(divisor[5]) );
  DFFX1_LVT divisor_reg_4_ ( .D(N327), .CLK(n289), .Q(divisor[4]) );
  DFFX1_LVT divisor_reg_3_ ( .D(N326), .CLK(n289), .Q(divisor[3]) );
  DFFX1_LVT divisor_reg_2_ ( .D(N325), .CLK(n289), .Q(divisor[2]), .QN(n205)
         );
  DFFX1_LVT divisor_reg_1_ ( .D(N324), .CLK(n289), .Q(divisor[1]) );
  DFFX1_LVT divisor_reg_0_ ( .D(N323), .CLK(n289), .Q(divisor[0]) );
  DFFX1_LVT remainder_reg_32_ ( .D(N426), .CLK(n285), .Q(n_T_51[32]), .QN(n261) );
  DFFX1_LVT remainder_reg_33_ ( .D(N427), .CLK(n285), .Q(n_T_51[33]), .QN(n260) );
  DFFX1_LVT remainder_reg_34_ ( .D(N428), .CLK(n280), .Q(n_T_51[34]), .QN(n259) );
  DFFX1_LVT remainder_reg_35_ ( .D(N429), .CLK(n280), .Q(n_T_51[35]), .QN(n258) );
  DFFX1_LVT remainder_reg_36_ ( .D(N430), .CLK(n280), .Q(n_T_51[36]), .QN(n257) );
  DFFX1_LVT remainder_reg_37_ ( .D(N431), .CLK(n280), .Q(n_T_51[37]), .QN(n256) );
  DFFX1_LVT remainder_reg_38_ ( .D(N432), .CLK(n280), .Q(n_T_51[38]), .QN(n255) );
  DFFX1_LVT remainder_reg_39_ ( .D(N433), .CLK(n280), .Q(n_T_51[39]), .QN(n254) );
  DFFX1_LVT remainder_reg_40_ ( .D(N434), .CLK(n280), .Q(n_T_51[40]), .QN(n188) );
  DFFX1_LVT remainder_reg_41_ ( .D(N435), .CLK(n280), .Q(n_T_51[41]), .QN(n252) );
  DFFX1_LVT remainder_reg_42_ ( .D(N436), .CLK(n280), .Q(n_T_51[42]), .QN(n251) );
  DFFX1_LVT remainder_reg_43_ ( .D(N437), .CLK(n280), .Q(n_T_51[43]), .QN(n250) );
  DFFX1_LVT remainder_reg_44_ ( .D(N438), .CLK(n280), .Q(n_T_51[44]), .QN(n249) );
  DFFX1_LVT remainder_reg_45_ ( .D(N439), .CLK(n280), .Q(n_T_51[45]), .QN(n248) );
  DFFX1_LVT remainder_reg_46_ ( .D(N440), .CLK(n279), .Q(n_T_51[46]), .QN(n247) );
  DFFX1_LVT remainder_reg_47_ ( .D(N441), .CLK(n279), .Q(n_T_51[47]), .QN(n246) );
  DFFX1_LVT remainder_reg_48_ ( .D(N442), .CLK(n279), .Q(n_T_51[48]), .QN(n243) );
  DFFX1_LVT remainder_reg_49_ ( .D(N443), .CLK(n279), .Q(n_T_51[49]), .QN(n182) );
  DFFX1_LVT remainder_reg_50_ ( .D(N444), .CLK(n279), .Q(n_T_51[50]), .QN(n241) );
  DFFX1_LVT remainder_reg_51_ ( .D(N445), .CLK(n279), .Q(n_T_51[51]), .QN(n240) );
  DFFX1_LVT remainder_reg_52_ ( .D(N446), .CLK(n279), .Q(n_T_51[52]), .QN(n239) );
  DFFX1_LVT remainder_reg_53_ ( .D(N447), .CLK(n279), .Q(n_T_51[53]), .QN(n238) );
  DFFX1_LVT remainder_reg_54_ ( .D(N448), .CLK(n279), .Q(n_T_51[54]), .QN(n237) );
  DFFX1_LVT remainder_reg_55_ ( .D(N449), .CLK(n279), .Q(n_T_51[55]), .QN(n236) );
  DFFX1_LVT remainder_reg_56_ ( .D(N450), .CLK(n279), .Q(n_T_51[56]), .QN(n234) );
  DFFX1_LVT remainder_reg_57_ ( .D(N451), .CLK(n279), .Q(n_T_51[57]), .QN(n233) );
  DFFX1_LVT remainder_reg_58_ ( .D(N452), .CLK(n276), .Q(n_T_51[58]), .QN(n232) );
  DFFX1_LVT remainder_reg_59_ ( .D(N453), .CLK(n276), .Q(n_T_51[59]), .QN(n231) );
  DFFX1_LVT remainder_reg_60_ ( .D(N454), .CLK(n276), .Q(n_T_51[60]), .QN(n187) );
  DFFX1_LVT remainder_reg_61_ ( .D(N455), .CLK(n276), .Q(n_T_51[61]), .QN(n229) );
  DFFX1_LVT remainder_reg_62_ ( .D(N456), .CLK(n276), .Q(n_T_51[62]), .QN(n228) );
  DFFX1_LVT remainder_reg_63_ ( .D(N457), .CLK(n276), .Q(n_T_51[63]), .QN(n149) );
  DFFX1_LVT remainder_reg_64_ ( .D(N458), .CLK(n276), .Q(n_T_59_8_) );
  DFFX1_LVT remainder_reg_65_ ( .D(N459), .CLK(n276), .Q(n_T_51[64]) );
  DFFX1_LVT remainder_reg_66_ ( .D(N460), .CLK(n276), .Q(n_T_51[65]) );
  DFFX1_LVT remainder_reg_67_ ( .D(N461), .CLK(n276), .Q(n_T_51[66]) );
  DFFX1_LVT remainder_reg_68_ ( .D(N462), .CLK(n276), .Q(n_T_51[67]) );
  DFFX1_LVT remainder_reg_69_ ( .D(N463), .CLK(n276), .Q(n_T_51[68]) );
  DFFX1_LVT remainder_reg_70_ ( .D(N464), .CLK(n271), .Q(n_T_51[69]) );
  DFFX1_LVT remainder_reg_71_ ( .D(N465), .CLK(n271), .Q(n_T_51[70]) );
  DFFX1_LVT remainder_reg_72_ ( .D(N466), .CLK(n271), .Q(n_T_51[71]) );
  DFFX1_LVT remainder_reg_73_ ( .D(N467), .CLK(n271), .Q(n_T_51[72]) );
  DFFX1_LVT remainder_reg_74_ ( .D(N468), .CLK(n271), .Q(n_T_51[73]) );
  DFFX1_LVT remainder_reg_75_ ( .D(N469), .CLK(n271), .Q(n_T_51[74]) );
  DFFX1_LVT remainder_reg_76_ ( .D(N470), .CLK(n271), .Q(n_T_51[75]) );
  DFFX1_LVT remainder_reg_77_ ( .D(N471), .CLK(n271), .Q(n_T_51[76]) );
  DFFX1_LVT remainder_reg_78_ ( .D(N472), .CLK(n271), .Q(n_T_51[77]) );
  DFFX1_LVT remainder_reg_79_ ( .D(N473), .CLK(n271), .Q(n_T_51[78]) );
  DFFX1_LVT remainder_reg_80_ ( .D(N474), .CLK(n271), .Q(n_T_51[79]) );
  DFFX1_LVT remainder_reg_81_ ( .D(N475), .CLK(n271), .Q(n_T_51[80]) );
  DFFX1_LVT remainder_reg_82_ ( .D(N476), .CLK(n265), .Q(n_T_51[81]) );
  DFFX1_LVT remainder_reg_83_ ( .D(N477), .CLK(n265), .Q(n_T_51[82]) );
  DFFX1_LVT remainder_reg_84_ ( .D(N478), .CLK(n265), .Q(n_T_51[83]) );
  DFFX1_LVT remainder_reg_85_ ( .D(N479), .CLK(n265), .Q(n_T_51[84]) );
  DFFX1_LVT remainder_reg_86_ ( .D(N480), .CLK(n265), .Q(n_T_51[85]) );
  DFFX1_LVT remainder_reg_87_ ( .D(N481), .CLK(n265), .Q(n_T_51[86]) );
  DFFX1_LVT remainder_reg_88_ ( .D(N482), .CLK(n265), .Q(n_T_51[87]) );
  DFFX1_LVT remainder_reg_89_ ( .D(N483), .CLK(n265), .Q(n_T_51[88]) );
  DFFX1_LVT remainder_reg_90_ ( .D(N484), .CLK(n265), .Q(n_T_51[89]) );
  DFFX1_LVT remainder_reg_91_ ( .D(N485), .CLK(n265), .Q(n_T_51[90]) );
  DFFX1_LVT remainder_reg_92_ ( .D(N486), .CLK(n265), .Q(n_T_51[91]) );
  DFFX1_LVT remainder_reg_93_ ( .D(N487), .CLK(n265), .Q(n_T_51[92]) );
  DFFX1_LVT remainder_reg_94_ ( .D(N488), .CLK(n262), .Q(n_T_51[93]) );
  DFFX1_LVT remainder_reg_95_ ( .D(N489), .CLK(n262), .Q(n_T_51[94]) );
  DFFX1_LVT remainder_reg_96_ ( .D(N490), .CLK(n262), .Q(n_T_51[95]) );
  DFFX1_LVT remainder_reg_97_ ( .D(N491), .CLK(n262), .Q(n_T_51[96]) );
  DFFX1_LVT remainder_reg_98_ ( .D(N492), .CLK(n262), .Q(n_T_51[97]) );
  DFFX1_LVT remainder_reg_99_ ( .D(N494), .CLK(n262), .Q(n_T_51[98]) );
  DFFX1_LVT remainder_reg_100_ ( .D(N495), .CLK(n262), .Q(n_T_51[99]) );
  DFFX1_LVT remainder_reg_101_ ( .D(N496), .CLK(n262), .Q(n_T_51[100]) );
  DFFX1_LVT remainder_reg_102_ ( .D(N497), .CLK(n262), .Q(n_T_51[101]) );
  DFFX1_LVT remainder_reg_103_ ( .D(N498), .CLK(n262), .Q(n_T_51[102]) );
  DFFX1_LVT remainder_reg_104_ ( .D(N499), .CLK(n262), .Q(n_T_51[103]) );
  DFFX1_LVT remainder_reg_105_ ( .D(N500), .CLK(n262), .Q(n_T_51[104]) );
  DFFX1_LVT remainder_reg_106_ ( .D(N501), .CLK(n253), .Q(n_T_51[105]) );
  DFFX1_LVT remainder_reg_107_ ( .D(N502), .CLK(n253), .Q(n_T_51[106]) );
  DFFX1_LVT remainder_reg_108_ ( .D(N503), .CLK(n253), .Q(n_T_51[107]) );
  DFFX1_LVT remainder_reg_109_ ( .D(N504), .CLK(n253), .Q(n_T_51[108]) );
  DFFX1_LVT remainder_reg_110_ ( .D(N505), .CLK(n253), .Q(n_T_51[109]) );
  DFFX1_LVT remainder_reg_111_ ( .D(N506), .CLK(n253), .Q(n_T_51[110]) );
  DFFX1_LVT remainder_reg_112_ ( .D(N507), .CLK(n253), .Q(n_T_51[111]) );
  DFFX1_LVT remainder_reg_113_ ( .D(N508), .CLK(n253), .Q(n_T_51[112]) );
  DFFX1_LVT remainder_reg_114_ ( .D(N509), .CLK(n253), .Q(n_T_51[113]) );
  DFFX1_LVT remainder_reg_115_ ( .D(N510), .CLK(n253), .Q(n_T_51[114]) );
  DFFX1_LVT remainder_reg_116_ ( .D(N511), .CLK(n253), .Q(n_T_51[115]) );
  DFFX1_LVT remainder_reg_117_ ( .D(N512), .CLK(n253), .Q(n_T_51[116]) );
  DFFX1_LVT remainder_reg_118_ ( .D(N513), .CLK(n245), .Q(n_T_51[117]) );
  DFFX1_LVT remainder_reg_119_ ( .D(N514), .CLK(n245), .Q(n_T_51[118]) );
  DFFX1_LVT remainder_reg_120_ ( .D(N515), .CLK(n245), .Q(n_T_51[119]) );
  DFFX1_LVT remainder_reg_121_ ( .D(N516), .CLK(n245), .Q(n_T_51[120]) );
  DFFX1_LVT remainder_reg_122_ ( .D(N517), .CLK(n245), .Q(n_T_51[121]) );
  DFFX1_LVT remainder_reg_123_ ( .D(N518), .CLK(n245), .Q(n_T_51[122]) );
  DFFX1_LVT remainder_reg_124_ ( .D(N519), .CLK(n245), .Q(n_T_51[123]) );
  DFFX1_LVT remainder_reg_125_ ( .D(N520), .CLK(n245), .Q(n_T_51[124]) );
  DFFX1_LVT remainder_reg_126_ ( .D(N521), .CLK(n245), .Q(n_T_51[125]) );
  DFFX1_LVT remainder_reg_127_ ( .D(N522), .CLK(n245), .Q(n_T_51[126]) );
  DFFX1_LVT remainder_reg_128_ ( .D(N523), .CLK(n245), .Q(n_T_51[127]) );
  DFFSSRX1_LVT remainder_reg_129_ ( .D(n230), .SETB(n_T_65[72]), .RSTB(1'b1), 
        .CLK(n245), .QN(n_T_51[128]) );
  DFFX1_LVT resHi_reg ( .D(n794), .CLK(net34700), .Q(resHi) );
  DFFX1_LVT count_reg_0_ ( .D(N294), .CLK(net34695), .Q(n300), .QN(n204) );
  OA21X1_LVT isHi_reg_U2 ( .A1(io_req_bits_fn[2]), .A2(n786), .A3(n785), .Y(
        n145) );
  DFFX1_LVT isHi_reg ( .D(n145), .CLK(net34690), .Q(n189), .QN(isHi) );
  AO221X1_LVT U3 ( .A1(1'b1), .A2(n132), .A3(n_T_87[52]), .A4(n679), .A5(n133), 
        .Y(n135) );
  AO221X1_LVT U4 ( .A1(1'b1), .A2(n135), .A3(n_T_51[51]), .A4(n227), .A5(n136), 
        .Y(N446) );
  AO221X1_LVT U5 ( .A1(1'b1), .A2(n120), .A3(n_T_87[32]), .A4(n679), .A5(n121), 
        .Y(n123) );
  AO221X1_LVT U6 ( .A1(1'b1), .A2(n123), .A3(n_T_51[31]), .A4(n227), .A5(n124), 
        .Y(N426) );
  AO221X1_LVT U7 ( .A1(1'b1), .A2(n117), .A3(n225), .A4(n_T_442[1]), .A5(n118), 
        .Y(N395) );
  AO221X1_LVT U8 ( .A1(1'b1), .A2(n105), .A3(n225), .A4(n_T_442[4]), .A5(n106), 
        .Y(N398) );
  AO221X1_LVT U9 ( .A1(1'b1), .A2(n97), .A3(n227), .A4(n_T_51[15]), .A5(n98), 
        .Y(n100) );
  AO221X1_LVT U10 ( .A1(1'b1), .A2(n92), .A3(n225), .A4(n_T_442[2]), .A5(n93), 
        .Y(N396) );
  AO221X1_LVT U11 ( .A1(1'b1), .A2(n87), .A3(n157), .A4(n_T_442[24]), .A5(n88), 
        .Y(N418) );
  AO221X1_LVT U12 ( .A1(1'b1), .A2(n977), .A3(n_T_51[63]), .A4(n224), .A5(N293), .Y(N493) );
  AO221X1_LVT U13 ( .A1(1'b1), .A2(n77), .A3(n_T_87[40]), .A4(n679), .A5(n78), 
        .Y(n80) );
  AO221X1_LVT U14 ( .A1(1'b1), .A2(n80), .A3(n_T_51[39]), .A4(n227), .A5(n81), 
        .Y(N434) );
  AO221X1_LVT U15 ( .A1(1'b1), .A2(n72), .A3(n225), .A4(n_T_442[12]), .A5(n73), 
        .Y(N406) );
  AO221X1_LVT U16 ( .A1(1'b1), .A2(n65), .A3(n_T_87[48]), .A4(n679), .A5(n66), 
        .Y(n68) );
  AO221X1_LVT U17 ( .A1(1'b1), .A2(n68), .A3(n_T_51[47]), .A4(n227), .A5(n69), 
        .Y(N442) );
  AO221X1_LVT U18 ( .A1(1'b1), .A2(n971), .A3(n999), .A4(n795), .A5(n970), .Y(
        n58) );
  AO221X1_LVT U19 ( .A1(1'b1), .A2(n44), .A3(n_T_87[56]), .A4(n679), .A5(n45), 
        .Y(n47) );
  AO221X1_LVT U20 ( .A1(1'b1), .A2(n47), .A3(n224), .A4(negated_remainder[56]), 
        .A5(n48), .Y(N450) );
  AO222X1_LVT U21 ( .A1(n753), .A2(n224), .A3(n680), .A4(1'b1), .A5(n29), .A6(
        n235), .Y(N283) );
  AO221X1_LVT U22 ( .A1(1'b1), .A2(n12), .A3(n1003), .A4(n15), .A5(n22), .Y(
        n_T_429[1]) );
  OA221X1_LVT U23 ( .A1(n975), .A2(n30), .A3(n777), .A4(n997), .A5(n776), .Y(
        n31) );
  INVX1_LVT U24 ( .A(n209), .Y(n146) );
  AOI222X1_LVT U25 ( .A1(n_T_51[23]), .A2(n775), .A3(n749), .A4(n_T_51[19]), 
        .A5(n_T_51[27]), .A6(n776), .Y(n2) );
  AND2X1_LVT U26 ( .A1(n263), .A2(n2), .Y(n755) );
  NAND2X0_LVT U27 ( .A1(subtractor[46]), .A2(n754), .Y(n3) );
  NAND2X0_LVT U28 ( .A1(n655), .A2(io_req_bits_in2[46]), .Y(n4) );
  NAND3X0_LVT U29 ( .A1(n3), .A2(n633), .A3(n4), .Y(N369) );
  NAND2X0_LVT U30 ( .A1(subtractor[40]), .A2(n754), .Y(n5) );
  NAND2X0_LVT U31 ( .A1(n655), .A2(io_req_bits_in2[40]), .Y(n6) );
  NAND3X0_LVT U32 ( .A1(n5), .A2(n633), .A3(n6), .Y(N363) );
  NAND2X0_LVT U33 ( .A1(subtractor[50]), .A2(n754), .Y(n7) );
  NAND2X0_LVT U34 ( .A1(n655), .A2(io_req_bits_in2[50]), .Y(n8) );
  NAND3X0_LVT U35 ( .A1(n7), .A2(n633), .A3(n8), .Y(N373) );
  OA21X1_LVT U36 ( .A1(n232), .A2(n746), .A3(n228), .Y(n9) );
  NAND2X0_LVT U37 ( .A1(n773), .A2(n_T_51[54]), .Y(n10) );
  NAND2X0_LVT U38 ( .A1(n747), .A2(n_T_51[50]), .Y(n11) );
  NAND4X0_LVT U39 ( .A1(n9), .A2(n758), .A3(n10), .A4(n11), .Y(n12) );
  AOI22X1_LVT U40 ( .A1(n775), .A2(n_T_51[22]), .A3(n_T_51[18]), .A4(n749), 
        .Y(n13) );
  OR2X1_LVT U41 ( .A1(n268), .A2(n748), .Y(n14) );
  NAND4X0_LVT U42 ( .A1(n264), .A2(n755), .A3(n13), .A4(n14), .Y(n15) );
  AOI22X1_LVT U43 ( .A1(n_T_51[34]), .A2(n742), .A3(n_T_51[38]), .A4(n741), 
        .Y(n16) );
  OR2X1_LVT U44 ( .A1(n251), .A2(n740), .Y(n17) );
  NAND4X0_LVT U45 ( .A1(n247), .A2(n756), .A3(n16), .A4(n17), .Y(n18) );
  AOI22X1_LVT U46 ( .A1(n304), .A2(n745), .A3(n_T_51[6]), .A4(n744), .Y(n19)
         );
  OR2X1_LVT U47 ( .A1(n286), .A2(n743), .Y(n20) );
  NAND4X0_LVT U48 ( .A1(n282), .A2(n757), .A3(n19), .A4(n20), .Y(n21) );
  AO22X1_LVT U49 ( .A1(n1002), .A2(n18), .A3(n1001), .A4(n21), .Y(n22) );
  NAND2X0_LVT U51 ( .A1(subtractor[47]), .A2(n754), .Y(n24) );
  NAND2X0_LVT U52 ( .A1(n655), .A2(io_req_bits_in2[47]), .Y(n25) );
  NAND3X0_LVT U53 ( .A1(n24), .A2(n633), .A3(n25), .Y(N370) );
  AOI222X1_LVT U54 ( .A1(n_T_51[51]), .A2(n747), .A3(n_T_51[55]), .A4(n773), 
        .A5(n_T_51[59]), .A6(n774), .Y(n26) );
  AND2X1_LVT U55 ( .A1(n149), .A2(n26), .Y(n758) );
  NAND2X0_LVT U56 ( .A1(subtractor[54]), .A2(n754), .Y(n27) );
  NAND2X0_LVT U57 ( .A1(n655), .A2(io_req_bits_in2[54]), .Y(n28) );
  NAND3X0_LVT U58 ( .A1(n27), .A2(n633), .A3(n28), .Y(N377) );
  AND2X1_LVT U59 ( .A1(n309), .A2(io_req_bits_fn[2]), .Y(n29) );
  OA21X1_LVT U60 ( .A1(n1000), .A2(n781), .A3(n780), .Y(n30) );
  INVX0_LVT U61 ( .A(n773), .Y(n32) );
  OA22X1_LVT U62 ( .A1(n_T_430_5_), .A2(n31), .A3(n779), .A4(n32), .Y(n33) );
  NAND2X0_LVT U63 ( .A1(n971), .A2(n772), .Y(n34) );
  AO21X1_LVT U64 ( .A1(n771), .A2(n34), .A3(n972), .Y(n35) );
  NAND3X0_LVT U65 ( .A1(n774), .A2(n33), .A3(n35), .Y(n_T_429[2]) );
  NAND2X0_LVT U66 ( .A1(subtractor[53]), .A2(n754), .Y(n36) );
  NAND2X0_LVT U67 ( .A1(n655), .A2(io_req_bits_in2[53]), .Y(n37) );
  NAND3X0_LVT U68 ( .A1(n36), .A2(n633), .A3(n37), .Y(N376) );
  NAND2X0_LVT U69 ( .A1(subtractor[41]), .A2(n754), .Y(n38) );
  NAND2X0_LVT U70 ( .A1(n655), .A2(io_req_bits_in2[41]), .Y(n39) );
  NAND3X0_LVT U71 ( .A1(n38), .A2(n633), .A3(n39), .Y(N364) );
  NAND2X0_LVT U72 ( .A1(subtractor[55]), .A2(n754), .Y(n40) );
  NAND2X0_LVT U73 ( .A1(n655), .A2(io_req_bits_in2[55]), .Y(n41) );
  NAND3X0_LVT U74 ( .A1(n40), .A2(n633), .A3(n41), .Y(N378) );
  AOI222X1_LVT U76 ( .A1(n_T_51[39]), .A2(n741), .A3(n_T_51[35]), .A4(n742), 
        .A5(n_T_51[43]), .A6(n771), .Y(n43) );
  AND2X1_LVT U77 ( .A1(n246), .A2(n43), .Y(n756) );
  INVX0_LVT U78 ( .A(n658), .Y(n44) );
  AO22X1_LVT U79 ( .A1(n_T_65[0]), .A2(n223), .A3(io_req_bits_in1[56]), .A4(
        n655), .Y(n45) );
  AO22X1_LVT U81 ( .A1(n_T_51[55]), .A2(n227), .A3(n225), .A4(n_T_442[56]), 
        .Y(n48) );
  NAND2X0_LVT U82 ( .A1(subtractor[58]), .A2(n754), .Y(n49) );
  NAND2X0_LVT U83 ( .A1(n655), .A2(io_req_bits_in2[58]), .Y(n50) );
  NAND3X0_LVT U84 ( .A1(n49), .A2(n633), .A3(n50), .Y(N381) );
  OA22X1_LVT U85 ( .A1(n773), .A2(n789), .A3(n775), .A4(n788), .Y(n51) );
  OA22X1_LVT U86 ( .A1(n148), .A2(n210), .A3(n973), .A4(n974), .Y(n52) );
  NOR4X0_LVT U87 ( .A1(n302), .A2(n305), .A3(n304), .A4(n52), .Y(n53) );
  AND4X1_LVT U88 ( .A1(n781), .A2(n189), .A3(n296), .A4(n53), .Y(n54) );
  NAND2X0_LVT U89 ( .A1(n732), .A2(n779), .Y(n55) );
  NAND3X0_LVT U90 ( .A1(n55), .A2(n148), .A3(n210), .Y(n56) );
  NAND2X0_LVT U92 ( .A1(n210), .A2(n58), .Y(n59) );
  AND4X1_LVT U93 ( .A1(n51), .A2(n54), .A3(n56), .A4(n59), .Y(n60) );
  NAND2X0_LVT U94 ( .A1(n1000), .A2(n800), .Y(n61) );
  NAND4X0_LVT U95 ( .A1(n790), .A2(n980), .A3(n60), .A4(n61), .Y(n338) );
  NAND2X0_LVT U96 ( .A1(subtractor[49]), .A2(n754), .Y(n62) );
  NAND2X0_LVT U97 ( .A1(n655), .A2(io_req_bits_in2[49]), .Y(n63) );
  NAND3X0_LVT U98 ( .A1(n62), .A2(n633), .A3(n63), .Y(N372) );
  INVX0_LVT U99 ( .A(subtractor[64]), .Y(n64) );
  NAND2X0_LVT U100 ( .A1(n343), .A2(n64), .Y(n207) );
  AO22X1_LVT U101 ( .A1(n209), .A2(result[22]), .A3(result[54]), .A4(n146), 
        .Y(io_resp_bits_data[22]) );
  INVX0_LVT U102 ( .A(n658), .Y(n65) );
  AO22X1_LVT U103 ( .A1(n_T_51[56]), .A2(n223), .A3(io_req_bits_in1[48]), .A4(
        n655), .Y(n66) );
  AO22X1_LVT U105 ( .A1(n224), .A2(negated_remainder[48]), .A3(n225), .A4(
        n_T_442[48]), .Y(n69) );
  NAND2X0_LVT U106 ( .A1(subtractor[57]), .A2(n754), .Y(n70) );
  NAND2X0_LVT U107 ( .A1(n655), .A2(io_req_bits_in2[57]), .Y(n71) );
  NAND3X0_LVT U108 ( .A1(n70), .A2(n633), .A3(n71), .Y(N380) );
  AO222X1_LVT U109 ( .A1(n_T_51[20]), .A2(n223), .A3(n679), .A4(n_T_87[12]), 
        .A5(io_req_bits_in1[12]), .A6(n235), .Y(n72) );
  AO22X1_LVT U110 ( .A1(n224), .A2(negated_remainder[12]), .A3(n_T_51[11]), 
        .A4(n227), .Y(n73) );
  AND4X1_LVT U112 ( .A1(n_T_69[4]), .A2(n613), .A3(n_T_71_39_), .A4(n614), .Y(
        n75) );
  AND3X1_LVT U113 ( .A1(n204), .A2(neg_out), .A3(n75), .Y(n76) );
  AO222X1_LVT U114 ( .A1(n783), .A2(n76), .A3(n157), .A4(n_T_442[64]), .A5(
        n227), .A6(n_T_51[63]), .Y(N458) );
  INVX0_LVT U115 ( .A(n658), .Y(n77) );
  AO22X1_LVT U116 ( .A1(n_T_51[48]), .A2(n223), .A3(io_req_bits_in1[40]), .A4(
        n655), .Y(n78) );
  AO22X1_LVT U118 ( .A1(n224), .A2(negated_remainder[40]), .A3(n225), .A4(
        n_T_442[40]), .Y(n81) );
  NAND2X0_LVT U119 ( .A1(subtractor[63]), .A2(n754), .Y(n82) );
  NAND2X0_LVT U120 ( .A1(n655), .A2(io_req_bits_in2[63]), .Y(n83) );
  NAND3X0_LVT U121 ( .A1(n82), .A2(n633), .A3(n83), .Y(N386) );
  NAND2X0_LVT U123 ( .A1(subtractor[60]), .A2(n754), .Y(n85) );
  NAND2X0_LVT U124 ( .A1(n655), .A2(io_req_bits_in2[60]), .Y(n86) );
  NAND3X0_LVT U125 ( .A1(n85), .A2(n633), .A3(n86), .Y(N383) );
  AO222X1_LVT U126 ( .A1(n_T_51[32]), .A2(n223), .A3(n679), .A4(n_T_87[24]), 
        .A5(io_req_bits_in1[24]), .A6(n235), .Y(n87) );
  AO22X1_LVT U127 ( .A1(n224), .A2(negated_remainder[24]), .A3(n_T_51[23]), 
        .A4(n227), .Y(n88) );
  INVX0_LVT U129 ( .A(n286), .Y(n90) );
  INVX0_LVT U130 ( .A(n201), .Y(n91) );
  AO222X1_LVT U131 ( .A1(n90), .A2(n91), .A3(negated_remainder[2]), .A4(n224), 
        .A5(n235), .A6(io_req_bits_in1[2]), .Y(n92) );
  AO22X1_LVT U132 ( .A1(n679), .A2(n_T_87[2]), .A3(n_T_51[1]), .A4(n227), .Y(
        n93) );
  NAND2X0_LVT U134 ( .A1(subtractor[61]), .A2(n754), .Y(n95) );
  NAND2X0_LVT U135 ( .A1(n655), .A2(io_req_bits_in2[61]), .Y(n96) );
  NAND3X0_LVT U136 ( .A1(n95), .A2(n633), .A3(n96), .Y(N384) );
  AO22X1_LVT U137 ( .A1(n_T_51[24]), .A2(n223), .A3(io_req_bits_in1[16]), .A4(
        n235), .Y(n97) );
  AO22X1_LVT U138 ( .A1(n679), .A2(n_T_87[16]), .A3(n224), .A4(
        negated_remainder[16]), .Y(n98) );
  AO21X1_LVT U140 ( .A1(n_T_442[16]), .A2(n225), .A3(n100), .Y(N410) );
  AO22X1_LVT U141 ( .A1(n209), .A2(result[11]), .A3(result[43]), .A4(n146), 
        .Y(io_resp_bits_data[11]) );
  NAND2X0_LVT U142 ( .A1(subtractor[43]), .A2(n754), .Y(n101) );
  NAND2X0_LVT U143 ( .A1(n655), .A2(io_req_bits_in2[43]), .Y(n102) );
  NAND3X0_LVT U144 ( .A1(n101), .A2(n633), .A3(n102), .Y(N366) );
  NAND2X0_LVT U145 ( .A1(n655), .A2(io_req_bits_in2[62]), .Y(n103) );
  NAND2X0_LVT U146 ( .A1(subtractor[62]), .A2(n754), .Y(n104) );
  NAND3X0_LVT U147 ( .A1(n104), .A2(n633), .A3(n103), .Y(N385) );
  AO222X1_LVT U148 ( .A1(n_T_51[12]), .A2(n223), .A3(n224), .A4(
        negated_remainder[4]), .A5(io_req_bits_in1[4]), .A6(n235), .Y(n105) );
  AO22X1_LVT U149 ( .A1(n679), .A2(n_T_87[4]), .A3(n305), .A4(n227), .Y(n106)
         );
  AOI222X1_LVT U151 ( .A1(n_T_51[8]), .A2(n223), .A3(n224), .A4(result[0]), 
        .A5(io_req_bits_in1[0]), .A6(n235), .Y(n108) );
  AOI22X1_LVT U152 ( .A1(n_T_87[0]), .A2(n679), .A3(n157), .A4(n_T_442[0]), 
        .Y(n109) );
  NAND3X0_LVT U153 ( .A1(n108), .A2(n207), .A3(n109), .Y(N394) );
  INVX0_LVT U154 ( .A(n344), .Y(n110) );
  AND3X1_LVT U155 ( .A1(n342), .A2(n343), .A3(n110), .Y(n157) );
  NAND2X0_LVT U156 ( .A1(subtractor[32]), .A2(n754), .Y(n111) );
  NAND2X0_LVT U157 ( .A1(n655), .A2(io_req_bits_in2[32]), .Y(n112) );
  NAND3X0_LVT U158 ( .A1(n111), .A2(n633), .A3(n112), .Y(N355) );
  NAND2X0_LVT U159 ( .A1(subtractor[44]), .A2(n754), .Y(n113) );
  NAND2X0_LVT U160 ( .A1(n655), .A2(io_req_bits_in2[44]), .Y(n114) );
  NAND3X0_LVT U161 ( .A1(n113), .A2(n633), .A3(n114), .Y(N367) );
  NAND2X0_LVT U162 ( .A1(subtractor[51]), .A2(n754), .Y(n115) );
  NAND2X0_LVT U163 ( .A1(n655), .A2(io_req_bits_in2[51]), .Y(n116) );
  NAND3X0_LVT U164 ( .A1(n115), .A2(n633), .A3(n116), .Y(N374) );
  AO222X1_LVT U165 ( .A1(n223), .A2(n_T_51[9]), .A3(n235), .A4(
        io_req_bits_in1[1]), .A5(negated_remainder[1]), .A6(n224), .Y(n117) );
  AO22X1_LVT U166 ( .A1(n679), .A2(n_T_87[1]), .A3(n302), .A4(n227), .Y(n118)
         );
  INVX0_LVT U168 ( .A(n658), .Y(n120) );
  AO22X1_LVT U169 ( .A1(n_T_51[40]), .A2(n223), .A3(io_req_bits_in1[32]), .A4(
        n655), .Y(n121) );
  AO22X1_LVT U171 ( .A1(n224), .A2(negated_remainder[32]), .A3(n225), .A4(
        n_T_442[32]), .Y(n124) );
  NAND2X0_LVT U172 ( .A1(subtractor[35]), .A2(n754), .Y(n125) );
  NAND2X0_LVT U173 ( .A1(n655), .A2(io_req_bits_in2[35]), .Y(n126) );
  NAND3X0_LVT U174 ( .A1(n125), .A2(n633), .A3(n126), .Y(N358) );
  NAND2X0_LVT U175 ( .A1(subtractor[52]), .A2(n754), .Y(n127) );
  NAND2X0_LVT U176 ( .A1(n655), .A2(io_req_bits_in2[52]), .Y(n128) );
  NAND3X0_LVT U177 ( .A1(n127), .A2(n633), .A3(n128), .Y(N375) );
  NAND2X0_LVT U178 ( .A1(subtractor[56]), .A2(n754), .Y(n129) );
  NAND2X0_LVT U179 ( .A1(n655), .A2(io_req_bits_in2[56]), .Y(n130) );
  NAND3X0_LVT U180 ( .A1(n129), .A2(n633), .A3(n130), .Y(N379) );
  INVX0_LVT U181 ( .A(n1000), .Y(n131) );
  AND2X1_LVT U182 ( .A1(n781), .A2(n131), .Y(n745) );
  INVX0_LVT U183 ( .A(n658), .Y(n132) );
  AO22X1_LVT U184 ( .A1(n_T_51[60]), .A2(n223), .A3(io_req_bits_in1[52]), .A4(
        n655), .Y(n133) );
  AO22X1_LVT U186 ( .A1(n224), .A2(negated_remainder[52]), .A3(n225), .A4(
        n_T_442[52]), .Y(n136) );
  NAND2X0_LVT U187 ( .A1(subtractor[48]), .A2(n754), .Y(n137) );
  NAND2X0_LVT U188 ( .A1(n655), .A2(io_req_bits_in2[48]), .Y(n138) );
  NAND3X0_LVT U189 ( .A1(n137), .A2(n633), .A3(n138), .Y(N371) );
  NAND2X0_LVT U190 ( .A1(n655), .A2(io_req_bits_in2[59]), .Y(n139) );
  NAND2X0_LVT U191 ( .A1(subtractor[59]), .A2(n754), .Y(n140) );
  NAND3X0_LVT U192 ( .A1(n140), .A2(n633), .A3(n139), .Y(N382) );
  NAND2X0_LVT U193 ( .A1(n_T_69[8]), .A2(n803), .Y(n141) );
  HADDX1_LVT U194 ( .A0(n141), .B0(n155), .SO(n_T_97_6_) );
  NAND2X4_LVT U195 ( .A1(n616), .A2(n615), .Y(n633) );
  NAND2X4_LVT U196 ( .A1(io_req_bits_in1[31]), .A2(n337), .Y(n658) );
  INVX1_LVT U197 ( .A(n655), .Y(n222) );
  INVX1_LVT U198 ( .A(n1000), .Y(n744) );
  INVX1_LVT U199 ( .A(io_req_bits_fn[1]), .Y(n785) );
  INVX1_LVT U200 ( .A(io_req_bits_fn[0]), .Y(n786) );
  INVX1_LVT U201 ( .A(io_req_bits_dw), .Y(n787) );
  INVX1_LVT U202 ( .A(io_req_bits_fn[2]), .Y(n784) );
  INVX1_LVT U203 ( .A(reset), .Y(n309) );
  INVX0_LVT U204 ( .A(n_T_434[5]), .Y(n170) );
  INVX0_LVT U205 ( .A(n_T_434[4]), .Y(n169) );
  INVX0_LVT U206 ( .A(n_T_434[3]), .Y(n168) );
  INVX0_LVT U207 ( .A(subtractor[64]), .Y(n310) );
  INVX0_LVT U208 ( .A(n753), .Y(n327) );
  NOR2X1_LVT U209 ( .A1(n320), .A2(io_kill), .Y(n753) );
  INVX0_LVT U210 ( .A(n957), .Y(n963) );
  INVX0_LVT U211 ( .A(n763), .Y(n968) );
  INVX0_LVT U212 ( .A(n338), .Y(n333) );
  NOR2X1_LVT U213 ( .A1(n_T_273_5_), .A2(n940), .Y(n763) );
  NOR4X0_LVT U214 ( .A1(n974), .A2(n973), .A3(n997), .A4(n_T_430_5_), .Y(n1001) );
  INVX0_LVT U215 ( .A(n956), .Y(n969) );
  MUX21X1_LVT U216 ( .A1(io_req_bits_in2[31]), .A2(io_req_bits_in2[63]), .S0(
        io_req_bits_dw), .Y(n324) );
  INVX0_LVT U217 ( .A(n1002), .Y(n972) );
  INVX0_LVT U218 ( .A(n615), .Y(n312) );
  INVX0_LVT U219 ( .A(n966), .Y(n723) );
  INVX0_LVT U220 ( .A(n967), .Y(n216) );
  INVX0_LVT U221 ( .A(n777), .Y(n974) );
  INVX0_LVT U222 ( .A(n788), .Y(n605) );
  INVX0_LVT U223 ( .A(n331), .Y(n614) );
  NOR2X1_LVT U224 ( .A1(divisor[43]), .A2(divisor[41]), .Y(n686) );
  NOR2X1_LVT U225 ( .A1(divisor[11]), .A2(divisor[9]), .Y(n699) );
  NOR2X1_LVT U226 ( .A1(divisor[27]), .A2(divisor[25]), .Y(n687) );
  NBUFFX2_LVT U227 ( .A(net34684), .Y(n299) );
  NBUFFX2_LVT U228 ( .A(net34684), .Y(n289) );
  NBUFFX2_LVT U229 ( .A(net34684), .Y(n294) );
  NBUFFX2_LVT U230 ( .A(net34684), .Y(n297) );
  NBUFFX2_LVT U231 ( .A(net34684), .Y(n295) );
  NBUFFX2_LVT U232 ( .A(net34684), .Y(n298) );
  NBUFFX2_LVT U233 ( .A(net34705), .Y(n288) );
  NBUFFX2_LVT U234 ( .A(net34705), .Y(n287) );
  NBUFFX2_LVT U235 ( .A(net34705), .Y(n285) );
  NBUFFX2_LVT U236 ( .A(net34705), .Y(n280) );
  NBUFFX2_LVT U237 ( .A(net34705), .Y(n279) );
  NBUFFX2_LVT U238 ( .A(net34705), .Y(n276) );
  NBUFFX2_LVT U239 ( .A(net34705), .Y(n271) );
  NBUFFX2_LVT U240 ( .A(net34705), .Y(n265) );
  NBUFFX2_LVT U241 ( .A(net34705), .Y(n253) );
  NBUFFX2_LVT U242 ( .A(net34705), .Y(n262) );
  NBUFFX2_LVT U243 ( .A(net34705), .Y(n245) );
  INVX1_LVT U244 ( .A(n207), .Y(n226) );
  AND2X1_LVT U245 ( .A1(subtractor[64]), .A2(n227), .Y(n931) );
  AND2X1_LVT U246 ( .A1(n235), .A2(io_req_bits_dw), .Y(n655) );
  AND2X1_LVT U247 ( .A1(n789), .A2(n605), .Y(n_T_85[5]) );
  INVX1_LVT U248 ( .A(n201), .Y(n223) );
  INVX1_LVT U249 ( .A(n200), .Y(n227) );
  OAI21X1_LVT U250 ( .A1(n980), .A2(n344), .A3(n343), .Y(n200) );
  INVX1_LVT U251 ( .A(n_T_434[0]), .Y(n171) );
  INVX1_LVT U252 ( .A(n_T_434[1]), .Y(n166) );
  INVX1_LVT U253 ( .A(n_T_434[2]), .Y(n167) );
  NBUFFX2_LVT U254 ( .A(n157), .Y(n225) );
  OR3X1_LVT U255 ( .A1(n970), .A2(n972), .A3(n998), .Y(n_T_430_5_) );
  INVX1_LVT U256 ( .A(n775), .Y(n997) );
  NBUFFX2_LVT U257 ( .A(n_T_59_8_), .Y(n301) );
  AND2X1_LVT U258 ( .A1(n224), .A2(n217), .Y(n754) );
  AND2X1_LVT U259 ( .A1(n333), .A2(n783), .Y(n679) );
  OR2X1_LVT U260 ( .A1(n_T_69[9]), .A2(n321), .Y(n980) );
  AND2X1_LVT U261 ( .A1(n774), .A2(n683), .Y(n773) );
  AND2X1_LVT U262 ( .A1(n750), .A2(n220), .Y(n783) );
  INVX1_LVT U263 ( .A(n203), .Y(n224) );
  INVX1_LVT U264 ( .A(n199), .Y(n235) );
  MUX21X1_LVT U265 ( .A1(n_T_51[16]), .A2(n_T_51[80]), .S0(n308), .Y(
        result[16]) );
  MUX21X1_LVT U266 ( .A1(n_T_51[24]), .A2(n_T_51[88]), .S0(n308), .Y(
        result[24]) );
  MUX21X1_LVT U267 ( .A1(n_T_51[51]), .A2(n_T_51[115]), .S0(n308), .Y(
        result[51]) );
  MUX21X1_LVT U268 ( .A1(n_T_51[56]), .A2(n_T_51[120]), .S0(n308), .Y(
        result[56]) );
  MUX21X1_LVT U269 ( .A1(n_T_51[33]), .A2(n_T_51[97]), .S0(n308), .Y(
        result[33]) );
  MUX21X1_LVT U270 ( .A1(n_T_51[37]), .A2(n_T_51[101]), .S0(n308), .Y(
        result[37]) );
  MUX21X1_LVT U271 ( .A1(n_T_51[48]), .A2(n_T_51[112]), .S0(n308), .Y(
        result[48]) );
  MUX21X1_LVT U272 ( .A1(n_T_51[47]), .A2(n_T_51[111]), .S0(n308), .Y(
        result[47]) );
  MUX21X1_LVT U273 ( .A1(n_T_51[57]), .A2(n_T_51[121]), .S0(n308), .Y(
        result[57]) );
  MUX21X1_LVT U274 ( .A1(n_T_51[58]), .A2(n_T_51[122]), .S0(n308), .Y(
        result[58]) );
  MUX21X1_LVT U275 ( .A1(n_T_51[14]), .A2(n_T_51[78]), .S0(n308), .Y(
        result[14]) );
  MUX21X1_LVT U276 ( .A1(n_T_51[46]), .A2(n_T_51[110]), .S0(n308), .Y(
        result[46]) );
  MUX21X1_LVT U277 ( .A1(n_T_51[40]), .A2(n_T_51[104]), .S0(n308), .Y(
        result[40]) );
  MUX21X1_LVT U278 ( .A1(n_T_51[49]), .A2(n_T_51[113]), .S0(n308), .Y(
        result[49]) );
  MUX21X1_LVT U279 ( .A1(n_T_51[52]), .A2(n_T_51[116]), .S0(n308), .Y(
        result[52]) );
  MUX21X1_LVT U280 ( .A1(n_T_51[53]), .A2(n_T_51[117]), .S0(n308), .Y(
        result[53]) );
  MUX21X1_LVT U281 ( .A1(n_T_51[42]), .A2(n_T_51[106]), .S0(n308), .Y(
        result[42]) );
  INVX1_LVT U282 ( .A(n156), .Y(n242) );
  MUX21X1_LVT U283 ( .A1(n_T_51[45]), .A2(n_T_51[109]), .S0(n308), .Y(
        result[45]) );
  MUX21X1_LVT U284 ( .A1(n_T_51[39]), .A2(n_T_51[103]), .S0(n308), .Y(
        result[39]) );
  MUX21X1_LVT U285 ( .A1(n_T_51[38]), .A2(n_T_51[102]), .S0(n308), .Y(
        result[38]) );
  MUX21X1_LVT U286 ( .A1(n_T_51[41]), .A2(n_T_51[105]), .S0(n308), .Y(
        result[41]) );
  MUX21X1_LVT U287 ( .A1(n_T_51[44]), .A2(n_T_51[108]), .S0(n308), .Y(
        result[44]) );
  INVX1_LVT U288 ( .A(n208), .Y(n304) );
  MUX21X1_LVT U289 ( .A1(n_T_51[34]), .A2(n_T_51[98]), .S0(n308), .Y(
        result[34]) );
  MUX21X1_LVT U290 ( .A1(n_T_51[43]), .A2(n_T_51[107]), .S0(n308), .Y(
        result[43]) );
  MUX21X1_LVT U291 ( .A1(n_T_51[60]), .A2(n_T_51[124]), .S0(n308), .Y(
        result[60]) );
  MUX21X1_LVT U292 ( .A1(n_T_51[36]), .A2(n_T_51[100]), .S0(n308), .Y(
        result[36]) );
  MUX21X1_LVT U293 ( .A1(n_T_51[32]), .A2(n_T_51[96]), .S0(n308), .Y(
        result[32]) );
  MUX21X1_LVT U294 ( .A1(n_T_51[54]), .A2(n_T_51[118]), .S0(n308), .Y(
        result[54]) );
  MUX21X1_LVT U295 ( .A1(n_T_51[30]), .A2(n_T_51[94]), .S0(n308), .Y(
        result[30]) );
  MUX21X1_LVT U296 ( .A1(n_T_51[62]), .A2(n_T_51[126]), .S0(n308), .Y(
        result[62]) );
  AO22X1_LVT U297 ( .A1(n146), .A2(result[63]), .A3(n209), .A4(result[31]), 
        .Y(io_resp_bits_data[31]) );
  MUX21X1_LVT U298 ( .A1(n_T_51[31]), .A2(n_T_51[95]), .S0(n308), .Y(
        result[31]) );
  MUX21X1_LVT U299 ( .A1(n_T_51[63]), .A2(n_T_51[127]), .S0(n308), .Y(
        result[63]) );
  MUX21X1_LVT U300 ( .A1(n_T_51[59]), .A2(n_T_51[123]), .S0(n308), .Y(
        result[59]) );
  MUX21X1_LVT U301 ( .A1(n_T_51[55]), .A2(n_T_51[119]), .S0(n308), .Y(
        result[55]) );
  MUX21X1_LVT U302 ( .A1(n_T_51[61]), .A2(n_T_51[125]), .S0(n308), .Y(
        result[61]) );
  MUX21X1_LVT U303 ( .A1(n_T_51[50]), .A2(n_T_51[114]), .S0(n308), .Y(
        result[50]) );
  NBUFFX2_LVT U304 ( .A(resHi), .Y(n308) );
  NAND2X0_LVT U305 ( .A1(n220), .A2(n244), .Y(n209) );
  INVX1_LVT U306 ( .A(n206), .Y(n244) );
  XOR2X2_LVT U307 ( .A1(n300), .A2(n_T_69[4]), .Y(n_T_85[4]) );
  NAND2X0_LVT U308 ( .A1(n150), .A2(n219), .Y(n203) );
  AND2X1_LVT U309 ( .A1(n750), .A2(n150), .Y(n343) );
  NAND2X0_LVT U310 ( .A1(io_req_valid), .A2(io_req_ready), .Y(n199) );
  NOR4X1_LVT U311 ( .A1(n978), .A2(n977), .A3(n235), .A4(n782), .Y(n979) );
  INVX1_LVT U312 ( .A(n804), .Y(n803) );
  INVX1_LVT U313 ( .A(n990), .Y(n1003) );
  INVX1_LVT U314 ( .A(n_T_430_5_), .Y(n976) );
  INVX1_LVT U315 ( .A(n_T_273_5_), .Y(n965) );
  AND4X1_LVT U316 ( .A1(n758), .A2(n983), .A3(n982), .A4(n981), .Y(n151) );
  NBUFFX2_LVT U317 ( .A(n_T_51[6]), .Y(n307) );
  AOI22X1_LVT U318 ( .A1(n976), .A2(n997), .A3(n1001), .A4(n1000), .Y(n158) );
  INVX1_LVT U319 ( .A(n783), .Y(n230) );
  NBUFFX2_LVT U320 ( .A(n_T_51[0]), .Y(n302) );
  NBUFFX2_LVT U321 ( .A(n_T_51[3]), .Y(n305) );
  NBUFFX2_LVT U322 ( .A(n_T_51[1]), .Y(n303) );
  NBUFFX2_LVT U323 ( .A(n_T_51[4]), .Y(n306) );
  NAND2X0_LVT U324 ( .A1(n783), .A2(n338), .Y(n201) );
  AOI22X1_LVT U325 ( .A1(n965), .A2(n964), .A3(n963), .A4(n962), .Y(n211) );
  AOI22X1_LVT U326 ( .A1(n1002), .A2(n995), .A3(n1003), .A4(n994), .Y(n213) );
  NAND2X0_LVT U327 ( .A1(n1001), .A2(n996), .Y(n214) );
  NAND3X0_LVT U328 ( .A1(n213), .A2(n151), .A3(n214), .Y(n_T_429[0]) );
  NAND2X0_LVT U329 ( .A1(n1002), .A2(n999), .Y(n215) );
  NAND3X0_LVT U330 ( .A1(n158), .A2(n773), .A3(n215), .Y(n_T_429[3]) );
  NAND2X0_LVT U331 ( .A1(n969), .A2(n966), .Y(n218) );
  NAND3X0_LVT U332 ( .A1(n211), .A2(n216), .A3(n218), .Y(n_T_272[3]) );
  NAND2X0_LVT U333 ( .A1(n210), .A2(n795), .Y(n221) );
  NAND3X0_LVT U334 ( .A1(n800), .A2(n805), .A3(n221), .Y(n798) );
  AND2X1_LVT U335 ( .A1(n184), .A2(n217), .Y(n750) );
  NAND3X0_LVT U336 ( .A1(n204), .A2(n148), .A3(n210), .Y(n789) );
  OR2X1_LVT U337 ( .A1(n_T_69[6]), .A2(n_T_69[7]), .Y(n331) );
  OR3X1_LVT U338 ( .A1(n_T_69[8]), .A2(n331), .A3(n789), .Y(n321) );
  INVX1_LVT U339 ( .A(n980), .Y(n342) );
  NAND4X0_LVT U340 ( .A1(n310), .A2(n342), .A3(n150), .A4(n189), .Y(n311) );
  AND3X1_LVT U341 ( .A1(n219), .A2(n220), .A3(n217), .Y(io_req_ready) );
  NAND3X0_LVT U342 ( .A1(n311), .A2(neg_out), .A3(n199), .Y(n318) );
  AND2X1_LVT U343 ( .A1(n235), .A2(n787), .Y(n615) );
  OA22X1_LVT U344 ( .A1(n222), .A2(io_req_bits_in1[63]), .A3(n312), .A4(
        io_req_bits_in1[31]), .Y(n316) );
  MUX21X1_LVT U345 ( .A1(io_req_bits_in1[31]), .A2(io_req_bits_in1[63]), .S0(
        io_req_bits_dw), .Y(n313) );
  AO21X1_LVT U346 ( .A1(n784), .A2(n785), .A3(n786), .Y(n336) );
  AND2X1_LVT U347 ( .A1(n313), .A2(n336), .Y(n325) );
  NAND2X0_LVT U348 ( .A1(n325), .A2(n235), .Y(n315) );
  NAND3X0_LVT U349 ( .A1(n324), .A2(n786), .A3(n785), .Y(n314) );
  MUX21X1_LVT U350 ( .A1(n316), .A2(n315), .S0(n314), .Y(n317) );
  NAND2X0_LVT U351 ( .A1(n318), .A2(n317), .Y(n793) );
  AND2X1_LVT U352 ( .A1(n184), .A2(n154), .Y(io_resp_valid) );
  NAND2X0_LVT U353 ( .A1(io_resp_ready), .A2(io_resp_valid), .Y(n319) );
  NAND3X0_LVT U354 ( .A1(n319), .A2(n199), .A3(n309), .Y(n320) );
  INVX1_LVT U355 ( .A(n321), .Y(n322) );
  AND3X1_LVT U356 ( .A1(n322), .A2(n_T_69[9]), .A3(n343), .Y(n782) );
  AND2X1_LVT U357 ( .A1(n753), .A2(n782), .Y(n680) );
  NAND2X0_LVT U358 ( .A1(n680), .A2(n212), .Y(n330) );
  MUX21X1_LVT U359 ( .A1(n785), .A2(n786), .S0(io_req_bits_fn[2]), .Y(n323) );
  AND2X1_LVT U360 ( .A1(n324), .A2(n323), .Y(n616) );
  OA21X1_LVT U361 ( .A1(n325), .A2(n616), .A3(io_req_bits_fn[2]), .Y(n326) );
  OR3X1_LVT U362 ( .A1(reset), .A2(n199), .A3(n326), .Y(n329) );
  AO21X1_LVT U363 ( .A1(n203), .A2(n230), .A3(n327), .Y(n328) );
  NAND3X0_LVT U364 ( .A1(n330), .A2(n329), .A3(n328), .Y(N284) );
  NAND2X0_LVT U365 ( .A1(n792), .A2(subtractor[64]), .Y(n344) );
  NAND2X0_LVT U366 ( .A1(n_T_69[4]), .A2(n300), .Y(n795) );
  OR2X1_LVT U367 ( .A1(n210), .A2(n795), .Y(n800) );
  INVX1_LVT U368 ( .A(n800), .Y(n778) );
  NOR2X0_LVT U369 ( .A1(n_T_69[9]), .A2(n_T_69[8]), .Y(n613) );
  NAND3X0_LVT U370 ( .A1(n778), .A2(n614), .A3(n613), .Y(n790) );
  AO222X1_LVT U371 ( .A1(n783), .A2(n_T_65[70]), .A3(subtractor[62]), .A4(n226), .A5(n_T_51[125]), .A6(n931), .Y(N522) );
  INVX1_LVT U372 ( .A(n790), .Y(n334) );
  AND4X1_LVT U373 ( .A1(n147), .A2(n186), .A3(n153), .A4(n286), .Y(n332) );
  AND4X1_LVT U374 ( .A1(n283), .A2(n281), .A3(n284), .A4(n282), .Y(n780) );
  NAND2X0_LVT U375 ( .A1(n332), .A2(n780), .Y(n1000) );
  AND4X1_LVT U376 ( .A1(n290), .A2(n293), .A3(n292), .A4(n291), .Y(n781) );
  AND4X1_LVT U377 ( .A1(n182), .A2(n243), .A3(n240), .A4(n241), .Y(n732) );
  AND4X1_LVT U378 ( .A1(n236), .A2(n239), .A3(n238), .A4(n237), .Y(n779) );
  AO21X1_LVT U379 ( .A1(n783), .A2(n334), .A3(n679), .Y(n978) );
  NOR2X0_LVT U380 ( .A1(n782), .A2(n978), .Y(n752) );
  INVX1_LVT U381 ( .A(n752), .Y(n335) );
  AO22X1_LVT U382 ( .A1(isHi), .A2(n335), .A3(n308), .A4(n979), .Y(n794) );
  NAND2X0_LVT U383 ( .A1(negated_remainder[58]), .A2(n224), .Y(n348) );
  NAND2X0_LVT U384 ( .A1(n_T_87[58]), .A2(n679), .Y(n341) );
  AND3X1_LVT U385 ( .A1(n235), .A2(n787), .A3(n336), .Y(n337) );
  NAND2X0_LVT U386 ( .A1(n223), .A2(n_T_65[2]), .Y(n340) );
  NAND2X0_LVT U387 ( .A1(n655), .A2(io_req_bits_in1[58]), .Y(n339) );
  AND4X1_LVT U388 ( .A1(n341), .A2(n658), .A3(n340), .A4(n339), .Y(n347) );
  NAND2X0_LVT U389 ( .A1(n_T_442[58]), .A2(n225), .Y(n346) );
  NAND2X0_LVT U390 ( .A1(n227), .A2(n_T_51[57]), .Y(n345) );
  NAND4X0_LVT U391 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(N452) );
  NAND2X0_LVT U392 ( .A1(negated_remainder[59]), .A2(n224), .Y(n355) );
  NAND2X0_LVT U393 ( .A1(n_T_65[3]), .A2(n223), .Y(n351) );
  NAND2X0_LVT U394 ( .A1(n_T_87[59]), .A2(n679), .Y(n350) );
  NAND2X0_LVT U395 ( .A1(n655), .A2(io_req_bits_in1[59]), .Y(n349) );
  AND4X1_LVT U396 ( .A1(n351), .A2(n658), .A3(n350), .A4(n349), .Y(n354) );
  NAND2X0_LVT U397 ( .A1(n227), .A2(n_T_51[58]), .Y(n353) );
  NAND2X0_LVT U398 ( .A1(n_T_442[59]), .A2(n157), .Y(n352) );
  NAND4X0_LVT U399 ( .A1(n355), .A2(n354), .A3(n353), .A4(n352), .Y(N453) );
  NAND2X0_LVT U400 ( .A1(negated_remainder[60]), .A2(n224), .Y(n362) );
  NAND2X0_LVT U401 ( .A1(n_T_65[4]), .A2(n223), .Y(n358) );
  NAND2X0_LVT U402 ( .A1(n_T_87[60]), .A2(n679), .Y(n357) );
  NAND2X0_LVT U403 ( .A1(n655), .A2(io_req_bits_in1[60]), .Y(n356) );
  AND4X1_LVT U404 ( .A1(n358), .A2(n658), .A3(n357), .A4(n356), .Y(n361) );
  NAND2X0_LVT U405 ( .A1(n227), .A2(n_T_51[59]), .Y(n360) );
  NAND2X0_LVT U406 ( .A1(n_T_442[60]), .A2(n225), .Y(n359) );
  NAND4X0_LVT U407 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .Y(N454) );
  NAND2X0_LVT U408 ( .A1(negated_remainder[61]), .A2(n224), .Y(n369) );
  NAND2X0_LVT U409 ( .A1(n_T_65[5]), .A2(n223), .Y(n365) );
  NAND2X0_LVT U410 ( .A1(n_T_87[61]), .A2(n679), .Y(n364) );
  NAND2X0_LVT U411 ( .A1(n655), .A2(io_req_bits_in1[61]), .Y(n363) );
  AND4X1_LVT U412 ( .A1(n365), .A2(n658), .A3(n364), .A4(n363), .Y(n368) );
  NAND2X0_LVT U413 ( .A1(n227), .A2(n_T_51[60]), .Y(n367) );
  NAND2X0_LVT U414 ( .A1(n_T_442[61]), .A2(n225), .Y(n366) );
  NAND4X0_LVT U415 ( .A1(n369), .A2(n368), .A3(n367), .A4(n366), .Y(N455) );
  NAND2X0_LVT U416 ( .A1(n_T_442[50]), .A2(n225), .Y(n376) );
  NAND2X0_LVT U417 ( .A1(n_T_87[50]), .A2(n679), .Y(n372) );
  NAND2X0_LVT U418 ( .A1(n223), .A2(n_T_51[58]), .Y(n371) );
  NAND2X0_LVT U419 ( .A1(n655), .A2(io_req_bits_in1[50]), .Y(n370) );
  AND4X1_LVT U420 ( .A1(n372), .A2(n658), .A3(n371), .A4(n370), .Y(n375) );
  NAND2X0_LVT U421 ( .A1(n227), .A2(n_T_51[49]), .Y(n374) );
  NAND2X0_LVT U422 ( .A1(negated_remainder[50]), .A2(n224), .Y(n373) );
  NAND4X0_LVT U423 ( .A1(n376), .A2(n375), .A3(n374), .A4(n373), .Y(N444) );
  NAND2X0_LVT U424 ( .A1(n_T_442[51]), .A2(n225), .Y(n383) );
  NAND2X0_LVT U425 ( .A1(n_T_87[51]), .A2(n679), .Y(n379) );
  NAND2X0_LVT U426 ( .A1(n223), .A2(n_T_51[59]), .Y(n378) );
  NAND2X0_LVT U427 ( .A1(n655), .A2(io_req_bits_in1[51]), .Y(n377) );
  AND4X1_LVT U428 ( .A1(n379), .A2(n658), .A3(n378), .A4(n377), .Y(n382) );
  NAND2X0_LVT U429 ( .A1(n227), .A2(n_T_51[50]), .Y(n381) );
  NAND2X0_LVT U430 ( .A1(negated_remainder[51]), .A2(n224), .Y(n380) );
  NAND4X0_LVT U431 ( .A1(n383), .A2(n382), .A3(n381), .A4(n380), .Y(N445) );
  NAND2X0_LVT U432 ( .A1(n_T_442[53]), .A2(n225), .Y(n390) );
  NAND2X0_LVT U433 ( .A1(n_T_87[53]), .A2(n679), .Y(n386) );
  NAND2X0_LVT U434 ( .A1(n223), .A2(n_T_51[61]), .Y(n385) );
  NAND2X0_LVT U435 ( .A1(n655), .A2(io_req_bits_in1[53]), .Y(n384) );
  AND4X1_LVT U436 ( .A1(n386), .A2(n658), .A3(n385), .A4(n384), .Y(n389) );
  NAND2X0_LVT U437 ( .A1(n227), .A2(n_T_51[52]), .Y(n388) );
  NAND2X0_LVT U438 ( .A1(negated_remainder[53]), .A2(n224), .Y(n387) );
  NAND4X0_LVT U439 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .Y(N447) );
  NAND2X0_LVT U440 ( .A1(n_T_442[54]), .A2(n157), .Y(n397) );
  NAND2X0_LVT U441 ( .A1(n_T_87[54]), .A2(n679), .Y(n393) );
  NAND2X0_LVT U442 ( .A1(n223), .A2(n_T_51[62]), .Y(n392) );
  NAND2X0_LVT U443 ( .A1(n655), .A2(io_req_bits_in1[54]), .Y(n391) );
  AND4X1_LVT U444 ( .A1(n393), .A2(n658), .A3(n392), .A4(n391), .Y(n396) );
  NAND2X0_LVT U445 ( .A1(n227), .A2(n_T_51[53]), .Y(n395) );
  NAND2X0_LVT U446 ( .A1(negated_remainder[54]), .A2(n224), .Y(n394) );
  NAND4X0_LVT U447 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .Y(N448) );
  NAND2X0_LVT U448 ( .A1(n_T_442[55]), .A2(n157), .Y(n404) );
  NAND2X0_LVT U449 ( .A1(n_T_87[55]), .A2(n679), .Y(n400) );
  NAND2X0_LVT U450 ( .A1(n223), .A2(n_T_51[63]), .Y(n399) );
  NAND2X0_LVT U451 ( .A1(n655), .A2(io_req_bits_in1[55]), .Y(n398) );
  AND4X1_LVT U452 ( .A1(n400), .A2(n658), .A3(n399), .A4(n398), .Y(n403) );
  NAND2X0_LVT U453 ( .A1(n227), .A2(n_T_51[54]), .Y(n402) );
  NAND2X0_LVT U454 ( .A1(negated_remainder[55]), .A2(n224), .Y(n401) );
  NAND4X0_LVT U455 ( .A1(n404), .A2(n403), .A3(n402), .A4(n401), .Y(N449) );
  NAND2X0_LVT U456 ( .A1(n_T_442[42]), .A2(n225), .Y(n411) );
  NAND2X0_LVT U457 ( .A1(n_T_87[42]), .A2(n679), .Y(n407) );
  NAND2X0_LVT U458 ( .A1(n223), .A2(n_T_51[50]), .Y(n406) );
  NAND2X0_LVT U459 ( .A1(n655), .A2(io_req_bits_in1[42]), .Y(n405) );
  AND4X1_LVT U460 ( .A1(n407), .A2(n658), .A3(n406), .A4(n405), .Y(n410) );
  NAND2X0_LVT U461 ( .A1(n227), .A2(n_T_51[41]), .Y(n409) );
  NAND2X0_LVT U462 ( .A1(negated_remainder[42]), .A2(n224), .Y(n408) );
  NAND4X0_LVT U463 ( .A1(n411), .A2(n410), .A3(n409), .A4(n408), .Y(N436) );
  NAND2X0_LVT U464 ( .A1(n_T_442[43]), .A2(n225), .Y(n418) );
  NAND2X0_LVT U465 ( .A1(n_T_87[43]), .A2(n679), .Y(n414) );
  NAND2X0_LVT U466 ( .A1(n223), .A2(n_T_51[51]), .Y(n413) );
  NAND2X0_LVT U467 ( .A1(n655), .A2(io_req_bits_in1[43]), .Y(n412) );
  AND4X1_LVT U468 ( .A1(n414), .A2(n658), .A3(n413), .A4(n412), .Y(n417) );
  NAND2X0_LVT U469 ( .A1(n227), .A2(n_T_51[42]), .Y(n416) );
  NAND2X0_LVT U470 ( .A1(negated_remainder[43]), .A2(n224), .Y(n415) );
  NAND4X0_LVT U471 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .Y(N437) );
  NAND2X0_LVT U472 ( .A1(n_T_442[44]), .A2(n225), .Y(n425) );
  NAND2X0_LVT U473 ( .A1(n_T_87[44]), .A2(n679), .Y(n421) );
  NAND2X0_LVT U474 ( .A1(n223), .A2(n_T_51[52]), .Y(n420) );
  NAND2X0_LVT U475 ( .A1(n655), .A2(io_req_bits_in1[44]), .Y(n419) );
  AND4X1_LVT U476 ( .A1(n421), .A2(n658), .A3(n420), .A4(n419), .Y(n424) );
  NAND2X0_LVT U477 ( .A1(n227), .A2(n_T_51[43]), .Y(n423) );
  NAND2X0_LVT U478 ( .A1(negated_remainder[44]), .A2(n224), .Y(n422) );
  NAND4X0_LVT U479 ( .A1(n425), .A2(n424), .A3(n423), .A4(n422), .Y(N438) );
  NAND2X0_LVT U480 ( .A1(n_T_442[45]), .A2(n225), .Y(n432) );
  NAND2X0_LVT U481 ( .A1(n_T_87[45]), .A2(n679), .Y(n428) );
  NAND2X0_LVT U482 ( .A1(n223), .A2(n_T_51[53]), .Y(n427) );
  NAND2X0_LVT U483 ( .A1(n655), .A2(io_req_bits_in1[45]), .Y(n426) );
  AND4X1_LVT U484 ( .A1(n428), .A2(n658), .A3(n427), .A4(n426), .Y(n431) );
  NAND2X0_LVT U485 ( .A1(n227), .A2(n_T_51[44]), .Y(n430) );
  NAND2X0_LVT U486 ( .A1(negated_remainder[45]), .A2(n224), .Y(n429) );
  NAND4X0_LVT U487 ( .A1(n432), .A2(n431), .A3(n430), .A4(n429), .Y(N439) );
  NAND2X0_LVT U488 ( .A1(n_T_442[46]), .A2(n225), .Y(n439) );
  NAND2X0_LVT U489 ( .A1(n_T_87[46]), .A2(n679), .Y(n435) );
  NAND2X0_LVT U490 ( .A1(n223), .A2(n_T_51[54]), .Y(n434) );
  NAND2X0_LVT U491 ( .A1(n655), .A2(io_req_bits_in1[46]), .Y(n433) );
  AND4X1_LVT U492 ( .A1(n435), .A2(n658), .A3(n434), .A4(n433), .Y(n438) );
  NAND2X0_LVT U493 ( .A1(n227), .A2(n_T_51[45]), .Y(n437) );
  NAND2X0_LVT U494 ( .A1(negated_remainder[46]), .A2(n224), .Y(n436) );
  NAND4X0_LVT U495 ( .A1(n439), .A2(n438), .A3(n437), .A4(n436), .Y(N440) );
  NAND2X0_LVT U496 ( .A1(n_T_442[47]), .A2(n225), .Y(n446) );
  NAND2X0_LVT U497 ( .A1(n_T_87[47]), .A2(n679), .Y(n442) );
  NAND2X0_LVT U498 ( .A1(n223), .A2(n_T_51[55]), .Y(n441) );
  NAND2X0_LVT U499 ( .A1(n655), .A2(io_req_bits_in1[47]), .Y(n440) );
  AND4X1_LVT U500 ( .A1(n442), .A2(n658), .A3(n441), .A4(n440), .Y(n445) );
  NAND2X0_LVT U501 ( .A1(n227), .A2(n_T_51[46]), .Y(n444) );
  NAND2X0_LVT U502 ( .A1(negated_remainder[47]), .A2(n224), .Y(n443) );
  NAND4X0_LVT U503 ( .A1(n446), .A2(n445), .A3(n444), .A4(n443), .Y(N441) );
  NAND2X0_LVT U504 ( .A1(n_T_442[34]), .A2(n225), .Y(n453) );
  NAND2X0_LVT U505 ( .A1(n_T_87[34]), .A2(n679), .Y(n449) );
  NAND2X0_LVT U506 ( .A1(n223), .A2(n_T_51[42]), .Y(n448) );
  NAND2X0_LVT U507 ( .A1(n655), .A2(io_req_bits_in1[34]), .Y(n447) );
  AND4X1_LVT U508 ( .A1(n449), .A2(n658), .A3(n448), .A4(n447), .Y(n452) );
  NAND2X0_LVT U509 ( .A1(n227), .A2(n_T_51[33]), .Y(n451) );
  NAND2X0_LVT U510 ( .A1(negated_remainder[34]), .A2(n224), .Y(n450) );
  NAND4X0_LVT U511 ( .A1(n453), .A2(n452), .A3(n451), .A4(n450), .Y(N428) );
  NAND2X0_LVT U512 ( .A1(n_T_442[35]), .A2(n157), .Y(n460) );
  NAND2X0_LVT U513 ( .A1(n_T_87[35]), .A2(n679), .Y(n456) );
  NAND2X0_LVT U514 ( .A1(n223), .A2(n_T_51[43]), .Y(n455) );
  NAND2X0_LVT U515 ( .A1(n655), .A2(io_req_bits_in1[35]), .Y(n454) );
  AND4X1_LVT U516 ( .A1(n456), .A2(n658), .A3(n455), .A4(n454), .Y(n459) );
  NAND2X0_LVT U517 ( .A1(n227), .A2(n_T_51[34]), .Y(n458) );
  NAND2X0_LVT U518 ( .A1(negated_remainder[35]), .A2(n224), .Y(n457) );
  NAND4X0_LVT U519 ( .A1(n460), .A2(n459), .A3(n458), .A4(n457), .Y(N429) );
  NAND2X0_LVT U520 ( .A1(n_T_442[36]), .A2(n225), .Y(n467) );
  NAND2X0_LVT U521 ( .A1(n_T_87[36]), .A2(n679), .Y(n463) );
  NAND2X0_LVT U522 ( .A1(n223), .A2(n_T_51[44]), .Y(n462) );
  NAND2X0_LVT U523 ( .A1(n655), .A2(io_req_bits_in1[36]), .Y(n461) );
  AND4X1_LVT U524 ( .A1(n463), .A2(n658), .A3(n462), .A4(n461), .Y(n466) );
  NAND2X0_LVT U525 ( .A1(n227), .A2(n_T_51[35]), .Y(n465) );
  NAND2X0_LVT U526 ( .A1(negated_remainder[36]), .A2(n224), .Y(n464) );
  NAND4X0_LVT U527 ( .A1(n467), .A2(n466), .A3(n465), .A4(n464), .Y(N430) );
  NAND2X0_LVT U528 ( .A1(n_T_442[37]), .A2(n157), .Y(n474) );
  NAND2X0_LVT U529 ( .A1(n_T_87[37]), .A2(n679), .Y(n470) );
  NAND2X0_LVT U530 ( .A1(n223), .A2(n_T_51[45]), .Y(n469) );
  NAND2X0_LVT U531 ( .A1(n655), .A2(io_req_bits_in1[37]), .Y(n468) );
  AND4X1_LVT U532 ( .A1(n470), .A2(n658), .A3(n469), .A4(n468), .Y(n473) );
  NAND2X0_LVT U533 ( .A1(n227), .A2(n_T_51[36]), .Y(n472) );
  NAND2X0_LVT U534 ( .A1(negated_remainder[37]), .A2(n224), .Y(n471) );
  NAND4X0_LVT U535 ( .A1(n474), .A2(n473), .A3(n472), .A4(n471), .Y(N431) );
  NAND2X0_LVT U536 ( .A1(n_T_442[38]), .A2(n225), .Y(n481) );
  NAND2X0_LVT U537 ( .A1(n_T_87[38]), .A2(n679), .Y(n477) );
  NAND2X0_LVT U538 ( .A1(n223), .A2(n_T_51[46]), .Y(n476) );
  NAND2X0_LVT U539 ( .A1(n655), .A2(io_req_bits_in1[38]), .Y(n475) );
  AND4X1_LVT U540 ( .A1(n477), .A2(n658), .A3(n476), .A4(n475), .Y(n480) );
  NAND2X0_LVT U541 ( .A1(n227), .A2(n_T_51[37]), .Y(n479) );
  NAND2X0_LVT U542 ( .A1(negated_remainder[38]), .A2(n224), .Y(n478) );
  NAND4X0_LVT U543 ( .A1(n481), .A2(n480), .A3(n479), .A4(n478), .Y(N432) );
  NAND2X0_LVT U544 ( .A1(n_T_442[39]), .A2(n225), .Y(n488) );
  NAND2X0_LVT U545 ( .A1(n_T_87[39]), .A2(n679), .Y(n484) );
  NAND2X0_LVT U546 ( .A1(n223), .A2(n_T_51[47]), .Y(n483) );
  NAND2X0_LVT U547 ( .A1(n655), .A2(io_req_bits_in1[39]), .Y(n482) );
  AND4X1_LVT U548 ( .A1(n484), .A2(n658), .A3(n483), .A4(n482), .Y(n487) );
  NAND2X0_LVT U549 ( .A1(n227), .A2(n_T_51[38]), .Y(n486) );
  NAND2X0_LVT U550 ( .A1(negated_remainder[39]), .A2(n224), .Y(n485) );
  NAND4X0_LVT U551 ( .A1(n488), .A2(n487), .A3(n486), .A4(n485), .Y(N433) );
  MUX21X1_LVT U552 ( .A1(n_T_51[35]), .A2(n_T_51[99]), .S0(n308), .Y(
        result[35]) );
  NAND2X0_LVT U553 ( .A1(n225), .A2(n_T_442[26]), .Y(n493) );
  AO22X1_LVT U554 ( .A1(n235), .A2(io_req_bits_in1[26]), .A3(n223), .A4(
        n_T_51[34]), .Y(n489) );
  AOI21X1_LVT U555 ( .A1(n679), .A2(n_T_87[26]), .A3(n489), .Y(n492) );
  NAND2X0_LVT U556 ( .A1(n227), .A2(n_T_51[25]), .Y(n491) );
  NAND2X0_LVT U557 ( .A1(negated_remainder[26]), .A2(n224), .Y(n490) );
  NAND4X0_LVT U558 ( .A1(n493), .A2(n492), .A3(n491), .A4(n490), .Y(N420) );
  NAND2X0_LVT U559 ( .A1(n225), .A2(n_T_442[27]), .Y(n498) );
  AO22X1_LVT U560 ( .A1(n235), .A2(io_req_bits_in1[27]), .A3(n223), .A4(
        n_T_51[35]), .Y(n494) );
  AOI21X1_LVT U561 ( .A1(n679), .A2(n_T_87[27]), .A3(n494), .Y(n497) );
  NAND2X0_LVT U562 ( .A1(n227), .A2(n_T_51[26]), .Y(n496) );
  NAND2X0_LVT U563 ( .A1(negated_remainder[27]), .A2(n224), .Y(n495) );
  NAND4X0_LVT U564 ( .A1(n498), .A2(n497), .A3(n496), .A4(n495), .Y(N421) );
  NAND2X0_LVT U565 ( .A1(n225), .A2(n_T_442[28]), .Y(n503) );
  AO22X1_LVT U566 ( .A1(n235), .A2(io_req_bits_in1[28]), .A3(n223), .A4(
        n_T_51[36]), .Y(n499) );
  AOI21X1_LVT U567 ( .A1(n679), .A2(n_T_87[28]), .A3(n499), .Y(n502) );
  NAND2X0_LVT U568 ( .A1(n227), .A2(n_T_51[27]), .Y(n501) );
  NAND2X0_LVT U569 ( .A1(negated_remainder[28]), .A2(n224), .Y(n500) );
  NAND4X0_LVT U570 ( .A1(n503), .A2(n502), .A3(n501), .A4(n500), .Y(N422) );
  NAND2X0_LVT U571 ( .A1(n225), .A2(n_T_442[29]), .Y(n508) );
  AO22X1_LVT U572 ( .A1(n235), .A2(io_req_bits_in1[29]), .A3(n223), .A4(
        n_T_51[37]), .Y(n504) );
  AOI21X1_LVT U573 ( .A1(n679), .A2(n_T_87[29]), .A3(n504), .Y(n507) );
  NAND2X0_LVT U574 ( .A1(n227), .A2(n_T_51[28]), .Y(n506) );
  NAND2X0_LVT U575 ( .A1(negated_remainder[29]), .A2(n224), .Y(n505) );
  NAND4X0_LVT U576 ( .A1(n508), .A2(n507), .A3(n506), .A4(n505), .Y(N423) );
  NAND2X0_LVT U577 ( .A1(n225), .A2(n_T_442[30]), .Y(n513) );
  AO22X1_LVT U578 ( .A1(n235), .A2(io_req_bits_in1[30]), .A3(n223), .A4(
        n_T_51[38]), .Y(n509) );
  AOI21X1_LVT U579 ( .A1(n679), .A2(n_T_87[30]), .A3(n509), .Y(n512) );
  NAND2X0_LVT U580 ( .A1(n227), .A2(n_T_51[29]), .Y(n511) );
  NAND2X0_LVT U581 ( .A1(negated_remainder[30]), .A2(n224), .Y(n510) );
  NAND4X0_LVT U582 ( .A1(n513), .A2(n512), .A3(n511), .A4(n510), .Y(N424) );
  NAND2X0_LVT U583 ( .A1(n225), .A2(n_T_442[31]), .Y(n518) );
  AO22X1_LVT U584 ( .A1(n235), .A2(io_req_bits_in1[31]), .A3(n223), .A4(
        n_T_51[39]), .Y(n514) );
  AOI21X1_LVT U585 ( .A1(n679), .A2(n_T_87[31]), .A3(n514), .Y(n517) );
  NAND2X0_LVT U586 ( .A1(n227), .A2(n_T_51[30]), .Y(n516) );
  NAND2X0_LVT U587 ( .A1(negated_remainder[31]), .A2(n224), .Y(n515) );
  NAND4X0_LVT U588 ( .A1(n518), .A2(n517), .A3(n516), .A4(n515), .Y(N425) );
  MUX21X1_LVT U589 ( .A1(n_T_51[29]), .A2(n_T_51[93]), .S0(n308), .Y(
        result[29]) );
  MUX21X1_LVT U590 ( .A1(n_T_51[28]), .A2(n_T_51[92]), .S0(n308), .Y(
        result[28]) );
  MUX21X1_LVT U591 ( .A1(n_T_51[27]), .A2(n_T_51[91]), .S0(n308), .Y(
        result[27]) );
  MUX21X1_LVT U592 ( .A1(n_T_51[26]), .A2(n_T_51[90]), .S0(n308), .Y(
        result[26]) );
  MUX21X1_LVT U593 ( .A1(n_T_51[25]), .A2(n_T_51[89]), .S0(n308), .Y(
        result[25]) );
  NAND2X0_LVT U594 ( .A1(n225), .A2(n_T_442[18]), .Y(n523) );
  AO22X1_LVT U595 ( .A1(n235), .A2(io_req_bits_in1[18]), .A3(n223), .A4(
        n_T_51[26]), .Y(n519) );
  AOI21X1_LVT U596 ( .A1(n679), .A2(n_T_87[18]), .A3(n519), .Y(n522) );
  NAND2X0_LVT U597 ( .A1(n227), .A2(n_T_51[17]), .Y(n521) );
  NAND2X0_LVT U598 ( .A1(negated_remainder[18]), .A2(n224), .Y(n520) );
  NAND4X0_LVT U599 ( .A1(n523), .A2(n522), .A3(n521), .A4(n520), .Y(N412) );
  NAND2X0_LVT U600 ( .A1(n225), .A2(n_T_442[19]), .Y(n528) );
  AO22X1_LVT U601 ( .A1(n235), .A2(io_req_bits_in1[19]), .A3(n223), .A4(
        n_T_51[27]), .Y(n524) );
  AOI21X1_LVT U602 ( .A1(n679), .A2(n_T_87[19]), .A3(n524), .Y(n527) );
  NAND2X0_LVT U603 ( .A1(n227), .A2(n_T_51[18]), .Y(n526) );
  NAND2X0_LVT U604 ( .A1(negated_remainder[19]), .A2(n224), .Y(n525) );
  NAND4X0_LVT U605 ( .A1(n528), .A2(n527), .A3(n526), .A4(n525), .Y(N413) );
  NAND2X0_LVT U606 ( .A1(n225), .A2(n_T_442[20]), .Y(n533) );
  AO22X1_LVT U607 ( .A1(n235), .A2(io_req_bits_in1[20]), .A3(n223), .A4(
        n_T_51[28]), .Y(n529) );
  AOI21X1_LVT U608 ( .A1(n679), .A2(n_T_87[20]), .A3(n529), .Y(n532) );
  NAND2X0_LVT U609 ( .A1(n227), .A2(n_T_51[19]), .Y(n531) );
  NAND2X0_LVT U610 ( .A1(negated_remainder[20]), .A2(n224), .Y(n530) );
  NAND4X0_LVT U611 ( .A1(n533), .A2(n532), .A3(n531), .A4(n530), .Y(N414) );
  NAND2X0_LVT U612 ( .A1(n225), .A2(n_T_442[21]), .Y(n538) );
  AO22X1_LVT U613 ( .A1(n235), .A2(io_req_bits_in1[21]), .A3(n223), .A4(
        n_T_51[29]), .Y(n534) );
  AOI21X1_LVT U614 ( .A1(n679), .A2(n_T_87[21]), .A3(n534), .Y(n537) );
  NAND2X0_LVT U615 ( .A1(n227), .A2(n_T_51[20]), .Y(n536) );
  NAND2X0_LVT U616 ( .A1(negated_remainder[21]), .A2(n224), .Y(n535) );
  NAND4X0_LVT U617 ( .A1(n538), .A2(n537), .A3(n536), .A4(n535), .Y(N415) );
  NAND2X0_LVT U618 ( .A1(n225), .A2(n_T_442[22]), .Y(n543) );
  AO22X1_LVT U619 ( .A1(n235), .A2(io_req_bits_in1[22]), .A3(n223), .A4(
        n_T_51[30]), .Y(n539) );
  AOI21X1_LVT U620 ( .A1(n679), .A2(n_T_87[22]), .A3(n539), .Y(n542) );
  NAND2X0_LVT U621 ( .A1(n227), .A2(n_T_51[21]), .Y(n541) );
  NAND2X0_LVT U622 ( .A1(negated_remainder[22]), .A2(n224), .Y(n540) );
  NAND4X0_LVT U623 ( .A1(n543), .A2(n542), .A3(n541), .A4(n540), .Y(N416) );
  NAND2X0_LVT U624 ( .A1(n225), .A2(n_T_442[23]), .Y(n548) );
  AO22X1_LVT U625 ( .A1(n235), .A2(io_req_bits_in1[23]), .A3(n223), .A4(
        n_T_51[31]), .Y(n544) );
  AOI21X1_LVT U626 ( .A1(n679), .A2(n_T_87[23]), .A3(n544), .Y(n547) );
  NAND2X0_LVT U627 ( .A1(n227), .A2(n_T_51[22]), .Y(n546) );
  NAND2X0_LVT U628 ( .A1(negated_remainder[23]), .A2(n224), .Y(n545) );
  NAND4X0_LVT U629 ( .A1(n548), .A2(n547), .A3(n546), .A4(n545), .Y(N417) );
  MUX21X1_LVT U630 ( .A1(n_T_51[23]), .A2(n_T_51[87]), .S0(resHi), .Y(
        result[23]) );
  MUX21X1_LVT U631 ( .A1(n_T_51[22]), .A2(n_T_51[86]), .S0(resHi), .Y(
        result[22]) );
  MUX21X1_LVT U632 ( .A1(n_T_51[21]), .A2(n_T_51[85]), .S0(n308), .Y(
        result[21]) );
  MUX21X1_LVT U633 ( .A1(n_T_51[20]), .A2(n_T_51[84]), .S0(resHi), .Y(
        result[20]) );
  MUX21X1_LVT U634 ( .A1(n_T_51[19]), .A2(n_T_51[83]), .S0(n308), .Y(
        result[19]) );
  MUX21X1_LVT U635 ( .A1(n_T_51[18]), .A2(n_T_51[82]), .S0(n308), .Y(
        result[18]) );
  MUX21X1_LVT U636 ( .A1(n_T_51[17]), .A2(n_T_51[81]), .S0(n308), .Y(
        result[17]) );
  NAND2X0_LVT U637 ( .A1(n225), .A2(n_T_442[10]), .Y(n553) );
  AO22X1_LVT U638 ( .A1(n235), .A2(io_req_bits_in1[10]), .A3(n223), .A4(
        n_T_51[18]), .Y(n549) );
  AOI21X1_LVT U639 ( .A1(n679), .A2(n_T_87[10]), .A3(n549), .Y(n552) );
  NAND2X0_LVT U640 ( .A1(n227), .A2(n_T_51[9]), .Y(n551) );
  NAND2X0_LVT U641 ( .A1(negated_remainder[10]), .A2(n224), .Y(n550) );
  NAND4X0_LVT U642 ( .A1(n553), .A2(n552), .A3(n551), .A4(n550), .Y(N404) );
  NAND2X0_LVT U643 ( .A1(n225), .A2(n_T_442[11]), .Y(n558) );
  AO22X1_LVT U644 ( .A1(n235), .A2(io_req_bits_in1[11]), .A3(n223), .A4(
        n_T_51[19]), .Y(n554) );
  AOI21X1_LVT U645 ( .A1(n679), .A2(n_T_87[11]), .A3(n554), .Y(n557) );
  NAND2X0_LVT U646 ( .A1(n227), .A2(n_T_51[10]), .Y(n556) );
  NAND2X0_LVT U647 ( .A1(negated_remainder[11]), .A2(n224), .Y(n555) );
  NAND4X0_LVT U648 ( .A1(n558), .A2(n557), .A3(n556), .A4(n555), .Y(N405) );
  NAND2X0_LVT U649 ( .A1(n225), .A2(n_T_442[13]), .Y(n563) );
  AO22X1_LVT U650 ( .A1(n235), .A2(io_req_bits_in1[13]), .A3(n223), .A4(
        n_T_51[21]), .Y(n559) );
  AOI21X1_LVT U651 ( .A1(n679), .A2(n_T_87[13]), .A3(n559), .Y(n562) );
  NAND2X0_LVT U652 ( .A1(n227), .A2(n_T_51[12]), .Y(n561) );
  NAND2X0_LVT U653 ( .A1(negated_remainder[13]), .A2(n224), .Y(n560) );
  NAND4X0_LVT U654 ( .A1(n563), .A2(n562), .A3(n561), .A4(n560), .Y(N407) );
  NAND2X0_LVT U655 ( .A1(n225), .A2(n_T_442[14]), .Y(n568) );
  AO22X1_LVT U656 ( .A1(n235), .A2(io_req_bits_in1[14]), .A3(n223), .A4(
        n_T_51[22]), .Y(n564) );
  AOI21X1_LVT U657 ( .A1(n679), .A2(n_T_87[14]), .A3(n564), .Y(n567) );
  NAND2X0_LVT U658 ( .A1(n227), .A2(n_T_51[13]), .Y(n566) );
  NAND2X0_LVT U659 ( .A1(negated_remainder[14]), .A2(n224), .Y(n565) );
  NAND4X0_LVT U660 ( .A1(n568), .A2(n567), .A3(n566), .A4(n565), .Y(N408) );
  NAND2X0_LVT U661 ( .A1(n157), .A2(n_T_442[15]), .Y(n573) );
  AO22X1_LVT U662 ( .A1(n235), .A2(io_req_bits_in1[15]), .A3(n223), .A4(
        n_T_51[23]), .Y(n569) );
  AOI21X1_LVT U663 ( .A1(n679), .A2(n_T_87[15]), .A3(n569), .Y(n572) );
  NAND2X0_LVT U664 ( .A1(n227), .A2(n_T_51[14]), .Y(n571) );
  NAND2X0_LVT U665 ( .A1(negated_remainder[15]), .A2(n224), .Y(n570) );
  NAND4X0_LVT U666 ( .A1(n573), .A2(n572), .A3(n571), .A4(n570), .Y(N409) );
  MUX21X1_LVT U667 ( .A1(n_T_51[15]), .A2(n_T_51[79]), .S0(n308), .Y(
        result[15]) );
  MUX21X1_LVT U668 ( .A1(n_T_51[13]), .A2(n_T_51[77]), .S0(n308), .Y(
        result[13]) );
  MUX21X1_LVT U669 ( .A1(n_T_51[12]), .A2(n_T_51[76]), .S0(n308), .Y(
        result[12]) );
  MUX21X1_LVT U670 ( .A1(n_T_51[11]), .A2(n_T_51[75]), .S0(resHi), .Y(
        result[11]) );
  MUX21X1_LVT U671 ( .A1(n_T_51[10]), .A2(n_T_51[74]), .S0(resHi), .Y(
        result[10]) );
  MUX21X1_LVT U672 ( .A1(n_T_51[9]), .A2(n_T_51[73]), .S0(n308), .Y(result[9])
         );
  NAND2X0_LVT U673 ( .A1(n225), .A2(n_T_442[3]), .Y(n578) );
  AO22X1_LVT U674 ( .A1(n235), .A2(io_req_bits_in1[3]), .A3(
        negated_remainder[3]), .A4(n224), .Y(n574) );
  AOI21X1_LVT U675 ( .A1(n_T_51[11]), .A2(n223), .A3(n574), .Y(n577) );
  NAND2X0_LVT U676 ( .A1(n227), .A2(n304), .Y(n576) );
  NAND2X0_LVT U677 ( .A1(n_T_87[3]), .A2(n679), .Y(n575) );
  NAND4X0_LVT U678 ( .A1(n578), .A2(n577), .A3(n576), .A4(n575), .Y(N397) );
  NAND2X0_LVT U679 ( .A1(n225), .A2(n_T_442[5]), .Y(n583) );
  AO22X1_LVT U680 ( .A1(io_req_bits_in1[5]), .A2(n235), .A3(n223), .A4(
        n_T_51[13]), .Y(n579) );
  AOI21X1_LVT U681 ( .A1(n679), .A2(n_T_87[5]), .A3(n579), .Y(n582) );
  NAND2X0_LVT U682 ( .A1(n227), .A2(n_T_51[4]), .Y(n581) );
  NAND2X0_LVT U683 ( .A1(negated_remainder[5]), .A2(n224), .Y(n580) );
  NAND4X0_LVT U684 ( .A1(n583), .A2(n582), .A3(n581), .A4(n580), .Y(N399) );
  NAND2X0_LVT U685 ( .A1(n225), .A2(n_T_442[6]), .Y(n588) );
  AO22X1_LVT U686 ( .A1(io_req_bits_in1[6]), .A2(n235), .A3(n223), .A4(
        n_T_51[14]), .Y(n584) );
  AOI21X1_LVT U687 ( .A1(n679), .A2(n_T_87[6]), .A3(n584), .Y(n587) );
  NAND2X0_LVT U688 ( .A1(n227), .A2(n_T_51[5]), .Y(n586) );
  NAND2X0_LVT U689 ( .A1(negated_remainder[6]), .A2(n224), .Y(n585) );
  NAND4X0_LVT U690 ( .A1(n588), .A2(n587), .A3(n586), .A4(n585), .Y(N400) );
  NAND2X0_LVT U691 ( .A1(n157), .A2(n_T_442[7]), .Y(n593) );
  AO22X1_LVT U692 ( .A1(io_req_bits_in1[7]), .A2(n235), .A3(n223), .A4(
        n_T_51[15]), .Y(n589) );
  AOI21X1_LVT U693 ( .A1(n679), .A2(n_T_87[7]), .A3(n589), .Y(n592) );
  NAND2X0_LVT U694 ( .A1(n227), .A2(n_T_51[6]), .Y(n591) );
  NAND2X0_LVT U695 ( .A1(negated_remainder[7]), .A2(n224), .Y(n590) );
  NAND4X0_LVT U696 ( .A1(n593), .A2(n592), .A3(n591), .A4(n590), .Y(N401) );
  NAND2X0_LVT U697 ( .A1(n225), .A2(n_T_442[8]), .Y(n598) );
  AO22X1_LVT U698 ( .A1(n235), .A2(io_req_bits_in1[8]), .A3(n223), .A4(
        n_T_51[16]), .Y(n594) );
  AOI21X1_LVT U699 ( .A1(n679), .A2(n_T_87[8]), .A3(n594), .Y(n597) );
  NAND2X0_LVT U700 ( .A1(n227), .A2(n_T_51[7]), .Y(n596) );
  NAND2X0_LVT U701 ( .A1(negated_remainder[8]), .A2(n224), .Y(n595) );
  NAND4X0_LVT U702 ( .A1(n598), .A2(n597), .A3(n596), .A4(n595), .Y(N402) );
  MUX21X1_LVT U703 ( .A1(n_T_51[8]), .A2(n_T_51[72]), .S0(resHi), .Y(result[8]) );
  MUX21X1_LVT U704 ( .A1(n_T_51[7]), .A2(n_T_51[71]), .S0(n308), .Y(result[7])
         );
  MUX21X1_LVT U705 ( .A1(n_T_51[6]), .A2(n_T_51[70]), .S0(resHi), .Y(result[6]) );
  MUX21X1_LVT U706 ( .A1(n_T_51[5]), .A2(n_T_51[69]), .S0(n308), .Y(result[5])
         );
  MUX21X1_LVT U707 ( .A1(n_T_51[4]), .A2(n_T_51[68]), .S0(n308), .Y(result[4])
         );
  MUX21X1_LVT U708 ( .A1(n305), .A2(n_T_51[67]), .S0(n308), .Y(result[3]) );
  MUX21X1_LVT U709 ( .A1(n304), .A2(n_T_51[66]), .S0(n308), .Y(result[2]) );
  MUX21X1_LVT U710 ( .A1(n_T_51[1]), .A2(n_T_51[65]), .S0(n308), .Y(result[1])
         );
  MUX21X1_LVT U711 ( .A1(n302), .A2(n_T_51[64]), .S0(n308), .Y(result[0]) );
  NAND2X0_LVT U712 ( .A1(n_T_65[6]), .A2(n223), .Y(n601) );
  NAND2X0_LVT U713 ( .A1(n_T_87[62]), .A2(n679), .Y(n600) );
  NAND2X0_LVT U714 ( .A1(n655), .A2(io_req_bits_in1[62]), .Y(n599) );
  NAND4X0_LVT U715 ( .A1(n601), .A2(n658), .A3(n600), .A4(n599), .Y(n602) );
  AO21X1_LVT U716 ( .A1(n227), .A2(n_T_51[61]), .A3(n602), .Y(n603) );
  AO21X1_LVT U717 ( .A1(n225), .A2(n_T_442[62]), .A3(n603), .Y(n604) );
  AO21X1_LVT U718 ( .A1(negated_remainder[62]), .A2(n224), .A3(n604), .Y(N456)
         );
  OA21X1_LVT U719 ( .A1(n300), .A2(n_T_69[4]), .A3(n_T_71_39_), .Y(n788) );
  NAND2X0_LVT U720 ( .A1(negated_remainder[63]), .A2(n224), .Y(n612) );
  NAND2X0_LVT U721 ( .A1(n_T_65[7]), .A2(n223), .Y(n608) );
  NAND2X0_LVT U722 ( .A1(n_T_87[63]), .A2(n679), .Y(n607) );
  NAND2X0_LVT U723 ( .A1(n655), .A2(io_req_bits_in1[63]), .Y(n606) );
  AND4X1_LVT U724 ( .A1(n608), .A2(n607), .A3(n606), .A4(n658), .Y(n611) );
  NAND2X0_LVT U725 ( .A1(n227), .A2(n_T_51[62]), .Y(n610) );
  NAND2X0_LVT U726 ( .A1(n_T_442[63]), .A2(n225), .Y(n609) );
  NAND4X0_LVT U727 ( .A1(n612), .A2(n611), .A3(n610), .A4(n609), .Y(N457) );
  AO22X1_LVT U728 ( .A1(n235), .A2(n616), .A3(subtractor[64]), .A4(n754), .Y(
        N387) );
  NAND2X0_LVT U729 ( .A1(subtractor[45]), .A2(n754), .Y(n618) );
  NAND2X0_LVT U730 ( .A1(io_req_bits_in2[45]), .A2(n655), .Y(n617) );
  NAND3X0_LVT U731 ( .A1(n618), .A2(n633), .A3(n617), .Y(N368) );
  NAND2X0_LVT U732 ( .A1(subtractor[42]), .A2(n754), .Y(n620) );
  NAND2X0_LVT U733 ( .A1(io_req_bits_in2[42]), .A2(n655), .Y(n619) );
  NAND3X0_LVT U734 ( .A1(n620), .A2(n633), .A3(n619), .Y(N365) );
  NAND2X0_LVT U735 ( .A1(subtractor[39]), .A2(n754), .Y(n622) );
  NAND2X0_LVT U736 ( .A1(io_req_bits_in2[39]), .A2(n655), .Y(n621) );
  NAND3X0_LVT U737 ( .A1(n622), .A2(n633), .A3(n621), .Y(N362) );
  NAND2X0_LVT U738 ( .A1(subtractor[38]), .A2(n754), .Y(n624) );
  NAND2X0_LVT U739 ( .A1(io_req_bits_in2[38]), .A2(n655), .Y(n623) );
  NAND3X0_LVT U740 ( .A1(n624), .A2(n633), .A3(n623), .Y(N361) );
  NAND2X0_LVT U741 ( .A1(subtractor[37]), .A2(n754), .Y(n626) );
  NAND2X0_LVT U742 ( .A1(io_req_bits_in2[37]), .A2(n655), .Y(n625) );
  NAND3X0_LVT U743 ( .A1(n626), .A2(n633), .A3(n625), .Y(N360) );
  NAND2X0_LVT U744 ( .A1(subtractor[36]), .A2(n754), .Y(n628) );
  NAND2X0_LVT U745 ( .A1(io_req_bits_in2[36]), .A2(n655), .Y(n627) );
  NAND3X0_LVT U746 ( .A1(n628), .A2(n633), .A3(n627), .Y(N359) );
  NAND2X0_LVT U747 ( .A1(subtractor[34]), .A2(n754), .Y(n630) );
  NAND2X0_LVT U748 ( .A1(io_req_bits_in2[34]), .A2(n655), .Y(n629) );
  NAND3X0_LVT U749 ( .A1(n630), .A2(n633), .A3(n629), .Y(N357) );
  NAND2X0_LVT U750 ( .A1(subtractor[33]), .A2(n754), .Y(n632) );
  NAND2X0_LVT U751 ( .A1(io_req_bits_in2[33]), .A2(n655), .Y(n631) );
  NAND3X0_LVT U752 ( .A1(n632), .A2(n633), .A3(n631), .Y(N356) );
  AO22X1_LVT U753 ( .A1(n235), .A2(io_req_bits_in2[31]), .A3(subtractor[31]), 
        .A4(n754), .Y(N354) );
  AO22X1_LVT U754 ( .A1(n235), .A2(io_req_bits_in2[30]), .A3(subtractor[30]), 
        .A4(n754), .Y(N353) );
  AO22X1_LVT U755 ( .A1(n235), .A2(io_req_bits_in2[29]), .A3(subtractor[29]), 
        .A4(n754), .Y(N352) );
  AO22X1_LVT U756 ( .A1(n235), .A2(io_req_bits_in2[28]), .A3(subtractor[28]), 
        .A4(n754), .Y(N351) );
  AO22X1_LVT U757 ( .A1(n235), .A2(io_req_bits_in2[27]), .A3(subtractor[27]), 
        .A4(n754), .Y(N350) );
  AO22X1_LVT U758 ( .A1(n235), .A2(io_req_bits_in2[26]), .A3(subtractor[26]), 
        .A4(n754), .Y(N349) );
  AO22X1_LVT U759 ( .A1(n235), .A2(io_req_bits_in2[25]), .A3(subtractor[25]), 
        .A4(n754), .Y(N348) );
  AO22X1_LVT U760 ( .A1(n235), .A2(io_req_bits_in2[24]), .A3(subtractor[24]), 
        .A4(n754), .Y(N347) );
  AO22X1_LVT U761 ( .A1(n235), .A2(io_req_bits_in2[23]), .A3(subtractor[23]), 
        .A4(n754), .Y(N346) );
  AO22X1_LVT U762 ( .A1(n235), .A2(io_req_bits_in2[22]), .A3(subtractor[22]), 
        .A4(n754), .Y(N345) );
  AO22X1_LVT U763 ( .A1(n235), .A2(io_req_bits_in2[21]), .A3(subtractor[21]), 
        .A4(n754), .Y(N344) );
  AO22X1_LVT U764 ( .A1(n235), .A2(io_req_bits_in2[20]), .A3(subtractor[20]), 
        .A4(n754), .Y(N343) );
  AO22X1_LVT U765 ( .A1(n235), .A2(io_req_bits_in2[19]), .A3(subtractor[19]), 
        .A4(n754), .Y(N342) );
  AO22X1_LVT U766 ( .A1(n235), .A2(io_req_bits_in2[18]), .A3(subtractor[18]), 
        .A4(n754), .Y(N341) );
  AO22X1_LVT U767 ( .A1(n235), .A2(io_req_bits_in2[17]), .A3(subtractor[17]), 
        .A4(n754), .Y(N340) );
  AO22X1_LVT U768 ( .A1(n235), .A2(io_req_bits_in2[16]), .A3(subtractor[16]), 
        .A4(n754), .Y(N339) );
  AO22X1_LVT U769 ( .A1(n235), .A2(io_req_bits_in2[15]), .A3(subtractor[15]), 
        .A4(n754), .Y(N338) );
  AO22X1_LVT U770 ( .A1(n235), .A2(io_req_bits_in2[14]), .A3(subtractor[14]), 
        .A4(n754), .Y(N337) );
  AO22X1_LVT U771 ( .A1(n235), .A2(io_req_bits_in2[13]), .A3(subtractor[13]), 
        .A4(n754), .Y(N336) );
  AO22X1_LVT U772 ( .A1(n235), .A2(io_req_bits_in2[12]), .A3(subtractor[12]), 
        .A4(n754), .Y(N335) );
  AO22X1_LVT U773 ( .A1(n235), .A2(io_req_bits_in2[11]), .A3(subtractor[11]), 
        .A4(n754), .Y(N334) );
  AO22X1_LVT U774 ( .A1(n235), .A2(io_req_bits_in2[10]), .A3(subtractor[10]), 
        .A4(n754), .Y(N333) );
  AO22X1_LVT U775 ( .A1(n235), .A2(io_req_bits_in2[9]), .A3(subtractor[9]), 
        .A4(n754), .Y(N332) );
  AO22X1_LVT U776 ( .A1(n235), .A2(io_req_bits_in2[8]), .A3(subtractor[8]), 
        .A4(n754), .Y(N331) );
  AO22X1_LVT U777 ( .A1(n235), .A2(io_req_bits_in2[7]), .A3(subtractor[7]), 
        .A4(n754), .Y(N330) );
  AO22X1_LVT U778 ( .A1(n235), .A2(io_req_bits_in2[6]), .A3(subtractor[6]), 
        .A4(n754), .Y(N329) );
  AO22X1_LVT U779 ( .A1(n235), .A2(io_req_bits_in2[5]), .A3(subtractor[5]), 
        .A4(n754), .Y(N328) );
  AO22X1_LVT U780 ( .A1(n235), .A2(io_req_bits_in2[4]), .A3(subtractor[4]), 
        .A4(n754), .Y(N327) );
  AO22X1_LVT U781 ( .A1(n235), .A2(io_req_bits_in2[3]), .A3(subtractor[3]), 
        .A4(n754), .Y(N326) );
  AO22X1_LVT U782 ( .A1(io_req_bits_in2[2]), .A2(n235), .A3(subtractor[2]), 
        .A4(n754), .Y(N325) );
  AO22X1_LVT U783 ( .A1(n754), .A2(subtractor[1]), .A3(io_req_bits_in2[1]), 
        .A4(n235), .Y(N324) );
  AO22X1_LVT U784 ( .A1(n754), .A2(subtractor[0]), .A3(io_req_bits_in2[0]), 
        .A4(n235), .Y(N323) );
  NAND2X0_LVT U785 ( .A1(negated_remainder[57]), .A2(n224), .Y(n640) );
  NAND2X0_LVT U786 ( .A1(n_T_87[57]), .A2(n679), .Y(n636) );
  NAND2X0_LVT U787 ( .A1(n223), .A2(n_T_65[1]), .Y(n635) );
  NAND2X0_LVT U788 ( .A1(n655), .A2(io_req_bits_in1[57]), .Y(n634) );
  AND4X1_LVT U789 ( .A1(n636), .A2(n658), .A3(n635), .A4(n634), .Y(n639) );
  NAND2X0_LVT U790 ( .A1(n_T_442[57]), .A2(n225), .Y(n638) );
  NAND2X0_LVT U791 ( .A1(n227), .A2(n_T_51[56]), .Y(n637) );
  NAND4X0_LVT U792 ( .A1(n640), .A2(n639), .A3(n638), .A4(n637), .Y(N451) );
  NAND2X0_LVT U793 ( .A1(n_T_442[49]), .A2(n157), .Y(n647) );
  NAND2X0_LVT U794 ( .A1(n_T_87[49]), .A2(n679), .Y(n643) );
  NAND2X0_LVT U795 ( .A1(n223), .A2(n_T_51[57]), .Y(n642) );
  NAND2X0_LVT U796 ( .A1(n655), .A2(io_req_bits_in1[49]), .Y(n641) );
  AND4X1_LVT U797 ( .A1(n643), .A2(n658), .A3(n642), .A4(n641), .Y(n646) );
  NAND2X0_LVT U798 ( .A1(n227), .A2(n_T_51[48]), .Y(n645) );
  NAND2X0_LVT U799 ( .A1(negated_remainder[49]), .A2(n224), .Y(n644) );
  NAND4X0_LVT U800 ( .A1(n647), .A2(n646), .A3(n645), .A4(n644), .Y(N443) );
  NAND2X0_LVT U801 ( .A1(n_T_442[41]), .A2(n157), .Y(n654) );
  NAND2X0_LVT U802 ( .A1(n_T_87[41]), .A2(n679), .Y(n650) );
  NAND2X0_LVT U803 ( .A1(n223), .A2(n_T_51[49]), .Y(n649) );
  NAND2X0_LVT U804 ( .A1(n655), .A2(io_req_bits_in1[41]), .Y(n648) );
  AND4X1_LVT U805 ( .A1(n650), .A2(n658), .A3(n649), .A4(n648), .Y(n653) );
  NAND2X0_LVT U806 ( .A1(n227), .A2(n_T_51[40]), .Y(n652) );
  NAND2X0_LVT U807 ( .A1(negated_remainder[41]), .A2(n224), .Y(n651) );
  NAND4X0_LVT U808 ( .A1(n654), .A2(n653), .A3(n652), .A4(n651), .Y(N435) );
  NAND2X0_LVT U809 ( .A1(n_T_442[33]), .A2(n225), .Y(n663) );
  NAND2X0_LVT U810 ( .A1(n_T_87[33]), .A2(n679), .Y(n659) );
  NAND2X0_LVT U811 ( .A1(n223), .A2(n_T_51[41]), .Y(n657) );
  NAND2X0_LVT U812 ( .A1(n655), .A2(io_req_bits_in1[33]), .Y(n656) );
  AND4X1_LVT U813 ( .A1(n659), .A2(n658), .A3(n657), .A4(n656), .Y(n662) );
  NAND2X0_LVT U814 ( .A1(n227), .A2(n_T_51[32]), .Y(n661) );
  NAND2X0_LVT U815 ( .A1(negated_remainder[33]), .A2(n224), .Y(n660) );
  NAND4X0_LVT U816 ( .A1(n663), .A2(n662), .A3(n661), .A4(n660), .Y(N427) );
  NAND2X0_LVT U817 ( .A1(n225), .A2(n_T_442[25]), .Y(n668) );
  AO22X1_LVT U818 ( .A1(n235), .A2(io_req_bits_in1[25]), .A3(n223), .A4(
        n_T_51[33]), .Y(n664) );
  AOI21X1_LVT U819 ( .A1(n679), .A2(n_T_87[25]), .A3(n664), .Y(n667) );
  NAND2X0_LVT U820 ( .A1(n227), .A2(n_T_51[24]), .Y(n666) );
  NAND2X0_LVT U821 ( .A1(negated_remainder[25]), .A2(n224), .Y(n665) );
  NAND4X0_LVT U822 ( .A1(n668), .A2(n667), .A3(n666), .A4(n665), .Y(N419) );
  NAND2X0_LVT U823 ( .A1(n225), .A2(n_T_442[17]), .Y(n673) );
  AO22X1_LVT U824 ( .A1(n235), .A2(io_req_bits_in1[17]), .A3(n223), .A4(
        n_T_51[25]), .Y(n669) );
  AOI21X1_LVT U825 ( .A1(n679), .A2(n_T_87[17]), .A3(n669), .Y(n672) );
  NAND2X0_LVT U826 ( .A1(n227), .A2(n_T_51[16]), .Y(n671) );
  NAND2X0_LVT U827 ( .A1(negated_remainder[17]), .A2(n224), .Y(n670) );
  NAND4X0_LVT U828 ( .A1(n673), .A2(n672), .A3(n671), .A4(n670), .Y(N411) );
  NAND2X0_LVT U829 ( .A1(n157), .A2(n_T_442[9]), .Y(n678) );
  AO22X1_LVT U830 ( .A1(n235), .A2(io_req_bits_in1[9]), .A3(n223), .A4(
        n_T_51[17]), .Y(n674) );
  AOI21X1_LVT U831 ( .A1(n679), .A2(n_T_87[9]), .A3(n674), .Y(n677) );
  NAND2X0_LVT U832 ( .A1(n227), .A2(n_T_51[8]), .Y(n676) );
  NAND2X0_LVT U833 ( .A1(negated_remainder[9]), .A2(n224), .Y(n675) );
  NAND4X0_LVT U834 ( .A1(n678), .A2(n677), .A3(n676), .A4(n675), .Y(N403) );
  AND2X1_LVT U835 ( .A1(n224), .A2(n154), .Y(n977) );
  OR2X1_LVT U836 ( .A1(n977), .A2(n978), .Y(n681) );
  AO21X1_LVT U837 ( .A1(n753), .A2(n681), .A3(n680), .Y(N285) );
  AO222X1_LVT U838 ( .A1(n783), .A2(n_T_65[71]), .A3(n931), .A4(n_T_51[126]), 
        .A5(subtractor[63]), .A6(n226), .Y(N523) );
  AO22X1_LVT U839 ( .A1(n157), .A2(n171), .A3(n805), .A4(n204), .Y(N294) );
  AND4X1_LVT U840 ( .A1(n272), .A2(n275), .A3(n274), .A4(n273), .Y(n777) );
  NAND4X0_LVT U841 ( .A1(n277), .A2(n278), .A3(n152), .A4(n183), .Y(n973) );
  AND4X1_LVT U842 ( .A1(n181), .A2(n264), .A3(n263), .A4(n266), .Y(n776) );
  AND4X1_LVT U843 ( .A1(n267), .A2(n270), .A3(n269), .A4(n268), .Y(n682) );
  AND2X1_LVT U844 ( .A1(n776), .A2(n682), .Y(n775) );
  AND4X1_LVT U845 ( .A1(n187), .A2(n149), .A3(n228), .A4(n229), .Y(n774) );
  AND4X1_LVT U846 ( .A1(n231), .A2(n234), .A3(n233), .A4(n232), .Y(n683) );
  NAND4X0_LVT U847 ( .A1(n259), .A2(n258), .A3(n261), .A4(n260), .Y(n970) );
  AND4X1_LVT U848 ( .A1(n188), .A2(n251), .A3(n250), .A4(n252), .Y(n772) );
  AND4X1_LVT U849 ( .A1(n248), .A2(n246), .A3(n249), .A4(n247), .Y(n771) );
  NAND2X0_LVT U850 ( .A1(n772), .A2(n771), .Y(n999) );
  NAND4X0_LVT U851 ( .A1(n254), .A2(n257), .A3(n256), .A4(n255), .Y(n971) );
  NOR2X0_LVT U852 ( .A1(divisor[57]), .A2(divisor[56]), .Y(n684) );
  NOR4X1_LVT U853 ( .A1(divisor[62]), .A2(divisor[61]), .A3(divisor[63]), .A4(
        divisor[60]), .Y(n769) );
  NAND4X0_LVT U854 ( .A1(n684), .A2(n769), .A3(n179), .A4(n180), .Y(n967) );
  NOR4X1_LVT U855 ( .A1(divisor[55]), .A2(divisor[54]), .A3(divisor[53]), .A4(
        divisor[52]), .Y(n770) );
  AND2X1_LVT U856 ( .A1(n216), .A2(n770), .Y(n717) );
  NOR4X1_LVT U857 ( .A1(divisor[51]), .A2(divisor[50]), .A3(divisor[49]), .A4(
        divisor[48]), .Y(n685) );
  NAND2X0_LVT U858 ( .A1(n717), .A2(n685), .Y(n956) );
  NOR4X1_LVT U859 ( .A1(divisor[46]), .A2(divisor[45]), .A3(divisor[47]), .A4(
        divisor[44]), .Y(n767) );
  NAND4X0_LVT U860 ( .A1(n686), .A2(n767), .A3(n185), .A4(n163), .Y(n966) );
  NOR4X1_LVT U861 ( .A1(divisor[38]), .A2(divisor[37]), .A3(divisor[39]), .A4(
        divisor[36]), .Y(n768) );
  AND2X1_LVT U862 ( .A1(n768), .A2(n723), .Y(n766) );
  NOR4X1_LVT U863 ( .A1(divisor[35]), .A2(divisor[34]), .A3(divisor[33]), .A4(
        divisor[32]), .Y(n932) );
  NOR4X1_LVT U864 ( .A1(divisor[31]), .A2(divisor[30]), .A3(divisor[29]), .A4(
        divisor[28]), .Y(n764) );
  NAND4X0_LVT U865 ( .A1(n687), .A2(n764), .A3(n196), .A4(n164), .Y(n964) );
  NOR4X1_LVT U866 ( .A1(divisor[22]), .A2(divisor[20]), .A3(divisor[23]), .A4(
        divisor[21]), .Y(n765) );
  INVX1_LVT U867 ( .A(n964), .Y(n728) );
  AND2X1_LVT U868 ( .A1(n765), .A2(n728), .Y(n727) );
  NOR4X1_LVT U869 ( .A1(divisor[18]), .A2(divisor[19]), .A3(divisor[17]), .A4(
        divisor[16]), .Y(n688) );
  AND2X1_LVT U870 ( .A1(n727), .A2(n688), .Y(n940) );
  NAND3X0_LVT U871 ( .A1(n727), .A2(divisor[17]), .A3(n161), .Y(n692) );
  NAND3X0_LVT U872 ( .A1(divisor[21]), .A2(n728), .A3(n190), .Y(n691) );
  NAND3X0_LVT U873 ( .A1(n764), .A2(divisor[25]), .A3(n196), .Y(n690) );
  NAND2X0_LVT U874 ( .A1(divisor[29]), .A2(n174), .Y(n689) );
  AND4X1_LVT U875 ( .A1(n692), .A2(n691), .A3(n690), .A4(n689), .Y(n694) );
  NAND3X0_LVT U876 ( .A1(n717), .A2(divisor[49]), .A3(n159), .Y(n693) );
  OA21X1_LVT U877 ( .A1(n694), .A2(n968), .A3(n693), .Y(n936) );
  NAND3X0_LVT U878 ( .A1(n216), .A2(divisor[53]), .A3(n195), .Y(n935) );
  NAND3X0_LVT U879 ( .A1(n769), .A2(divisor[57]), .A3(n179), .Y(n934) );
  NAND2X0_LVT U880 ( .A1(divisor[61]), .A2(n177), .Y(n933) );
  NAND2X0_LVT U881 ( .A1(n766), .A2(divisor[35]), .Y(n697) );
  NAND2X0_LVT U882 ( .A1(divisor[39]), .A2(n723), .Y(n696) );
  NAND2X0_LVT U883 ( .A1(n767), .A2(divisor[43]), .Y(n695) );
  AND4X1_LVT U884 ( .A1(n178), .A2(n697), .A3(n696), .A4(n695), .Y(n762) );
  NAND2X0_LVT U885 ( .A1(divisor[41]), .A2(n185), .Y(n698) );
  INVX1_LVT U886 ( .A(n767), .Y(n722) );
  OA22X1_LVT U887 ( .A1(divisor[46]), .A2(n173), .A3(n698), .A4(n722), .Y(n939) );
  NAND3X0_LVT U888 ( .A1(divisor[37]), .A2(n723), .A3(n192), .Y(n938) );
  NAND3X0_LVT U889 ( .A1(n766), .A2(divisor[33]), .A3(n160), .Y(n937) );
  NOR4X1_LVT U890 ( .A1(divisor[14]), .A2(divisor[13]), .A3(divisor[15]), .A4(
        divisor[12]), .Y(n761) );
  NAND4X0_LVT U891 ( .A1(n699), .A2(n761), .A3(n202), .A4(n165), .Y(n962) );
  NOR4X1_LVT U892 ( .A1(divisor[6]), .A2(divisor[7]), .A3(divisor[5]), .A4(
        divisor[4]), .Y(n760) );
  INVX1_LVT U893 ( .A(n962), .Y(n714) );
  AND2X1_LVT U894 ( .A1(n760), .A2(n714), .Y(n713) );
  NAND2X0_LVT U895 ( .A1(n713), .A2(divisor[3]), .Y(n702) );
  NAND2X0_LVT U896 ( .A1(divisor[7]), .A2(n714), .Y(n701) );
  NAND2X0_LVT U897 ( .A1(n761), .A2(divisor[11]), .Y(n700) );
  AND4X1_LVT U898 ( .A1(n162), .A2(n702), .A3(n701), .A4(n700), .Y(n759) );
  NAND2X0_LVT U899 ( .A1(divisor[9]), .A2(n202), .Y(n703) );
  INVX1_LVT U900 ( .A(n761), .Y(n715) );
  OA22X1_LVT U901 ( .A1(divisor[14]), .A2(n172), .A3(n703), .A4(n715), .Y(n943) );
  NAND3X0_LVT U902 ( .A1(divisor[5]), .A2(n714), .A3(n191), .Y(n942) );
  NAND3X0_LVT U903 ( .A1(n713), .A2(n205), .A3(divisor[1]), .Y(n941) );
  NAND2X0_LVT U904 ( .A1(n727), .A2(divisor[19]), .Y(n706) );
  NAND2X0_LVT U905 ( .A1(divisor[23]), .A2(n728), .Y(n705) );
  NAND2X0_LVT U906 ( .A1(n764), .A2(divisor[27]), .Y(n704) );
  NAND4X0_LVT U907 ( .A1(n176), .A2(n706), .A3(n705), .A4(n704), .Y(n711) );
  NAND2X0_LVT U908 ( .A1(divisor[51]), .A2(n717), .Y(n709) );
  NAND2X0_LVT U909 ( .A1(n216), .A2(divisor[55]), .Y(n708) );
  NAND2X0_LVT U910 ( .A1(n769), .A2(divisor[59]), .Y(n707) );
  NAND4X0_LVT U911 ( .A1(n175), .A2(n709), .A3(n708), .A4(n707), .Y(n710) );
  AO21X1_LVT U912 ( .A1(n763), .A2(n711), .A3(n710), .Y(n955) );
  INVX1_LVT U913 ( .A(n205), .Y(n712) );
  AO22X1_LVT U914 ( .A1(divisor[6]), .A2(n714), .A3(n713), .A4(n712), .Y(n950)
         );
  OR2X1_LVT U915 ( .A1(n202), .A2(n715), .Y(n716) );
  NAND3X0_LVT U916 ( .A1(n759), .A2(n193), .A3(n716), .Y(n949) );
  NAND2X0_LVT U917 ( .A1(n717), .A2(divisor[50]), .Y(n721) );
  NAND2X0_LVT U918 ( .A1(n216), .A2(divisor[54]), .Y(n720) );
  INVX1_LVT U919 ( .A(n179), .Y(n718) );
  NAND2X0_LVT U920 ( .A1(n769), .A2(n718), .Y(n719) );
  NAND4X0_LVT U921 ( .A1(n177), .A2(n721), .A3(n720), .A4(n719), .Y(n948) );
  OA21X1_LVT U922 ( .A1(n185), .A2(n722), .A3(n194), .Y(n726) );
  NAND2X0_LVT U923 ( .A1(divisor[38]), .A2(n723), .Y(n725) );
  NAND2X0_LVT U924 ( .A1(n766), .A2(divisor[34]), .Y(n724) );
  NAND4X0_LVT U925 ( .A1(n762), .A2(n726), .A3(n725), .A4(n724), .Y(n952) );
  NAND2X0_LVT U926 ( .A1(n727), .A2(divisor[18]), .Y(n731) );
  NAND2X0_LVT U927 ( .A1(divisor[22]), .A2(n728), .Y(n730) );
  NAND2X0_LVT U928 ( .A1(n764), .A2(divisor[26]), .Y(n729) );
  NAND4X0_LVT U929 ( .A1(n174), .A2(n731), .A3(n730), .A4(n729), .Y(n951) );
  AND2X1_LVT U930 ( .A1(n773), .A2(n779), .Y(n747) );
  AND2X1_LVT U931 ( .A1(n747), .A2(n732), .Y(n1002) );
  OR2X1_LVT U932 ( .A1(n971), .A2(n999), .Y(n998) );
  NAND2X0_LVT U933 ( .A1(n232), .A2(n_T_51[57]), .Y(n733) );
  INVX1_LVT U934 ( .A(n774), .Y(n746) );
  OA22X1_LVT U935 ( .A1(n229), .A2(n_T_51[62]), .A3(n733), .A4(n746), .Y(n983)
         );
  NAND3X0_LVT U936 ( .A1(n237), .A2(n773), .A3(n_T_51[53]), .Y(n982) );
  NAND3X0_LVT U937 ( .A1(n241), .A2(n_T_51[49]), .A3(n747), .Y(n981) );
  NAND2X0_LVT U938 ( .A1(n744), .A2(n_T_51[7]), .Y(n736) );
  NAND2X0_LVT U939 ( .A1(n305), .A2(n745), .Y(n735) );
  NAND2X0_LVT U940 ( .A1(n780), .A2(n_T_51[11]), .Y(n734) );
  AND4X1_LVT U941 ( .A1(n281), .A2(n736), .A3(n735), .A4(n734), .Y(n757) );
  INVX1_LVT U942 ( .A(n780), .Y(n743) );
  NAND2X0_LVT U943 ( .A1(n286), .A2(n_T_51[9]), .Y(n737) );
  OA22X1_LVT U944 ( .A1(n283), .A2(n_T_51[14]), .A3(n743), .A4(n737), .Y(n986)
         );
  NAND3X0_LVT U945 ( .A1(n291), .A2(n744), .A3(n_T_51[5]), .Y(n985) );
  NAND3X0_LVT U946 ( .A1(n745), .A2(n_T_51[1]), .A3(n208), .Y(n984) );
  INVX1_LVT U947 ( .A(n999), .Y(n741) );
  INVX1_LVT U948 ( .A(n998), .Y(n742) );
  NAND2X0_LVT U949 ( .A1(n251), .A2(n_T_51[41]), .Y(n738) );
  INVX1_LVT U950 ( .A(n771), .Y(n740) );
  OA22X1_LVT U951 ( .A1(n248), .A2(n_T_51[46]), .A3(n738), .A4(n740), .Y(n989)
         );
  NAND3X0_LVT U952 ( .A1(n255), .A2(n741), .A3(n_T_51[37]), .Y(n988) );
  NAND3X0_LVT U953 ( .A1(n742), .A2(n259), .A3(n_T_51[33]), .Y(n987) );
  AND2X1_LVT U954 ( .A1(n777), .A2(n775), .Y(n749) );
  INVX1_LVT U955 ( .A(n776), .Y(n748) );
  NAND2X0_LVT U956 ( .A1(n268), .A2(n_T_51[25]), .Y(n739) );
  OA22X1_LVT U957 ( .A1(n181), .A2(n_T_51[30]), .A3(n748), .A4(n739), .Y(n993)
         );
  NAND3X0_LVT U958 ( .A1(n273), .A2(n775), .A3(n_T_51[21]), .Y(n992) );
  NAND3X0_LVT U959 ( .A1(n749), .A2(n277), .A3(n_T_51[17]), .Y(n991) );
  INVX1_LVT U960 ( .A(n750), .Y(n751) );
  NAND2X0_LVT U961 ( .A1(n751), .A2(n199), .Y(N293) );
  NAND3X0_LVT U962 ( .A1(n753), .A2(n752), .A3(n203), .Y(N282) );
  AO21X1_LVT U963 ( .A1(n754), .A2(divisor[63]), .A3(n235), .Y(N322) );
  NAND3X0_LVT U964 ( .A1(n_T_69[6]), .A2(n_T_69[7]), .A3(n778), .Y(n804) );
  AND4X1_LVT U967 ( .A1(n_T_434[3]), .A2(n_T_434[5]), .A3(n_T_434[4]), .A4(
        n_T_434[0]), .Y(n791) );
  NAND3X0_LVT U968 ( .A1(n_T_434[2]), .A2(n_T_434[1]), .A3(n791), .Y(n792) );
  NAND2X0_LVT U969 ( .A1(n230), .A2(n200), .Y(n805) );
  AO22X1_LVT U970 ( .A1(n_T_85[4]), .A2(n805), .A3(n157), .A4(n166), .Y(N295)
         );
  NAND2X0_LVT U971 ( .A1(n225), .A2(n167), .Y(n799) );
  NAND3X0_LVT U972 ( .A1(n235), .A2(n787), .A3(n784), .Y(n797) );
  NAND3X0_LVT U973 ( .A1(n799), .A2(n798), .A3(n797), .Y(N296) );
  AO22X1_LVT U974 ( .A1(n_T_69[6]), .A2(n800), .A3(n198), .A4(n778), .Y(n801)
         );
  AO22X1_LVT U975 ( .A1(n801), .A2(n805), .A3(n225), .A4(n168), .Y(N297) );
  OA221X1_LVT U976 ( .A1(n_T_69[7]), .A2(n_T_69[6]), .A3(n_T_69[7]), .A4(n778), 
        .A5(n804), .Y(n802) );
  AO22X1_LVT U977 ( .A1(n802), .A2(n805), .A3(n225), .A4(n169), .Y(N298) );
  AO22X1_LVT U978 ( .A1(n_T_69[8]), .A2(n804), .A3(n197), .A4(n803), .Y(n806)
         );
  AO22X1_LVT U979 ( .A1(n806), .A2(n805), .A3(n225), .A4(n170), .Y(N299) );
  AO22X1_LVT U980 ( .A1(n225), .A2(n_T_442[65]), .A3(n931), .A4(n301), .Y(n808) );
  AO22X1_LVT U981 ( .A1(n783), .A2(n_T_65[8]), .A3(n226), .A4(subtractor[0]), 
        .Y(n807) );
  OR2X1_LVT U982 ( .A1(n808), .A2(n807), .Y(N459) );
  AO22X1_LVT U983 ( .A1(n157), .A2(n_T_442[66]), .A3(n_T_51[64]), .A4(n931), 
        .Y(n810) );
  AO22X1_LVT U984 ( .A1(n783), .A2(n_T_65[9]), .A3(n226), .A4(subtractor[1]), 
        .Y(n809) );
  OR2X1_LVT U985 ( .A1(n810), .A2(n809), .Y(N460) );
  AO22X1_LVT U986 ( .A1(n225), .A2(n_T_442[67]), .A3(n931), .A4(n_T_51[65]), 
        .Y(n812) );
  AO22X1_LVT U987 ( .A1(n783), .A2(n_T_65[10]), .A3(n226), .A4(subtractor[2]), 
        .Y(n811) );
  OR2X1_LVT U988 ( .A1(n812), .A2(n811), .Y(N461) );
  AO22X1_LVT U989 ( .A1(n225), .A2(n_T_442[68]), .A3(n931), .A4(n_T_51[66]), 
        .Y(n814) );
  AO22X1_LVT U990 ( .A1(n783), .A2(n_T_65[11]), .A3(n226), .A4(subtractor[3]), 
        .Y(n813) );
  OR2X1_LVT U991 ( .A1(n814), .A2(n813), .Y(N462) );
  AO22X1_LVT U992 ( .A1(n225), .A2(n_T_442[69]), .A3(n931), .A4(n_T_51[67]), 
        .Y(n816) );
  AO22X1_LVT U993 ( .A1(n783), .A2(n_T_65[12]), .A3(n226), .A4(subtractor[4]), 
        .Y(n815) );
  OR2X1_LVT U994 ( .A1(n816), .A2(n815), .Y(N463) );
  AO22X1_LVT U995 ( .A1(n225), .A2(n_T_442[70]), .A3(n931), .A4(n_T_51[68]), 
        .Y(n818) );
  AO22X1_LVT U996 ( .A1(n783), .A2(n_T_65[13]), .A3(n226), .A4(subtractor[5]), 
        .Y(n817) );
  OR2X1_LVT U997 ( .A1(n818), .A2(n817), .Y(N464) );
  AO22X1_LVT U998 ( .A1(n225), .A2(n_T_442[71]), .A3(n931), .A4(n_T_51[69]), 
        .Y(n820) );
  AO22X1_LVT U999 ( .A1(n783), .A2(n_T_65[14]), .A3(n226), .A4(subtractor[6]), 
        .Y(n819) );
  OR2X1_LVT U1000 ( .A1(n820), .A2(n819), .Y(N465) );
  AO22X1_LVT U1001 ( .A1(n225), .A2(n_T_442[72]), .A3(n931), .A4(n_T_51[70]), 
        .Y(n822) );
  AO22X1_LVT U1002 ( .A1(n783), .A2(n_T_65[15]), .A3(n226), .A4(subtractor[7]), 
        .Y(n821) );
  OR2X1_LVT U1003 ( .A1(n822), .A2(n821), .Y(N466) );
  AO22X1_LVT U1004 ( .A1(n225), .A2(n_T_442[73]), .A3(n931), .A4(n_T_51[71]), 
        .Y(n824) );
  AO22X1_LVT U1005 ( .A1(n783), .A2(n_T_65[16]), .A3(n226), .A4(subtractor[8]), 
        .Y(n823) );
  OR2X1_LVT U1006 ( .A1(n824), .A2(n823), .Y(N467) );
  AO22X1_LVT U1007 ( .A1(n157), .A2(n_T_442[74]), .A3(n931), .A4(n_T_51[72]), 
        .Y(n826) );
  AO22X1_LVT U1008 ( .A1(n783), .A2(n_T_65[17]), .A3(n226), .A4(subtractor[9]), 
        .Y(n825) );
  OR2X1_LVT U1009 ( .A1(n826), .A2(n825), .Y(N468) );
  AO22X1_LVT U1010 ( .A1(n225), .A2(n_T_442[75]), .A3(n931), .A4(n_T_51[73]), 
        .Y(n828) );
  AO22X1_LVT U1011 ( .A1(n783), .A2(n_T_65[18]), .A3(n226), .A4(subtractor[10]), .Y(n827) );
  OR2X1_LVT U1012 ( .A1(n828), .A2(n827), .Y(N469) );
  AO22X1_LVT U1013 ( .A1(n225), .A2(n_T_442[76]), .A3(n931), .A4(n_T_51[74]), 
        .Y(n830) );
  AO22X1_LVT U1014 ( .A1(n783), .A2(n_T_65[19]), .A3(n226), .A4(subtractor[11]), .Y(n829) );
  OR2X1_LVT U1015 ( .A1(n830), .A2(n829), .Y(N470) );
  AO22X1_LVT U1016 ( .A1(n225), .A2(n_T_442[77]), .A3(n931), .A4(n_T_51[75]), 
        .Y(n832) );
  AO22X1_LVT U1017 ( .A1(n783), .A2(n_T_65[20]), .A3(n226), .A4(subtractor[12]), .Y(n831) );
  OR2X1_LVT U1018 ( .A1(n832), .A2(n831), .Y(N471) );
  AO22X1_LVT U1019 ( .A1(n225), .A2(n_T_442[78]), .A3(n931), .A4(n_T_51[76]), 
        .Y(n834) );
  AO22X1_LVT U1020 ( .A1(n783), .A2(n_T_65[21]), .A3(n226), .A4(subtractor[13]), .Y(n833) );
  OR2X1_LVT U1021 ( .A1(n834), .A2(n833), .Y(N472) );
  AO22X1_LVT U1022 ( .A1(n157), .A2(n_T_442[79]), .A3(n931), .A4(n_T_51[77]), 
        .Y(n836) );
  AO22X1_LVT U1023 ( .A1(n783), .A2(n_T_65[22]), .A3(n226), .A4(subtractor[14]), .Y(n835) );
  OR2X1_LVT U1024 ( .A1(n836), .A2(n835), .Y(N473) );
  AO22X1_LVT U1025 ( .A1(n225), .A2(n_T_442[80]), .A3(n931), .A4(n_T_51[78]), 
        .Y(n838) );
  AO22X1_LVT U1026 ( .A1(n783), .A2(n_T_65[23]), .A3(n226), .A4(subtractor[15]), .Y(n837) );
  OR2X1_LVT U1027 ( .A1(n838), .A2(n837), .Y(N474) );
  AO22X1_LVT U1028 ( .A1(n225), .A2(n_T_442[81]), .A3(n931), .A4(n_T_51[79]), 
        .Y(n840) );
  AO22X1_LVT U1029 ( .A1(n783), .A2(n_T_65[24]), .A3(n226), .A4(subtractor[16]), .Y(n839) );
  OR2X1_LVT U1030 ( .A1(n840), .A2(n839), .Y(N475) );
  AO22X1_LVT U1031 ( .A1(n225), .A2(n_T_442[82]), .A3(n931), .A4(n_T_51[80]), 
        .Y(n842) );
  AO22X1_LVT U1032 ( .A1(n783), .A2(n_T_65[25]), .A3(n226), .A4(subtractor[17]), .Y(n841) );
  OR2X1_LVT U1033 ( .A1(n842), .A2(n841), .Y(N476) );
  AO22X1_LVT U1034 ( .A1(n225), .A2(n_T_442[83]), .A3(n931), .A4(n_T_51[81]), 
        .Y(n844) );
  AO22X1_LVT U1035 ( .A1(n783), .A2(n_T_65[26]), .A3(n226), .A4(subtractor[18]), .Y(n843) );
  OR2X1_LVT U1036 ( .A1(n844), .A2(n843), .Y(N477) );
  AO22X1_LVT U1037 ( .A1(n225), .A2(n_T_442[84]), .A3(n931), .A4(n_T_51[82]), 
        .Y(n846) );
  AO22X1_LVT U1038 ( .A1(n783), .A2(n_T_65[27]), .A3(n226), .A4(subtractor[19]), .Y(n845) );
  OR2X1_LVT U1039 ( .A1(n846), .A2(n845), .Y(N478) );
  AO22X1_LVT U1040 ( .A1(n225), .A2(n_T_442[85]), .A3(n931), .A4(n_T_51[83]), 
        .Y(n848) );
  AO22X1_LVT U1041 ( .A1(n783), .A2(n_T_65[28]), .A3(n226), .A4(subtractor[20]), .Y(n847) );
  OR2X1_LVT U1042 ( .A1(n848), .A2(n847), .Y(N479) );
  AO22X1_LVT U1043 ( .A1(n225), .A2(n_T_442[86]), .A3(n931), .A4(n_T_51[84]), 
        .Y(n850) );
  AO22X1_LVT U1044 ( .A1(n783), .A2(n_T_65[29]), .A3(n226), .A4(subtractor[21]), .Y(n849) );
  OR2X1_LVT U1045 ( .A1(n850), .A2(n849), .Y(N480) );
  AO22X1_LVT U1046 ( .A1(n225), .A2(n_T_442[87]), .A3(n931), .A4(n_T_51[85]), 
        .Y(n852) );
  AO22X1_LVT U1047 ( .A1(n783), .A2(n_T_65[30]), .A3(n226), .A4(subtractor[22]), .Y(n851) );
  OR2X1_LVT U1048 ( .A1(n852), .A2(n851), .Y(N481) );
  AO22X1_LVT U1049 ( .A1(n157), .A2(n_T_442[88]), .A3(n931), .A4(n_T_51[86]), 
        .Y(n854) );
  AO22X1_LVT U1050 ( .A1(n783), .A2(n_T_65[31]), .A3(n226), .A4(subtractor[23]), .Y(n853) );
  OR2X1_LVT U1051 ( .A1(n854), .A2(n853), .Y(N482) );
  AO22X1_LVT U1052 ( .A1(n225), .A2(n_T_442[89]), .A3(n931), .A4(n_T_51[87]), 
        .Y(n856) );
  AO22X1_LVT U1053 ( .A1(n783), .A2(n_T_65[32]), .A3(n226), .A4(subtractor[24]), .Y(n855) );
  OR2X1_LVT U1054 ( .A1(n856), .A2(n855), .Y(N483) );
  AO22X1_LVT U1055 ( .A1(n157), .A2(n_T_442[90]), .A3(n931), .A4(n_T_51[88]), 
        .Y(n858) );
  AO22X1_LVT U1056 ( .A1(n783), .A2(n_T_65[33]), .A3(n226), .A4(subtractor[25]), .Y(n857) );
  OR2X1_LVT U1057 ( .A1(n858), .A2(n857), .Y(N484) );
  AO22X1_LVT U1058 ( .A1(n225), .A2(n_T_442[91]), .A3(n931), .A4(n_T_51[89]), 
        .Y(n860) );
  AO22X1_LVT U1059 ( .A1(n783), .A2(n_T_65[34]), .A3(n226), .A4(subtractor[26]), .Y(n859) );
  OR2X1_LVT U1060 ( .A1(n860), .A2(n859), .Y(N485) );
  AO22X1_LVT U1061 ( .A1(n225), .A2(n_T_442[92]), .A3(n931), .A4(n_T_51[90]), 
        .Y(n862) );
  AO22X1_LVT U1062 ( .A1(n783), .A2(n_T_65[35]), .A3(n226), .A4(subtractor[27]), .Y(n861) );
  OR2X1_LVT U1063 ( .A1(n862), .A2(n861), .Y(N486) );
  AO22X1_LVT U1064 ( .A1(n157), .A2(n_T_442[93]), .A3(n931), .A4(n_T_51[91]), 
        .Y(n864) );
  AO22X1_LVT U1065 ( .A1(n783), .A2(n_T_65[36]), .A3(n226), .A4(subtractor[28]), .Y(n863) );
  OR2X1_LVT U1066 ( .A1(n864), .A2(n863), .Y(N487) );
  AO22X1_LVT U1067 ( .A1(n225), .A2(n_T_442[94]), .A3(n931), .A4(n_T_51[92]), 
        .Y(n866) );
  AO22X1_LVT U1068 ( .A1(n783), .A2(n_T_65[37]), .A3(n226), .A4(subtractor[29]), .Y(n865) );
  OR2X1_LVT U1069 ( .A1(n866), .A2(n865), .Y(N488) );
  AO22X1_LVT U1070 ( .A1(n225), .A2(n_T_442[95]), .A3(n931), .A4(n_T_51[93]), 
        .Y(n868) );
  AO22X1_LVT U1071 ( .A1(n783), .A2(n_T_65[38]), .A3(n226), .A4(subtractor[30]), .Y(n867) );
  OR2X1_LVT U1072 ( .A1(n868), .A2(n867), .Y(N489) );
  AO22X1_LVT U1073 ( .A1(n157), .A2(n_T_442[96]), .A3(n931), .A4(n_T_51[94]), 
        .Y(n870) );
  AO22X1_LVT U1074 ( .A1(n783), .A2(n_T_65[39]), .A3(n226), .A4(subtractor[31]), .Y(n869) );
  OR2X1_LVT U1075 ( .A1(n870), .A2(n869), .Y(N490) );
  AO22X1_LVT U1076 ( .A1(n225), .A2(n_T_442[97]), .A3(n931), .A4(n_T_51[95]), 
        .Y(n872) );
  AO22X1_LVT U1077 ( .A1(n783), .A2(n_T_65[40]), .A3(n226), .A4(subtractor[32]), .Y(n871) );
  OR2X1_LVT U1078 ( .A1(n872), .A2(n871), .Y(N491) );
  AO22X1_LVT U1079 ( .A1(n225), .A2(n_T_442[98]), .A3(n931), .A4(n_T_51[96]), 
        .Y(n874) );
  AO22X1_LVT U1080 ( .A1(n783), .A2(n_T_65[41]), .A3(n226), .A4(subtractor[33]), .Y(n873) );
  OR2X1_LVT U1081 ( .A1(n874), .A2(n873), .Y(N492) );
  AO22X1_LVT U1082 ( .A1(n157), .A2(n_T_442[99]), .A3(n931), .A4(n_T_51[97]), 
        .Y(n876) );
  AO22X1_LVT U1083 ( .A1(n783), .A2(n_T_65[42]), .A3(n226), .A4(subtractor[34]), .Y(n875) );
  OR2X1_LVT U1084 ( .A1(n876), .A2(n875), .Y(N494) );
  AO22X1_LVT U1085 ( .A1(n225), .A2(n_T_442[100]), .A3(n931), .A4(n_T_51[98]), 
        .Y(n878) );
  AO22X1_LVT U1086 ( .A1(n783), .A2(n_T_65[43]), .A3(n226), .A4(subtractor[35]), .Y(n877) );
  OR2X1_LVT U1087 ( .A1(n878), .A2(n877), .Y(N495) );
  AO22X1_LVT U1088 ( .A1(n225), .A2(n_T_442[101]), .A3(n931), .A4(n_T_51[99]), 
        .Y(n880) );
  AO22X1_LVT U1089 ( .A1(n783), .A2(n_T_65[44]), .A3(n226), .A4(subtractor[36]), .Y(n879) );
  OR2X1_LVT U1090 ( .A1(n880), .A2(n879), .Y(N496) );
  AO22X1_LVT U1091 ( .A1(n157), .A2(n_T_442[102]), .A3(n931), .A4(n_T_51[100]), 
        .Y(n882) );
  AO22X1_LVT U1092 ( .A1(n783), .A2(n_T_65[45]), .A3(n226), .A4(subtractor[37]), .Y(n881) );
  OR2X1_LVT U1093 ( .A1(n882), .A2(n881), .Y(N497) );
  AO22X1_LVT U1094 ( .A1(n225), .A2(n_T_442[103]), .A3(n931), .A4(n_T_51[101]), 
        .Y(n884) );
  AO22X1_LVT U1095 ( .A1(n783), .A2(n_T_65[46]), .A3(n226), .A4(subtractor[38]), .Y(n883) );
  OR2X1_LVT U1096 ( .A1(n884), .A2(n883), .Y(N498) );
  AO22X1_LVT U1097 ( .A1(n225), .A2(n_T_442[104]), .A3(n931), .A4(n_T_51[102]), 
        .Y(n886) );
  AO22X1_LVT U1098 ( .A1(n783), .A2(n_T_65[47]), .A3(n226), .A4(subtractor[39]), .Y(n885) );
  OR2X1_LVT U1099 ( .A1(n886), .A2(n885), .Y(N499) );
  AO22X1_LVT U1100 ( .A1(n225), .A2(n_T_442[105]), .A3(n931), .A4(n_T_51[103]), 
        .Y(n888) );
  AO22X1_LVT U1101 ( .A1(n783), .A2(n_T_65[48]), .A3(n226), .A4(subtractor[40]), .Y(n887) );
  OR2X1_LVT U1102 ( .A1(n888), .A2(n887), .Y(N500) );
  AO22X1_LVT U1103 ( .A1(n225), .A2(n_T_442[106]), .A3(n931), .A4(n_T_51[104]), 
        .Y(n890) );
  AO22X1_LVT U1104 ( .A1(n783), .A2(n_T_65[49]), .A3(n226), .A4(subtractor[41]), .Y(n889) );
  OR2X1_LVT U1105 ( .A1(n890), .A2(n889), .Y(N501) );
  AO22X1_LVT U1106 ( .A1(n157), .A2(n_T_442[107]), .A3(n931), .A4(n_T_51[105]), 
        .Y(n892) );
  AO22X1_LVT U1107 ( .A1(n783), .A2(n_T_65[50]), .A3(n226), .A4(subtractor[42]), .Y(n891) );
  OR2X1_LVT U1108 ( .A1(n892), .A2(n891), .Y(N502) );
  AO22X1_LVT U1109 ( .A1(n225), .A2(n_T_442[108]), .A3(n931), .A4(n_T_51[106]), 
        .Y(n894) );
  AO22X1_LVT U1110 ( .A1(n783), .A2(n_T_65[51]), .A3(n226), .A4(subtractor[43]), .Y(n893) );
  OR2X1_LVT U1111 ( .A1(n894), .A2(n893), .Y(N503) );
  AO22X1_LVT U1112 ( .A1(n225), .A2(n_T_442[109]), .A3(n931), .A4(n_T_51[107]), 
        .Y(n896) );
  AO22X1_LVT U1113 ( .A1(n783), .A2(n_T_65[52]), .A3(n226), .A4(subtractor[44]), .Y(n895) );
  OR2X1_LVT U1114 ( .A1(n896), .A2(n895), .Y(N504) );
  AO22X1_LVT U1115 ( .A1(n225), .A2(n_T_442[110]), .A3(n931), .A4(n_T_51[108]), 
        .Y(n898) );
  AO22X1_LVT U1116 ( .A1(n783), .A2(n_T_65[53]), .A3(n226), .A4(subtractor[45]), .Y(n897) );
  OR2X1_LVT U1117 ( .A1(n898), .A2(n897), .Y(N505) );
  AO22X1_LVT U1118 ( .A1(n157), .A2(n_T_442[111]), .A3(n931), .A4(n_T_51[109]), 
        .Y(n900) );
  AO22X1_LVT U1119 ( .A1(n783), .A2(n_T_65[54]), .A3(n226), .A4(subtractor[46]), .Y(n899) );
  OR2X1_LVT U1120 ( .A1(n900), .A2(n899), .Y(N506) );
  AO22X1_LVT U1121 ( .A1(n225), .A2(n_T_442[112]), .A3(n931), .A4(n_T_51[110]), 
        .Y(n902) );
  AO22X1_LVT U1122 ( .A1(n783), .A2(n_T_65[55]), .A3(n226), .A4(subtractor[47]), .Y(n901) );
  OR2X1_LVT U1123 ( .A1(n902), .A2(n901), .Y(N507) );
  AO22X1_LVT U1124 ( .A1(n225), .A2(n_T_442[113]), .A3(n931), .A4(n_T_51[111]), 
        .Y(n904) );
  AO22X1_LVT U1125 ( .A1(n783), .A2(n_T_65[56]), .A3(n226), .A4(subtractor[48]), .Y(n903) );
  OR2X1_LVT U1126 ( .A1(n904), .A2(n903), .Y(N508) );
  AO22X1_LVT U1127 ( .A1(n225), .A2(n_T_442[114]), .A3(n931), .A4(n_T_51[112]), 
        .Y(n906) );
  AO22X1_LVT U1128 ( .A1(n783), .A2(n_T_65[57]), .A3(n226), .A4(subtractor[49]), .Y(n905) );
  OR2X1_LVT U1129 ( .A1(n906), .A2(n905), .Y(N509) );
  AO22X1_LVT U1130 ( .A1(n225), .A2(n_T_442[115]), .A3(n931), .A4(n_T_51[113]), 
        .Y(n908) );
  AO22X1_LVT U1131 ( .A1(n783), .A2(n_T_65[58]), .A3(n226), .A4(subtractor[50]), .Y(n907) );
  OR2X1_LVT U1132 ( .A1(n908), .A2(n907), .Y(N510) );
  AO22X1_LVT U1133 ( .A1(n225), .A2(n_T_442[116]), .A3(n931), .A4(n_T_51[114]), 
        .Y(n910) );
  AO22X1_LVT U1134 ( .A1(n783), .A2(n_T_65[59]), .A3(n226), .A4(subtractor[51]), .Y(n909) );
  OR2X1_LVT U1135 ( .A1(n910), .A2(n909), .Y(N511) );
  AO22X1_LVT U1136 ( .A1(n225), .A2(n_T_442[117]), .A3(n931), .A4(n_T_51[115]), 
        .Y(n912) );
  AO22X1_LVT U1137 ( .A1(n783), .A2(n_T_65[60]), .A3(n226), .A4(subtractor[52]), .Y(n911) );
  OR2X1_LVT U1138 ( .A1(n912), .A2(n911), .Y(N512) );
  AO22X1_LVT U1139 ( .A1(n157), .A2(n_T_442[118]), .A3(n931), .A4(n_T_51[116]), 
        .Y(n914) );
  AO22X1_LVT U1140 ( .A1(n783), .A2(n_T_65[61]), .A3(n226), .A4(subtractor[53]), .Y(n913) );
  OR2X1_LVT U1141 ( .A1(n914), .A2(n913), .Y(N513) );
  AO22X1_LVT U1142 ( .A1(n225), .A2(n_T_442[119]), .A3(n931), .A4(n_T_51[117]), 
        .Y(n916) );
  AO22X1_LVT U1143 ( .A1(n783), .A2(n_T_65[62]), .A3(n226), .A4(subtractor[54]), .Y(n915) );
  OR2X1_LVT U1144 ( .A1(n916), .A2(n915), .Y(N514) );
  AO22X1_LVT U1145 ( .A1(n225), .A2(n_T_442[120]), .A3(n931), .A4(n_T_51[118]), 
        .Y(n918) );
  AO22X1_LVT U1146 ( .A1(n783), .A2(n_T_65[63]), .A3(n226), .A4(subtractor[55]), .Y(n917) );
  OR2X1_LVT U1147 ( .A1(n918), .A2(n917), .Y(N515) );
  AO22X1_LVT U1148 ( .A1(n225), .A2(n_T_442[121]), .A3(n931), .A4(n_T_51[119]), 
        .Y(n920) );
  AO22X1_LVT U1149 ( .A1(n783), .A2(n_T_65[64]), .A3(n226), .A4(subtractor[56]), .Y(n919) );
  OR2X1_LVT U1150 ( .A1(n920), .A2(n919), .Y(N516) );
  AO22X1_LVT U1151 ( .A1(n225), .A2(n_T_442[122]), .A3(n931), .A4(n_T_51[120]), 
        .Y(n922) );
  AO22X1_LVT U1152 ( .A1(n783), .A2(n_T_65[65]), .A3(n226), .A4(subtractor[57]), .Y(n921) );
  OR2X1_LVT U1153 ( .A1(n922), .A2(n921), .Y(N517) );
  AO22X1_LVT U1154 ( .A1(n157), .A2(n_T_442[123]), .A3(n931), .A4(n_T_51[121]), 
        .Y(n924) );
  AO22X1_LVT U1155 ( .A1(n783), .A2(n_T_65[66]), .A3(n226), .A4(subtractor[58]), .Y(n923) );
  OR2X1_LVT U1156 ( .A1(n924), .A2(n923), .Y(N518) );
  AO22X1_LVT U1157 ( .A1(n157), .A2(n_T_442[124]), .A3(n931), .A4(n_T_51[122]), 
        .Y(n926) );
  AO22X1_LVT U1158 ( .A1(n783), .A2(n_T_65[67]), .A3(n226), .A4(subtractor[59]), .Y(n925) );
  OR2X1_LVT U1159 ( .A1(n926), .A2(n925), .Y(N519) );
  AO22X1_LVT U1160 ( .A1(n157), .A2(n_T_442[125]), .A3(n931), .A4(n_T_51[123]), 
        .Y(n928) );
  AO22X1_LVT U1161 ( .A1(n783), .A2(n_T_65[68]), .A3(n226), .A4(subtractor[60]), .Y(n927) );
  OR2X1_LVT U1162 ( .A1(n928), .A2(n927), .Y(N520) );
  AO22X1_LVT U1163 ( .A1(n157), .A2(n_T_442[126]), .A3(n931), .A4(n_T_51[124]), 
        .Y(n930) );
  AO22X1_LVT U1164 ( .A1(n783), .A2(n_T_65[69]), .A3(n226), .A4(subtractor[61]), .Y(n929) );
  OR2X1_LVT U1165 ( .A1(n930), .A2(n929), .Y(N521) );
  NAND3X0_LVT U1166 ( .A1(n969), .A2(n766), .A3(n932), .Y(n_T_273_5_) );
  NAND4X0_LVT U1167 ( .A1(n936), .A2(n935), .A3(n934), .A4(n933), .Y(n947) );
  NAND4X0_LVT U1168 ( .A1(n762), .A2(n939), .A3(n938), .A4(n937), .Y(n945) );
  NAND2X0_LVT U1169 ( .A1(n965), .A2(n940), .Y(n957) );
  NAND4X0_LVT U1170 ( .A1(n759), .A2(n943), .A3(n942), .A4(n941), .Y(n944) );
  AO22X1_LVT U1171 ( .A1(n969), .A2(n945), .A3(n963), .A4(n944), .Y(n946) );
  OR3X1_LVT U1172 ( .A1(n955), .A2(n947), .A3(n946), .Y(n_T_272[0]) );
  AO221X1_LVT U1173 ( .A1(n963), .A2(n950), .A3(n963), .A4(n949), .A5(n948), 
        .Y(n954) );
  AO22X1_LVT U1174 ( .A1(n969), .A2(n952), .A3(n763), .A4(n951), .Y(n953) );
  OR3X1_LVT U1175 ( .A1(n955), .A2(n954), .A3(n953), .Y(n_T_272[1]) );
  OA21X1_LVT U1176 ( .A1(n770), .A2(n967), .A3(n769), .Y(n961) );
  AO221X1_LVT U1177 ( .A1(n764), .A2(n765), .A3(n764), .A4(n964), .A5(
        n_T_273_5_), .Y(n960) );
  AO221X1_LVT U1178 ( .A1(n767), .A2(n768), .A3(n767), .A4(n966), .A5(n956), 
        .Y(n959) );
  AO221X1_LVT U1179 ( .A1(n761), .A2(n760), .A3(n761), .A4(n962), .A5(n957), 
        .Y(n958) );
  NAND4X0_LVT U1180 ( .A1(n961), .A2(n960), .A3(n959), .A4(n958), .Y(
        n_T_272[2]) );
  NAND2X0_LVT U1181 ( .A1(n969), .A2(n968), .Y(n_T_272[4]) );
  OR3X1_LVT U1182 ( .A1(n974), .A2(n973), .A3(n997), .Y(n975) );
  NAND2X0_LVT U1183 ( .A1(n976), .A2(n975), .Y(n990) );
  NAND2X0_LVT U1184 ( .A1(n1002), .A2(n990), .Y(n_T_429[4]) );
  AO22X1_LVT U1185 ( .A1(n146), .A2(result[32]), .A3(n209), .A4(result[0]), 
        .Y(io_resp_bits_data[0]) );
  AO22X1_LVT U1186 ( .A1(n146), .A2(result[42]), .A3(n209), .A4(result[10]), 
        .Y(io_resp_bits_data[10]) );
  AO22X1_LVT U1187 ( .A1(n146), .A2(result[44]), .A3(n209), .A4(result[12]), 
        .Y(io_resp_bits_data[12]) );
  AO22X1_LVT U1188 ( .A1(n146), .A2(result[45]), .A3(n209), .A4(result[13]), 
        .Y(io_resp_bits_data[13]) );
  AO22X1_LVT U1189 ( .A1(n146), .A2(result[46]), .A3(n209), .A4(result[14]), 
        .Y(io_resp_bits_data[14]) );
  AO22X1_LVT U1190 ( .A1(n146), .A2(result[47]), .A3(n209), .A4(result[15]), 
        .Y(io_resp_bits_data[15]) );
  AO22X1_LVT U1191 ( .A1(n146), .A2(result[48]), .A3(n209), .A4(result[16]), 
        .Y(io_resp_bits_data[16]) );
  AO22X1_LVT U1192 ( .A1(n146), .A2(result[49]), .A3(n209), .A4(result[17]), 
        .Y(io_resp_bits_data[17]) );
  AO22X1_LVT U1193 ( .A1(n146), .A2(result[50]), .A3(n209), .A4(result[18]), 
        .Y(io_resp_bits_data[18]) );
  AO22X1_LVT U1194 ( .A1(n146), .A2(result[51]), .A3(n209), .A4(result[19]), 
        .Y(io_resp_bits_data[19]) );
  AO22X1_LVT U1195 ( .A1(n146), .A2(result[33]), .A3(n209), .A4(result[1]), 
        .Y(io_resp_bits_data[1]) );
  AO22X1_LVT U1196 ( .A1(n146), .A2(result[52]), .A3(n209), .A4(result[20]), 
        .Y(io_resp_bits_data[20]) );
  AO22X1_LVT U1197 ( .A1(n146), .A2(result[53]), .A3(n209), .A4(result[21]), 
        .Y(io_resp_bits_data[21]) );
  AO22X1_LVT U1198 ( .A1(n146), .A2(result[55]), .A3(n209), .A4(result[23]), 
        .Y(io_resp_bits_data[23]) );
  AO22X1_LVT U1199 ( .A1(n146), .A2(result[56]), .A3(n209), .A4(result[24]), 
        .Y(io_resp_bits_data[24]) );
  AO22X1_LVT U1200 ( .A1(n146), .A2(result[57]), .A3(n209), .A4(result[25]), 
        .Y(io_resp_bits_data[25]) );
  AO22X1_LVT U1201 ( .A1(n146), .A2(result[58]), .A3(n209), .A4(result[26]), 
        .Y(io_resp_bits_data[26]) );
  AO22X1_LVT U1202 ( .A1(n146), .A2(result[59]), .A3(n209), .A4(result[27]), 
        .Y(io_resp_bits_data[27]) );
  AO22X1_LVT U1203 ( .A1(n146), .A2(result[60]), .A3(n209), .A4(result[28]), 
        .Y(io_resp_bits_data[28]) );
  AO22X1_LVT U1204 ( .A1(n146), .A2(result[61]), .A3(n209), .A4(result[29]), 
        .Y(io_resp_bits_data[29]) );
  AO22X1_LVT U1205 ( .A1(n146), .A2(result[34]), .A3(n209), .A4(result[2]), 
        .Y(io_resp_bits_data[2]) );
  AO22X1_LVT U1206 ( .A1(n146), .A2(result[62]), .A3(n209), .A4(result[30]), 
        .Y(io_resp_bits_data[30]) );
  AO22X1_LVT U1207 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[32]), .Y(io_resp_bits_data[32]) );
  AO22X1_LVT U1208 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[33]), .Y(io_resp_bits_data[33]) );
  AO22X1_LVT U1209 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[34]), .Y(io_resp_bits_data[34]) );
  AO22X1_LVT U1210 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[35]), .Y(io_resp_bits_data[35]) );
  AO22X1_LVT U1211 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[36]), .Y(io_resp_bits_data[36]) );
  AO22X1_LVT U1212 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[37]), .Y(io_resp_bits_data[37]) );
  AO22X1_LVT U1213 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[38]), .Y(io_resp_bits_data[38]) );
  AO22X1_LVT U1214 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[39]), .Y(io_resp_bits_data[39]) );
  AO22X1_LVT U1215 ( .A1(n146), .A2(result[35]), .A3(n209), .A4(result[3]), 
        .Y(io_resp_bits_data[3]) );
  AO22X1_LVT U1216 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[40]), .Y(io_resp_bits_data[40]) );
  AO22X1_LVT U1217 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[41]), .Y(io_resp_bits_data[41]) );
  AO22X1_LVT U1218 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[42]), .Y(io_resp_bits_data[42]) );
  AO22X1_LVT U1219 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[43]), .Y(io_resp_bits_data[43]) );
  AO22X1_LVT U1220 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[44]), .Y(io_resp_bits_data[44]) );
  AO22X1_LVT U1221 ( .A1(n156), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[45]), .Y(io_resp_bits_data[45]) );
  AO22X1_LVT U1222 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[46]), .Y(io_resp_bits_data[46]) );
  AO22X1_LVT U1223 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[47]), .Y(io_resp_bits_data[47]) );
  AO22X1_LVT U1224 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[48]), .Y(io_resp_bits_data[48]) );
  AO22X1_LVT U1225 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[49]), .Y(io_resp_bits_data[49]) );
  AO22X1_LVT U1226 ( .A1(n146), .A2(result[36]), .A3(n209), .A4(result[4]), 
        .Y(io_resp_bits_data[4]) );
  AO22X1_LVT U1227 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[50]), .Y(io_resp_bits_data[50]) );
  AO22X1_LVT U1228 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[51]), .Y(io_resp_bits_data[51]) );
  AO22X1_LVT U1229 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[52]), .Y(io_resp_bits_data[52]) );
  AO22X1_LVT U1230 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[53]), .Y(io_resp_bits_data[53]) );
  AO22X1_LVT U1231 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[54]), .Y(io_resp_bits_data[54]) );
  AO22X1_LVT U1232 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n206), .A4(
        result[55]), .Y(io_resp_bits_data[55]) );
  AO22X1_LVT U1233 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[56]), .Y(io_resp_bits_data[56]) );
  AO22X1_LVT U1234 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[57]), .Y(io_resp_bits_data[57]) );
  AO22X1_LVT U1235 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[58]), .Y(io_resp_bits_data[58]) );
  AO22X1_LVT U1236 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[59]), .Y(io_resp_bits_data[59]) );
  AO22X1_LVT U1237 ( .A1(n146), .A2(result[37]), .A3(n209), .A4(result[5]), 
        .Y(io_resp_bits_data[5]) );
  AO22X1_LVT U1238 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[60]), .Y(io_resp_bits_data[60]) );
  AO22X1_LVT U1239 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[61]), .Y(io_resp_bits_data[61]) );
  AO22X1_LVT U1240 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[62]), .Y(io_resp_bits_data[62]) );
  AO22X1_LVT U1241 ( .A1(n244), .A2(io_resp_bits_data[31]), .A3(n242), .A4(
        result[63]), .Y(io_resp_bits_data[63]) );
  AO22X1_LVT U1242 ( .A1(n146), .A2(result[38]), .A3(n209), .A4(result[6]), 
        .Y(io_resp_bits_data[6]) );
  AO22X1_LVT U1243 ( .A1(n146), .A2(result[39]), .A3(n209), .A4(result[7]), 
        .Y(io_resp_bits_data[7]) );
  AO22X1_LVT U1244 ( .A1(n146), .A2(result[40]), .A3(n209), .A4(result[8]), 
        .Y(io_resp_bits_data[8]) );
  AO22X1_LVT U1245 ( .A1(n146), .A2(result[41]), .A3(n209), .A4(result[9]), 
        .Y(io_resp_bits_data[9]) );
  NAND4X0_LVT U1246 ( .A1(n757), .A2(n986), .A3(n985), .A4(n984), .Y(n996) );
  NAND4X0_LVT U1247 ( .A1(n756), .A2(n989), .A3(n988), .A4(n987), .Y(n995) );
  NAND4X0_LVT U1248 ( .A1(n755), .A2(n993), .A3(n992), .A4(n991), .Y(n994) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Rocket_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_LVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module Rocket_DW01_add_J37_0 ( A, B, CI, SUM, CO );
  input [38:0] A;
  input [38:0] B;
  output [38:0] SUM;
  input CI;
  output CO;
  wire   n125, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309;
  assign SUM[0] = A[0];

  HADDX1_LVT U160 ( .A0(A[2]), .B0(n259), .C1(n125), .SO(SUM[2]) );
  INVX1_LVT U170 ( .A(n301), .Y(n255) );
  INVX1_LVT U171 ( .A(n268), .Y(n257) );
  INVX1_LVT U172 ( .A(n286), .Y(n252) );
  INVX1_LVT U173 ( .A(n280), .Y(n253) );
  INVX1_LVT U174 ( .A(n290), .Y(n254) );
  INVX1_LVT U175 ( .A(n305), .Y(n256) );
  INVX1_LVT U176 ( .A(n272), .Y(n258) );
  INVX1_LVT U177 ( .A(n267), .Y(n259) );
  INVX1_LVT U178 ( .A(A[33]), .Y(n260) );
  INVX1_LVT U179 ( .A(A[29]), .Y(n261) );
  INVX1_LVT U180 ( .A(A[25]), .Y(n262) );
  INVX1_LVT U181 ( .A(A[17]), .Y(n263) );
  INVX1_LVT U182 ( .A(A[13]), .Y(n264) );
  INVX1_LVT U183 ( .A(A[9]), .Y(n265) );
  INVX1_LVT U184 ( .A(A[5]), .Y(n266) );
  AO22X1_LVT U185 ( .A1(n257), .A2(n265), .A3(n268), .A4(A[9]), .Y(SUM[9]) );
  HADDX1_LVT U186 ( .A0(A[8]), .B0(n269), .SO(SUM[8]) );
  AND2X1_LVT U187 ( .A1(A[7]), .A2(n270), .Y(n269) );
  HADDX1_LVT U188 ( .A0(A[7]), .B0(n270), .SO(SUM[7]) );
  HADDX1_LVT U189 ( .A0(n271), .B0(A[6]), .SO(SUM[6]) );
  AND2X1_LVT U190 ( .A1(n258), .A2(A[5]), .Y(n271) );
  AO22X1_LVT U191 ( .A1(A[5]), .A2(n272), .A3(n266), .A4(n258), .Y(SUM[5]) );
  HADDX1_LVT U192 ( .A0(A[4]), .B0(n273), .SO(SUM[4]) );
  AND2X1_LVT U193 ( .A1(n125), .A2(A[3]), .Y(n273) );
  HADDX1_LVT U194 ( .A0(n125), .B0(A[3]), .SO(SUM[3]) );
  HADDX1_LVT U195 ( .A0(n274), .B0(A[38]), .SO(SUM[38]) );
  AND2X1_LVT U196 ( .A1(n275), .A2(A[37]), .Y(n274) );
  HADDX1_LVT U197 ( .A0(A[37]), .B0(n275), .SO(SUM[37]) );
  AND2X1_LVT U198 ( .A1(n253), .A2(n276), .Y(n275) );
  AND4X1_LVT U199 ( .A1(A[34]), .A2(A[33]), .A3(A[35]), .A4(A[36]), .Y(n276)
         );
  HADDX1_LVT U200 ( .A0(A[36]), .B0(n277), .SO(SUM[36]) );
  AND4X1_LVT U201 ( .A1(A[34]), .A2(n253), .A3(A[33]), .A4(A[35]), .Y(n277) );
  HADDX1_LVT U202 ( .A0(n278), .B0(A[35]), .SO(SUM[35]) );
  AND3X1_LVT U203 ( .A1(n253), .A2(A[34]), .A3(A[33]), .Y(n278) );
  HADDX1_LVT U204 ( .A0(n279), .B0(A[34]), .SO(SUM[34]) );
  AND2X1_LVT U205 ( .A1(A[33]), .A2(n253), .Y(n279) );
  AO22X1_LVT U206 ( .A1(n253), .A2(n260), .A3(n280), .A4(A[33]), .Y(SUM[33])
         );
  NAND3X0_LVT U207 ( .A1(A[32]), .A2(A[31]), .A3(n281), .Y(n280) );
  AND4X1_LVT U208 ( .A1(A[29]), .A2(A[30]), .A3(n282), .A4(n254), .Y(n281) );
  HADDX1_LVT U209 ( .A0(A[32]), .B0(n283), .SO(SUM[32]) );
  AND4X1_LVT U210 ( .A1(A[31]), .A2(A[29]), .A3(A[30]), .A4(n252), .Y(n283) );
  HADDX1_LVT U211 ( .A0(A[31]), .B0(n284), .SO(SUM[31]) );
  AND3X1_LVT U212 ( .A1(A[29]), .A2(A[30]), .A3(n252), .Y(n284) );
  HADDX1_LVT U213 ( .A0(n285), .B0(A[30]), .SO(SUM[30]) );
  AND2X1_LVT U214 ( .A1(n252), .A2(A[29]), .Y(n285) );
  AO22X1_LVT U215 ( .A1(A[29]), .A2(n286), .A3(n261), .A4(n252), .Y(SUM[29])
         );
  NAND2X0_LVT U216 ( .A1(n282), .A2(n254), .Y(n286) );
  AND4X1_LVT U217 ( .A1(A[25]), .A2(A[26]), .A3(A[28]), .A4(A[27]), .Y(n282)
         );
  HADDX1_LVT U218 ( .A0(A[28]), .B0(n287), .SO(SUM[28]) );
  AND4X1_LVT U219 ( .A1(A[25]), .A2(A[26]), .A3(A[27]), .A4(n254), .Y(n287) );
  HADDX1_LVT U220 ( .A0(A[27]), .B0(n288), .SO(SUM[27]) );
  AND3X1_LVT U221 ( .A1(A[25]), .A2(A[26]), .A3(n254), .Y(n288) );
  HADDX1_LVT U222 ( .A0(n289), .B0(A[26]), .SO(SUM[26]) );
  AND2X1_LVT U223 ( .A1(n254), .A2(A[25]), .Y(n289) );
  AO22X1_LVT U224 ( .A1(A[25]), .A2(n290), .A3(n262), .A4(n254), .Y(SUM[25])
         );
  NAND2X0_LVT U225 ( .A1(n291), .A2(n255), .Y(n290) );
  AND4X1_LVT U226 ( .A1(A[23]), .A2(A[24]), .A3(n292), .A4(n293), .Y(n291) );
  HADDX1_LVT U227 ( .A0(A[24]), .B0(n294), .SO(SUM[24]) );
  AND4X1_LVT U228 ( .A1(A[23]), .A2(n292), .A3(n293), .A4(n255), .Y(n294) );
  HADDX1_LVT U229 ( .A0(A[23]), .B0(n295), .SO(SUM[23]) );
  AND3X1_LVT U230 ( .A1(n292), .A2(n293), .A3(n255), .Y(n295) );
  AND2X1_LVT U231 ( .A1(A[21]), .A2(A[22]), .Y(n292) );
  HADDX1_LVT U232 ( .A0(n296), .B0(A[22]), .SO(SUM[22]) );
  AND3X1_LVT U233 ( .A1(n293), .A2(A[21]), .A3(n255), .Y(n296) );
  HADDX1_LVT U234 ( .A0(A[21]), .B0(n297), .SO(SUM[21]) );
  AND2X1_LVT U235 ( .A1(n293), .A2(n255), .Y(n297) );
  AND4X1_LVT U236 ( .A1(A[17]), .A2(A[18]), .A3(A[20]), .A4(A[19]), .Y(n293)
         );
  HADDX1_LVT U237 ( .A0(A[20]), .B0(n298), .SO(SUM[20]) );
  AND4X1_LVT U238 ( .A1(A[17]), .A2(A[18]), .A3(A[19]), .A4(n255), .Y(n298) );
  OA21X1_LVT U239 ( .A1(A[1]), .A2(B[1]), .A3(n267), .Y(SUM[1]) );
  NAND2X0_LVT U240 ( .A1(A[1]), .A2(B[1]), .Y(n267) );
  HADDX1_LVT U241 ( .A0(A[19]), .B0(n299), .SO(SUM[19]) );
  AND3X1_LVT U242 ( .A1(A[17]), .A2(A[18]), .A3(n255), .Y(n299) );
  HADDX1_LVT U243 ( .A0(n300), .B0(A[18]), .SO(SUM[18]) );
  AND2X1_LVT U244 ( .A1(n255), .A2(A[17]), .Y(n300) );
  AO22X1_LVT U245 ( .A1(A[17]), .A2(n301), .A3(n263), .A4(n255), .Y(SUM[17])
         );
  NAND3X0_LVT U246 ( .A1(A[15]), .A2(A[16]), .A3(n302), .Y(n301) );
  HADDX1_LVT U247 ( .A0(A[16]), .B0(n303), .SO(SUM[16]) );
  AND4X1_LVT U248 ( .A1(A[13]), .A2(A[14]), .A3(A[15]), .A4(n256), .Y(n303) );
  HADDX1_LVT U249 ( .A0(A[15]), .B0(n302), .SO(SUM[15]) );
  AND3X1_LVT U250 ( .A1(A[13]), .A2(A[14]), .A3(n256), .Y(n302) );
  HADDX1_LVT U251 ( .A0(n304), .B0(A[14]), .SO(SUM[14]) );
  AND2X1_LVT U252 ( .A1(n256), .A2(A[13]), .Y(n304) );
  AO22X1_LVT U253 ( .A1(A[13]), .A2(n305), .A3(n264), .A4(n256), .Y(SUM[13])
         );
  NAND2X0_LVT U254 ( .A1(n257), .A2(n306), .Y(n305) );
  AND4X1_LVT U255 ( .A1(A[9]), .A2(A[10]), .A3(A[12]), .A4(A[11]), .Y(n306) );
  HADDX1_LVT U256 ( .A0(A[12]), .B0(n307), .SO(SUM[12]) );
  AND4X1_LVT U257 ( .A1(n257), .A2(A[9]), .A3(A[10]), .A4(A[11]), .Y(n307) );
  HADDX1_LVT U258 ( .A0(A[11]), .B0(n308), .SO(SUM[11]) );
  AND3X1_LVT U259 ( .A1(n257), .A2(A[9]), .A3(A[10]), .Y(n308) );
  HADDX1_LVT U260 ( .A0(n309), .B0(A[10]), .SO(SUM[10]) );
  AND2X1_LVT U261 ( .A1(A[9]), .A2(n257), .Y(n309) );
  NAND3X0_LVT U262 ( .A1(A[7]), .A2(A[8]), .A3(n270), .Y(n268) );
  AND3X1_LVT U263 ( .A1(A[5]), .A2(A[6]), .A3(n258), .Y(n270) );
  NAND3X0_LVT U264 ( .A1(n125), .A2(A[3]), .A3(A[4]), .Y(n272) );
endmodule


module Rocket_DW01_add_J37_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n246, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504;
  assign SUM[0] = A[0];

  FADDX1_LVT U319 ( .A(B[2]), .B(A[2]), .CI(n408), .CO(n246), .S(SUM[2]) );
  OA22X1_LVT U329 ( .A1(B[15]), .A2(A[15]), .A3(B[16]), .A4(A[16]), .Y(n394)
         );
  AND4X1_LVT U330 ( .A1(n410), .A2(n484), .A3(n394), .A4(n488), .Y(n395) );
  OA221X1_LVT U331 ( .A1(n485), .A2(n488), .A3(n485), .A4(n486), .A5(n394), 
        .Y(n396) );
  AO222X1_LVT U332 ( .A1(B[16]), .A2(A[16]), .A3(B[16]), .A4(n487), .A5(A[16]), 
        .A6(n487), .Y(n397) );
  OR3X1_LVT U333 ( .A1(n395), .A2(n396), .A3(n397), .Y(n440) );
  AO21X1_LVT U334 ( .A1(n415), .A2(n414), .A3(n416), .Y(n398) );
  OA22X1_LVT U335 ( .A1(B[7]), .A2(A[7]), .A3(B[8]), .A4(A[8]), .Y(n399) );
  OR2X1_LVT U336 ( .A1(B[8]), .A2(A[8]), .Y(n400) );
  AO222X1_LVT U337 ( .A1(n398), .A2(n399), .A3(n400), .A4(n413), .A5(A[8]), 
        .A6(B[8]), .Y(n410) );
  AO222X1_LVT U338 ( .A1(B[14]), .A2(A[14]), .A3(B[14]), .A4(n492), .A5(A[14]), 
        .A6(n492), .Y(n485) );
  AO222X1_LVT U339 ( .A1(B[18]), .A2(A[18]), .A3(B[18]), .A4(n482), .A5(A[18]), 
        .A6(n482), .Y(n478) );
  AO21X1_LVT U340 ( .A1(n465), .A2(n464), .A3(n466), .Y(n401) );
  AO221X1_LVT U341 ( .A1(n403), .A2(A[23]), .A3(n403), .A4(A[24]), .A5(n401), 
        .Y(n450) );
  AO222X1_LVT U342 ( .A1(B[10]), .A2(A[10]), .A3(B[10]), .A4(n501), .A5(A[10]), 
        .A6(n501), .Y(n497) );
  AO222X1_LVT U343 ( .A1(B[6]), .A2(A[6]), .A3(B[6]), .A4(n418), .A5(A[6]), 
        .A6(n418), .Y(n416) );
  INVX1_LVT U344 ( .A(B[39]), .Y(n404) );
  INVX0_LVT U345 ( .A(n424), .Y(n407) );
  OA221X1_LVT U346 ( .A1(n439), .A2(n440), .A3(n439), .A4(n441), .A5(n442), 
        .Y(n429) );
  NBUFFX2_LVT U347 ( .A(B[21]), .Y(n403) );
  OR2X1_LVT U348 ( .A1(n403), .A2(A[38]), .Y(n402) );
  AND2X1_LVT U349 ( .A1(n405), .A2(n406), .Y(n422) );
  AND2X1_LVT U350 ( .A1(n425), .A2(n423), .Y(n405) );
  NAND2X0_LVT U351 ( .A1(n402), .A2(n407), .Y(n406) );
  INVX1_LVT U352 ( .A(n409), .Y(n408) );
  FADDX1_LVT U353 ( .A(A[9]), .B(B[9]), .CI(n410), .S(SUM[9]) );
  FADDX1_LVT U354 ( .A(B[8]), .B(A[8]), .CI(n411), .S(SUM[8]) );
  AO221X1_LVT U355 ( .A1(n412), .A2(B[7]), .A3(n412), .A4(A[7]), .A5(n413), 
        .Y(n411) );
  FADDX1_LVT U356 ( .A(B[7]), .B(A[7]), .CI(n412), .S(SUM[7]) );
  AO21X1_LVT U357 ( .A1(n414), .A2(n415), .A3(n416), .Y(n412) );
  FADDX1_LVT U358 ( .A(B[6]), .B(A[6]), .CI(n417), .S(SUM[6]) );
  OA22X1_LVT U359 ( .A1(n415), .A2(n418), .A3(B[5]), .A4(A[5]), .Y(n417) );
  FADDX1_LVT U360 ( .A(n415), .B(B[5]), .CI(A[5]), .S(SUM[5]) );
  FADDX1_LVT U361 ( .A(B[4]), .B(A[4]), .CI(n419), .S(SUM[4]) );
  AO21X1_LVT U362 ( .A1(n246), .A2(n420), .A3(n421), .Y(n419) );
  FADDX1_LVT U363 ( .A(n246), .B(A[3]), .CI(B[3]), .S(SUM[3]) );
  FADDX1_LVT U364 ( .A(n422), .B(A[39]), .CI(n404), .S(SUM[39]) );
  NAND2X0_LVT U365 ( .A1(B[39]), .A2(A[38]), .Y(n425) );
  FADDX1_LVT U366 ( .A(n403), .B(A[38]), .CI(n426), .S(SUM[38]) );
  NAND2X0_LVT U367 ( .A1(n423), .A2(n424), .Y(n426) );
  NAND3X0_LVT U368 ( .A1(n427), .A2(n428), .A3(n429), .Y(n424) );
  OR2X1_LVT U369 ( .A1(A[37]), .A2(n403), .Y(n428) );
  AOI21X1_LVT U370 ( .A1(B[21]), .A2(A[37]), .A3(n430), .Y(n423) );
  FADDX1_LVT U371 ( .A(B[39]), .B(A[37]), .CI(n431), .S(SUM[37]) );
  AO21X1_LVT U372 ( .A1(n427), .A2(n429), .A3(n430), .Y(n431) );
  AO221X1_LVT U373 ( .A1(B[39]), .A2(A[35]), .A3(B[39]), .A4(A[36]), .A5(n432), 
        .Y(n430) );
  OA221X1_LVT U374 ( .A1(B[39]), .A2(A[35]), .A3(B[39]), .A4(A[36]), .A5(n433), 
        .Y(n427) );
  FADDX1_LVT U375 ( .A(n403), .B(n434), .CI(A[36]), .S(SUM[36]) );
  OA22X1_LVT U376 ( .A1(n435), .A2(n436), .A3(B[39]), .A4(A[35]), .Y(n434) );
  AND2X1_LVT U377 ( .A1(n403), .A2(A[35]), .Y(n435) );
  FADDX1_LVT U378 ( .A(n403), .B(A[35]), .CI(n436), .S(SUM[35]) );
  AO21X1_LVT U379 ( .A1(n433), .A2(n429), .A3(n432), .Y(n436) );
  OA21X1_LVT U380 ( .A1(A[33]), .A2(A[34]), .A3(B[39]), .Y(n432) );
  AO21X1_LVT U381 ( .A1(A[33]), .A2(A[34]), .A3(B[21]), .Y(n433) );
  FADDX1_LVT U382 ( .A(B[21]), .B(A[34]), .CI(n437), .S(SUM[34]) );
  AO22X1_LVT U383 ( .A1(n403), .A2(A[33]), .A3(n429), .A4(n438), .Y(n437) );
  OR2X1_LVT U384 ( .A1(n403), .A2(A[33]), .Y(n438) );
  FADDX1_LVT U385 ( .A(n403), .B(A[33]), .CI(n429), .S(SUM[33]) );
  AND4X1_LVT U386 ( .A1(n443), .A2(n444), .A3(n445), .A4(n446), .Y(n442) );
  OR2X1_LVT U387 ( .A1(B[21]), .A2(A[32]), .Y(n446) );
  OR3X1_LVT U388 ( .A1(n447), .A2(n448), .A3(n449), .Y(n439) );
  AO221X1_LVT U389 ( .A1(B[39]), .A2(A[31]), .A3(B[39]), .A4(A[32]), .A5(n450), 
        .Y(n449) );
  FADDX1_LVT U390 ( .A(n403), .B(A[32]), .CI(n451), .S(SUM[32]) );
  AO22X1_LVT U391 ( .A1(B[39]), .A2(A[31]), .A3(n452), .A4(n445), .Y(n451) );
  OR2X1_LVT U392 ( .A1(B[21]), .A2(A[31]), .Y(n445) );
  FADDX1_LVT U393 ( .A(n403), .B(A[31]), .CI(n452), .S(SUM[31]) );
  OA21X1_LVT U394 ( .A1(n453), .A2(n447), .A3(n443), .Y(n452) );
  AO21X1_LVT U395 ( .A1(A[30]), .A2(A[29]), .A3(B[21]), .Y(n443) );
  OA21X1_LVT U396 ( .A1(A[30]), .A2(A[29]), .A3(n403), .Y(n447) );
  FADDX1_LVT U397 ( .A(B[21]), .B(A[30]), .CI(n454), .S(SUM[30]) );
  AO22X1_LVT U398 ( .A1(n403), .A2(A[29]), .A3(n453), .A4(n455), .Y(n454) );
  OR2X1_LVT U399 ( .A1(n403), .A2(A[29]), .Y(n455) );
  FADDX1_LVT U400 ( .A(B[21]), .B(A[29]), .CI(n453), .S(SUM[29]) );
  OA21X1_LVT U401 ( .A1(n456), .A2(n448), .A3(n444), .Y(n453) );
  OA221X1_LVT U402 ( .A1(n403), .A2(A[27]), .A3(B[39]), .A4(A[28]), .A5(n457), 
        .Y(n444) );
  AO221X1_LVT U403 ( .A1(n403), .A2(A[27]), .A3(n403), .A4(A[28]), .A5(n458), 
        .Y(n448) );
  FADDX1_LVT U404 ( .A(B[39]), .B(A[28]), .CI(n459), .S(SUM[28]) );
  AO22X1_LVT U405 ( .A1(B[39]), .A2(A[27]), .A3(n460), .A4(n461), .Y(n459) );
  OR2X1_LVT U406 ( .A1(n403), .A2(A[27]), .Y(n461) );
  FADDX1_LVT U407 ( .A(B[21]), .B(A[27]), .CI(n460), .S(SUM[27]) );
  OA21X1_LVT U408 ( .A1(n456), .A2(n458), .A3(n457), .Y(n460) );
  AO21X1_LVT U409 ( .A1(A[26]), .A2(A[25]), .A3(n403), .Y(n457) );
  OA21X1_LVT U410 ( .A1(A[26]), .A2(A[25]), .A3(B[39]), .Y(n458) );
  FADDX1_LVT U411 ( .A(B[39]), .B(A[26]), .CI(n462), .S(SUM[26]) );
  AO22X1_LVT U412 ( .A1(n403), .A2(A[25]), .A3(n456), .A4(n463), .Y(n462) );
  OR2X1_LVT U413 ( .A1(n403), .A2(A[25]), .Y(n463) );
  FADDX1_LVT U414 ( .A(B[39]), .B(A[25]), .CI(n456), .S(SUM[25]) );
  AO21X1_LVT U415 ( .A1(n441), .A2(n440), .A3(n450), .Y(n456) );
  AND2X1_LVT U416 ( .A1(n467), .A2(n464), .Y(n441) );
  OA221X1_LVT U417 ( .A1(n403), .A2(A[23]), .A3(n403), .A4(A[24]), .A5(n468), 
        .Y(n464) );
  FADDX1_LVT U418 ( .A(n403), .B(A[24]), .CI(n469), .S(SUM[24]) );
  AO22X1_LVT U419 ( .A1(B[39]), .A2(A[23]), .A3(n470), .A4(n471), .Y(n469) );
  OR2X1_LVT U420 ( .A1(n403), .A2(A[23]), .Y(n471) );
  FADDX1_LVT U421 ( .A(n403), .B(A[23]), .CI(n470), .S(SUM[23]) );
  OA21X1_LVT U422 ( .A1(n472), .A2(n466), .A3(n468), .Y(n470) );
  AO21X1_LVT U423 ( .A1(A[22]), .A2(A[21]), .A3(n403), .Y(n468) );
  OA21X1_LVT U424 ( .A1(A[22]), .A2(A[21]), .A3(n403), .Y(n466) );
  FADDX1_LVT U425 ( .A(B[39]), .B(A[22]), .CI(n473), .S(SUM[22]) );
  AO22X1_LVT U426 ( .A1(n403), .A2(A[21]), .A3(n472), .A4(n474), .Y(n473) );
  OR2X1_LVT U427 ( .A1(n403), .A2(A[21]), .Y(n474) );
  FADDX1_LVT U428 ( .A(B[39]), .B(A[21]), .CI(n472), .S(SUM[21]) );
  AO21X1_LVT U429 ( .A1(n467), .A2(n440), .A3(n465), .Y(n472) );
  AO222X1_LVT U430 ( .A1(B[39]), .A2(A[20]), .A3(n475), .A4(n476), .A5(n477), 
        .A6(n478), .Y(n465) );
  OR2X1_LVT U431 ( .A1(A[20]), .A2(n403), .Y(n476) );
  AND2X1_LVT U432 ( .A1(n477), .A2(n479), .Y(n467) );
  OA22X1_LVT U433 ( .A1(B[39]), .A2(A[20]), .A3(B[19]), .A4(A[19]), .Y(n477)
         );
  FADDX1_LVT U434 ( .A(n403), .B(A[20]), .CI(n480), .S(SUM[20]) );
  AO221X1_LVT U435 ( .A1(n481), .A2(B[19]), .A3(n481), .A4(A[19]), .A5(n475), 
        .Y(n480) );
  AND2X1_LVT U436 ( .A1(B[19]), .A2(A[19]), .Y(n475) );
  OA21X1_LVT U437 ( .A1(A[1]), .A2(B[1]), .A3(n409), .Y(SUM[1]) );
  NAND2X0_LVT U438 ( .A1(A[1]), .A2(B[1]), .Y(n409) );
  FADDX1_LVT U439 ( .A(B[19]), .B(A[19]), .CI(n481), .S(SUM[19]) );
  AO21X1_LVT U440 ( .A1(n479), .A2(n440), .A3(n478), .Y(n481) );
  OA22X1_LVT U441 ( .A1(B[18]), .A2(A[18]), .A3(B[17]), .A4(A[17]), .Y(n479)
         );
  FADDX1_LVT U442 ( .A(B[18]), .B(A[18]), .CI(n483), .S(SUM[18]) );
  OA22X1_LVT U443 ( .A1(B[17]), .A2(A[17]), .A3(n482), .A4(n440), .Y(n483) );
  AND2X1_LVT U444 ( .A1(B[17]), .A2(A[17]), .Y(n482) );
  FADDX1_LVT U445 ( .A(B[17]), .B(A[17]), .CI(n440), .S(SUM[17]) );
  FADDX1_LVT U446 ( .A(B[16]), .B(A[16]), .CI(n489), .S(SUM[16]) );
  OA22X1_LVT U447 ( .A1(n487), .A2(n490), .A3(B[15]), .A4(A[15]), .Y(n489) );
  AND2X1_LVT U448 ( .A1(B[15]), .A2(A[15]), .Y(n487) );
  FADDX1_LVT U449 ( .A(B[15]), .B(A[15]), .CI(n490), .S(SUM[15]) );
  AO21X1_LVT U450 ( .A1(n488), .A2(n491), .A3(n485), .Y(n490) );
  OA22X1_LVT U451 ( .A1(B[14]), .A2(A[14]), .A3(B[13]), .A4(A[13]), .Y(n488)
         );
  FADDX1_LVT U452 ( .A(B[14]), .B(A[14]), .CI(n493), .S(SUM[14]) );
  OA22X1_LVT U453 ( .A1(n492), .A2(n491), .A3(B[13]), .A4(A[13]), .Y(n493) );
  AND2X1_LVT U454 ( .A1(B[13]), .A2(A[13]), .Y(n492) );
  FADDX1_LVT U455 ( .A(B[13]), .B(A[13]), .CI(n491), .S(SUM[13]) );
  AO21X1_LVT U456 ( .A1(n484), .A2(n410), .A3(n486), .Y(n491) );
  AO222X1_LVT U457 ( .A1(B[12]), .A2(A[12]), .A3(n494), .A4(n495), .A5(n496), 
        .A6(n497), .Y(n486) );
  OR2X1_LVT U458 ( .A1(A[12]), .A2(B[12]), .Y(n495) );
  AND2X1_LVT U459 ( .A1(n496), .A2(n498), .Y(n484) );
  OA22X1_LVT U460 ( .A1(B[12]), .A2(A[12]), .A3(B[11]), .A4(A[11]), .Y(n496)
         );
  FADDX1_LVT U461 ( .A(B[12]), .B(A[12]), .CI(n499), .S(SUM[12]) );
  OA22X1_LVT U462 ( .A1(n494), .A2(n500), .A3(B[11]), .A4(A[11]), .Y(n499) );
  AND2X1_LVT U463 ( .A1(B[11]), .A2(A[11]), .Y(n494) );
  FADDX1_LVT U464 ( .A(B[11]), .B(A[11]), .CI(n500), .S(SUM[11]) );
  AO21X1_LVT U465 ( .A1(n498), .A2(n410), .A3(n497), .Y(n500) );
  OA22X1_LVT U466 ( .A1(A[9]), .A2(B[9]), .A3(B[10]), .A4(A[10]), .Y(n498) );
  FADDX1_LVT U467 ( .A(B[10]), .B(A[10]), .CI(n502), .S(SUM[10]) );
  AO221X1_LVT U468 ( .A1(n410), .A2(A[9]), .A3(n410), .A4(B[9]), .A5(n501), 
        .Y(n502) );
  AND2X1_LVT U469 ( .A1(A[9]), .A2(B[9]), .Y(n501) );
  AND2X1_LVT U470 ( .A1(B[7]), .A2(A[7]), .Y(n413) );
  AND2X1_LVT U471 ( .A1(B[5]), .A2(A[5]), .Y(n418) );
  OA22X1_LVT U472 ( .A1(B[6]), .A2(A[6]), .A3(B[5]), .A4(A[5]), .Y(n414) );
  OA222X1_LVT U473 ( .A1(n503), .A2(n246), .A3(n503), .A4(n504), .A5(n503), 
        .A6(n420), .Y(n415) );
  OR2X1_LVT U474 ( .A1(A[3]), .A2(B[3]), .Y(n420) );
  AO22X1_LVT U475 ( .A1(B[4]), .A2(A[4]), .A3(n421), .A4(n504), .Y(n503) );
  OR2X1_LVT U476 ( .A1(B[4]), .A2(A[4]), .Y(n504) );
  AND2X1_LVT U477 ( .A1(A[3]), .A2(B[3]), .Y(n421) );
endmodule


module Rocket ( clock, reset, io_interrupts_debug, io_interrupts_mtip, 
        io_interrupts_msip, io_interrupts_meip, io_interrupts_seip, 
        io_imem_might_request, io_imem_req_valid, io_imem_req_bits_pc, 
        io_imem_req_bits_speculative, io_imem_sfence_valid, 
        io_imem_sfence_bits_rs1, io_imem_sfence_bits_rs2, 
        io_imem_sfence_bits_addr, io_imem_resp_ready, io_imem_resp_valid, 
        io_imem_resp_bits_btb_taken, io_imem_resp_bits_btb_bridx, 
        io_imem_resp_bits_btb_entry, io_imem_resp_bits_btb_bht_history, 
        io_imem_resp_bits_pc, io_imem_resp_bits_data, 
        io_imem_resp_bits_xcpt_pf_inst, io_imem_resp_bits_xcpt_ae_inst, 
        io_imem_resp_bits_replay, io_imem_btb_update_valid, 
        io_imem_btb_update_bits_prediction_entry, io_imem_btb_update_bits_pc, 
        io_imem_btb_update_bits_isValid, io_imem_btb_update_bits_br_pc, 
        io_imem_btb_update_bits_cfiType, io_imem_bht_update_valid, 
        io_imem_bht_update_bits_prediction_history, io_imem_bht_update_bits_pc, 
        io_imem_bht_update_bits_branch, io_imem_bht_update_bits_taken, 
        io_imem_bht_update_bits_mispredict, io_imem_flush_icache, 
        io_dmem_req_ready, io_dmem_req_valid, io_dmem_req_bits_addr, 
        io_dmem_req_bits_tag, io_dmem_req_bits_cmd, io_dmem_req_bits_size, 
        io_dmem_req_bits_signed, io_dmem_req_bits_dprv, io_dmem_s1_kill, 
        io_dmem_s1_data_data, io_dmem_s2_nack, io_dmem_resp_valid, 
        io_dmem_resp_bits_tag, io_dmem_resp_bits_size, io_dmem_resp_bits_data, 
        io_dmem_resp_bits_replay, io_dmem_resp_bits_has_data, 
        io_dmem_resp_bits_data_word_bypass, io_dmem_replay_next, 
        io_dmem_s2_xcpt_ma_ld, io_dmem_s2_xcpt_ma_st, io_dmem_s2_xcpt_pf_ld, 
        io_dmem_s2_xcpt_pf_st, io_dmem_s2_xcpt_ae_ld, io_dmem_s2_xcpt_ae_st, 
        io_dmem_ordered, io_dmem_perf_release, io_dmem_perf_grant, 
        io_ptw_ptbr_mode, io_ptw_ptbr_ppn, io_ptw_sfence_valid, 
        io_ptw_sfence_bits_rs1, io_ptw_sfence_bits_rs2, 
        io_ptw_sfence_bits_addr, io_ptw_status_debug, io_ptw_status_dprv, 
        io_ptw_status_prv, io_ptw_status_mxr, io_ptw_status_sum, 
        io_ptw_pmp_0_cfg_l, io_ptw_pmp_0_cfg_a, io_ptw_pmp_0_cfg_x, 
        io_ptw_pmp_0_cfg_w, io_ptw_pmp_0_cfg_r, io_ptw_pmp_0_addr, 
        io_ptw_pmp_0_mask, io_ptw_pmp_1_cfg_l, io_ptw_pmp_1_cfg_a, 
        io_ptw_pmp_1_cfg_x, io_ptw_pmp_1_cfg_w, io_ptw_pmp_1_cfg_r, 
        io_ptw_pmp_1_addr, io_ptw_pmp_1_mask, io_ptw_pmp_2_cfg_l, 
        io_ptw_pmp_2_cfg_a, io_ptw_pmp_2_cfg_x, io_ptw_pmp_2_cfg_w, 
        io_ptw_pmp_2_cfg_r, io_ptw_pmp_2_addr, io_ptw_pmp_2_mask, 
        io_ptw_pmp_3_cfg_l, io_ptw_pmp_3_cfg_a, io_ptw_pmp_3_cfg_x, 
        io_ptw_pmp_3_cfg_w, io_ptw_pmp_3_cfg_r, io_ptw_pmp_3_addr, 
        io_ptw_pmp_3_mask, io_ptw_pmp_4_cfg_l, io_ptw_pmp_4_cfg_a, 
        io_ptw_pmp_4_cfg_x, io_ptw_pmp_4_cfg_w, io_ptw_pmp_4_cfg_r, 
        io_ptw_pmp_4_addr, io_ptw_pmp_4_mask, io_ptw_pmp_5_cfg_l, 
        io_ptw_pmp_5_cfg_a, io_ptw_pmp_5_cfg_x, io_ptw_pmp_5_cfg_w, 
        io_ptw_pmp_5_cfg_r, io_ptw_pmp_5_addr, io_ptw_pmp_5_mask, 
        io_ptw_pmp_6_cfg_l, io_ptw_pmp_6_cfg_a, io_ptw_pmp_6_cfg_x, 
        io_ptw_pmp_6_cfg_w, io_ptw_pmp_6_cfg_r, io_ptw_pmp_6_addr, 
        io_ptw_pmp_6_mask, io_ptw_pmp_7_cfg_l, io_ptw_pmp_7_cfg_a, 
        io_ptw_pmp_7_cfg_x, io_ptw_pmp_7_cfg_w, io_ptw_pmp_7_cfg_r, 
        io_ptw_pmp_7_addr, io_ptw_pmp_7_mask, io_ptw_customCSRs_csrs_0_value, 
        io_fpu_inst, io_fpu_fromint_data, io_fpu_fcsr_rm, 
        io_fpu_fcsr_flags_valid, io_fpu_fcsr_flags_bits, io_fpu_store_data, 
        io_fpu_toint_data, io_fpu_dmem_resp_val, io_fpu_dmem_resp_type, 
        io_fpu_dmem_resp_tag, io_fpu_dmem_resp_data, io_fpu_valid, 
        io_fpu_fcsr_rdy, io_fpu_nack_mem, io_fpu_illegal_rm, io_fpu_killx, 
        io_fpu_killm, io_fpu_dec_wen, io_fpu_dec_ren1, io_fpu_dec_ren2, 
        io_fpu_dec_ren3, io_fpu_sboard_set, io_fpu_sboard_clr, 
        io_fpu_sboard_clra, io_wfi );
  output [39:0] io_imem_req_bits_pc;
  output [38:0] io_imem_sfence_bits_addr;
  input [4:0] io_imem_resp_bits_btb_entry;
  input [7:0] io_imem_resp_bits_btb_bht_history;
  input [39:0] io_imem_resp_bits_pc;
  input [31:0] io_imem_resp_bits_data;
  output [4:0] io_imem_btb_update_bits_prediction_entry;
  output [38:0] io_imem_btb_update_bits_pc;
  output [38:0] io_imem_btb_update_bits_br_pc;
  output [1:0] io_imem_btb_update_bits_cfiType;
  output [7:0] io_imem_bht_update_bits_prediction_history;
  output [38:0] io_imem_bht_update_bits_pc;
  output [39:0] io_dmem_req_bits_addr;
  output [6:0] io_dmem_req_bits_tag;
  output [4:0] io_dmem_req_bits_cmd;
  output [1:0] io_dmem_req_bits_size;
  output [1:0] io_dmem_req_bits_dprv;
  output [63:0] io_dmem_s1_data_data;
  input [6:0] io_dmem_resp_bits_tag;
  input [1:0] io_dmem_resp_bits_size;
  input [63:0] io_dmem_resp_bits_data;
  input [63:0] io_dmem_resp_bits_data_word_bypass;
  output [3:0] io_ptw_ptbr_mode;
  output [43:0] io_ptw_ptbr_ppn;
  output [38:0] io_ptw_sfence_bits_addr;
  output [1:0] io_ptw_status_dprv;
  output [1:0] io_ptw_status_prv;
  output [1:0] io_ptw_pmp_0_cfg_a;
  output [29:0] io_ptw_pmp_0_addr;
  output [31:0] io_ptw_pmp_0_mask;
  output [1:0] io_ptw_pmp_1_cfg_a;
  output [29:0] io_ptw_pmp_1_addr;
  output [31:0] io_ptw_pmp_1_mask;
  output [1:0] io_ptw_pmp_2_cfg_a;
  output [29:0] io_ptw_pmp_2_addr;
  output [31:0] io_ptw_pmp_2_mask;
  output [1:0] io_ptw_pmp_3_cfg_a;
  output [29:0] io_ptw_pmp_3_addr;
  output [31:0] io_ptw_pmp_3_mask;
  output [1:0] io_ptw_pmp_4_cfg_a;
  output [29:0] io_ptw_pmp_4_addr;
  output [31:0] io_ptw_pmp_4_mask;
  output [1:0] io_ptw_pmp_5_cfg_a;
  output [29:0] io_ptw_pmp_5_addr;
  output [31:0] io_ptw_pmp_5_mask;
  output [1:0] io_ptw_pmp_6_cfg_a;
  output [29:0] io_ptw_pmp_6_addr;
  output [31:0] io_ptw_pmp_6_mask;
  output [1:0] io_ptw_pmp_7_cfg_a;
  output [29:0] io_ptw_pmp_7_addr;
  output [31:0] io_ptw_pmp_7_mask;
  output [63:0] io_ptw_customCSRs_csrs_0_value;
  output [31:0] io_fpu_inst;
  output [63:0] io_fpu_fromint_data;
  output [2:0] io_fpu_fcsr_rm;
  input [4:0] io_fpu_fcsr_flags_bits;
  input [63:0] io_fpu_store_data;
  input [63:0] io_fpu_toint_data;
  output [2:0] io_fpu_dmem_resp_type;
  output [4:0] io_fpu_dmem_resp_tag;
  output [63:0] io_fpu_dmem_resp_data;
  input [4:0] io_fpu_sboard_clra;
  input clock, reset, io_interrupts_debug, io_interrupts_mtip,
         io_interrupts_msip, io_interrupts_meip, io_interrupts_seip,
         io_imem_resp_valid, io_imem_resp_bits_btb_taken,
         io_imem_resp_bits_btb_bridx, io_imem_resp_bits_xcpt_pf_inst,
         io_imem_resp_bits_xcpt_ae_inst, io_imem_resp_bits_replay,
         io_dmem_req_ready, io_dmem_s2_nack, io_dmem_resp_valid,
         io_dmem_resp_bits_replay, io_dmem_resp_bits_has_data,
         io_dmem_replay_next, io_dmem_s2_xcpt_ma_ld, io_dmem_s2_xcpt_ma_st,
         io_dmem_s2_xcpt_pf_ld, io_dmem_s2_xcpt_pf_st, io_dmem_s2_xcpt_ae_ld,
         io_dmem_s2_xcpt_ae_st, io_dmem_ordered, io_dmem_perf_release,
         io_dmem_perf_grant, io_fpu_fcsr_flags_valid, io_fpu_fcsr_rdy,
         io_fpu_nack_mem, io_fpu_illegal_rm, io_fpu_dec_wen, io_fpu_dec_ren1,
         io_fpu_dec_ren2, io_fpu_dec_ren3, io_fpu_sboard_set,
         io_fpu_sboard_clr;
  output io_imem_might_request, io_imem_req_valid,
         io_imem_req_bits_speculative, io_imem_sfence_valid,
         io_imem_sfence_bits_rs1, io_imem_sfence_bits_rs2, io_imem_resp_ready,
         io_imem_btb_update_valid, io_imem_btb_update_bits_isValid,
         io_imem_bht_update_valid, io_imem_bht_update_bits_branch,
         io_imem_bht_update_bits_taken, io_imem_bht_update_bits_mispredict,
         io_imem_flush_icache, io_dmem_req_valid, io_dmem_req_bits_signed,
         io_dmem_s1_kill, io_ptw_sfence_valid, io_ptw_sfence_bits_rs1,
         io_ptw_sfence_bits_rs2, io_ptw_status_debug, io_ptw_status_mxr,
         io_ptw_status_sum, io_ptw_pmp_0_cfg_l, io_ptw_pmp_0_cfg_x,
         io_ptw_pmp_0_cfg_w, io_ptw_pmp_0_cfg_r, io_ptw_pmp_1_cfg_l,
         io_ptw_pmp_1_cfg_x, io_ptw_pmp_1_cfg_w, io_ptw_pmp_1_cfg_r,
         io_ptw_pmp_2_cfg_l, io_ptw_pmp_2_cfg_x, io_ptw_pmp_2_cfg_w,
         io_ptw_pmp_2_cfg_r, io_ptw_pmp_3_cfg_l, io_ptw_pmp_3_cfg_x,
         io_ptw_pmp_3_cfg_w, io_ptw_pmp_3_cfg_r, io_ptw_pmp_4_cfg_l,
         io_ptw_pmp_4_cfg_x, io_ptw_pmp_4_cfg_w, io_ptw_pmp_4_cfg_r,
         io_ptw_pmp_5_cfg_l, io_ptw_pmp_5_cfg_x, io_ptw_pmp_5_cfg_w,
         io_ptw_pmp_5_cfg_r, io_ptw_pmp_6_cfg_l, io_ptw_pmp_6_cfg_x,
         io_ptw_pmp_6_cfg_w, io_ptw_pmp_6_cfg_r, io_ptw_pmp_7_cfg_l,
         io_ptw_pmp_7_cfg_x, io_ptw_pmp_7_cfg_w, io_ptw_pmp_7_cfg_r,
         io_fpu_dmem_resp_val, io_fpu_valid, io_fpu_killx, io_fpu_killm,
         io_wfi;
  wire   io_imem_sfence_valid, io_imem_sfence_bits_rs1,
         io_imem_sfence_bits_rs2, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         ibuf_io_inst_0_valid, ibuf_io_inst_0_bits_replay,
         ibuf_io_inst_0_bits_rvc, csr_io_rw_cmd_2_, csr_io_decode_0_fp_illegal,
         csr_io_decode_0_fp_csr, csr_io_decode_0_read_illegal,
         csr_io_decode_0_write_illegal, csr_io_decode_0_write_flush,
         csr_io_decode_0_system_illegal, csr_io_csr_stall, csr_io_eret,
         csr_io_singleStep, csr_io_exception, csr_io_retire, csr_io_interrupt,
         csr_io_bp_0_control_action, csr_io_bp_0_control_m,
         csr_io_bp_0_control_s, csr_io_bp_0_control_u, csr_io_bp_0_control_x,
         csr_io_bp_0_control_w, csr_io_bp_0_control_r, bpu_io_xcpt_if,
         bpu_io_xcpt_ld, bpu_io_xcpt_st, bpu_io_debug_if, bpu_io_debug_ld,
         bpu_io_debug_st, alu_io_dw, alu_io_adder_out_39_, alu_io_cmp_out,
         div_io_req_ready, div_io_kill, div_io_resp_ready, div_io_resp_valid,
         wb_reg_replay, wb_reg_valid, wb_ctrl_mem, wb_reg_flush_pipe,
         ex_reg_valid, ex_reg_replay, ex_reg_xcpt_interrupt, mem_ctrl_jalr,
         mem_reg_sfence, n_T_844_10_, n_T_911_11, mem_reg_rvc, mem_reg_valid,
         id_ctrl_mem_cmd_2_, id_ctrl_wfd, id_ctrl_wxd, id_reg_fence,
         ex_reg_inst_31_, ex_ctrl_wxd, mem_ctrl_wxd, mem_ctrl_mem,
         ex_reg_rs_bypass_1, ex_ctrl_sel_alu1_0_, ex_reg_rvc, ex_ctrl_jalr,
         ex_ctrl_mem, ex_ctrl_div, ex_ctrl_wfd, mem_reg_slow_bypass,
         mem_ctrl_wfd, wb_ctrl_wxd, wb_ctrl_div, wb_ctrl_wfd, blocked,
         id_reg_pause, n_GEN_9, n_T_731, do_bypass_1, n_T_760, ex_reg_load_use,
         mem_reg_replay, mem_reg_xcpt_interrupt, mem_pc_valid, mem_reg_xcpt,
         mem_reg_flush_pipe, ex_ctrl_rxs2, mem_reg_load, mem_reg_store,
         wb_ctrl_fence_i, wb_reg_sfence, n_T_1057, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N271, N274, N275, N279, N282, N283,
         N284, N286, N290, ex_ctrl_jal, N303, N304, N369, N370, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503,
         N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514,
         N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N526,
         N529, N530, N533, N535, N536, N598, N599, N600, N601, N602, N603,
         N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658,
         N659, N660, N661, N672, N673, N678, N679, N682, N683, N684, N685,
         N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696,
         N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707,
         N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729,
         N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740,
         N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751,
         N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, net34469, net34475, net34480, net34485,
         net34490, net34495, net34500, net34505, net34510, net34515, net34520,
         net34525, net34530, net34535, net34540, net34545, net34550, net34555,
         net34560, net34565, net34570, net34575, net34580, net34585, net34590,
         net34595, net34600, net34605, net34610, net34615, net34620, net34625,
         net34630, net34635, net34640, net34645, net34650, net34655, net34660,
         net34665, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n66, n67, n68, n69, n71, n72, n73, n74, n75, n76, n80, n98, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n308, n309, n310, n312, n313, n314,
         n315, n317, n318, n319, n320, n322, n323, n326, n369, n370, n406,
         n407, n546, n555, n559, n560, n561, n569, n570, n572, n576, n586,
         n588, n589, n590, n591, n592, n594, n595, n596, n598, n711, n882,
         n996, n997, n1262, n1279, n1281, n1431, n1531, n1532, n1589, n1612,
         n1628, n1699, n1820, n1821, n1822, n1823, n1828, n1829, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1855, n1856, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2238, n2239, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2501, n2507, n2510, n2512,
         n2514, n2515, n2516, n2518, n2521, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2541, n2542, n2543, n2544, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3046, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9417, n9418,
         n9421, n9422, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346;
  wire   [39:0] ibuf_io_pc;
  wire   [4:0] ibuf_io_btb_resp_entry;
  wire   [7:0] ibuf_io_btb_resp_bht_history;
  wire   [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire   [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire   [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire   [30:0] ibuf_io_inst_0_bits_raw;
  wire   [11:0] csr_io_rw_addr;
  wire   [63:0] csr_io_rw_rdata;
  wire   [12:0] csr_io_status_isa;
  wire   [39:1] csr_io_evec;
  wire   [39:0] csr_io_pc;
  wire   [39:0] csr_io_tval;
  wire   [31:0] csr_io_time;
  wire   [3:0] csr_io_interrupt_cause;
  wire   [1:0] csr_io_bp_0_control_tmatch;
  wire   [38:0] csr_io_bp_0_address;
  wire   [3:0] alu_io_fn;
  wire   [63:0] alu_io_in2;
  wire   [63:0] alu_io_in1;
  wire   [63:0] alu_io_out;
  wire   [63:0] div_io_resp_bits_data;
  wire   [4:0] div_io_resp_bits_tag;
  wire   [1942:0] n_T_427;
  wire   [63:0] n_T_427__T_1136_data;
  wire   [63:0] n_T_918;
  wire   [11:1] n_T_849;
  wire   [7:0] n_T_904;
  wire   [4:1] n_T_911;
  wire   [19:1] n_T_914;
  wire   [39:0] mem_reg_pc;
  wire   [39:0] mem_br_target;
  wire   [2:0] id_ctrl_sel_imm;
  wire   [4:1] wb_waddr;
  wire   [63:1] n_T_628;
  wire   [63:1] n_T_635;
  wire   [2:0] ex_ctrl_sel_imm;
  wire   [10:0] n_T_642;
  wire   [7:0] n_T_648;
  wire   [39:0] n_T_698;
  wire   [63:0] n_T_702;
  wire   [1:0] ex_ctrl_sel_alu2;
  wire   [2:0] ex_ctrl_csr;
  wire   [2:0] mem_ctrl_csr;
  wire   [31:1] n_T_1187;
  wire   [31:0] n_T_1298;
  wire   [1:0] n_T_726;
  wire   [1:0] n_T_728;
  wire   [2:0] wb_ctrl_csr;
  wire   [63:2] id_rs_1;
  wire   [63:0] wb_cause;
  wire   [63:0] wb_reg_cause;
  wire   [63:39] n_T_1165;
  wire   [63:0] mem_reg_rs2;
  wire   [63:0] mem_reg_cause;
  assign io_ptw_sfence_valid = io_imem_sfence_valid;
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1;
  assign io_ptw_sfence_bits_rs2 = io_imem_sfence_bits_rs2;
  assign io_ptw_sfence_bits_addr[38] = io_imem_sfence_bits_addr[38];
  assign io_ptw_sfence_bits_addr[37] = io_imem_sfence_bits_addr[37];
  assign io_ptw_sfence_bits_addr[36] = io_imem_sfence_bits_addr[36];
  assign io_ptw_sfence_bits_addr[35] = io_imem_sfence_bits_addr[35];
  assign io_ptw_sfence_bits_addr[34] = io_imem_sfence_bits_addr[34];
  assign io_ptw_sfence_bits_addr[33] = io_imem_sfence_bits_addr[33];
  assign io_ptw_sfence_bits_addr[32] = io_imem_sfence_bits_addr[32];
  assign io_ptw_sfence_bits_addr[31] = io_imem_sfence_bits_addr[31];
  assign io_ptw_sfence_bits_addr[30] = io_imem_sfence_bits_addr[30];
  assign io_ptw_sfence_bits_addr[29] = io_imem_sfence_bits_addr[29];
  assign io_ptw_sfence_bits_addr[28] = io_imem_sfence_bits_addr[28];
  assign io_ptw_sfence_bits_addr[27] = io_imem_sfence_bits_addr[27];
  assign io_ptw_sfence_bits_addr[26] = io_imem_sfence_bits_addr[26];
  assign io_ptw_sfence_bits_addr[25] = io_imem_sfence_bits_addr[25];
  assign io_ptw_sfence_bits_addr[24] = io_imem_sfence_bits_addr[24];
  assign io_ptw_sfence_bits_addr[23] = io_imem_sfence_bits_addr[23];
  assign io_ptw_sfence_bits_addr[22] = io_imem_sfence_bits_addr[22];
  assign io_ptw_sfence_bits_addr[21] = io_imem_sfence_bits_addr[21];
  assign io_ptw_sfence_bits_addr[20] = io_imem_sfence_bits_addr[20];
  assign io_ptw_sfence_bits_addr[19] = io_imem_sfence_bits_addr[19];
  assign io_ptw_sfence_bits_addr[18] = io_imem_sfence_bits_addr[18];
  assign io_ptw_sfence_bits_addr[17] = io_imem_sfence_bits_addr[17];
  assign io_ptw_sfence_bits_addr[16] = io_imem_sfence_bits_addr[16];
  assign io_ptw_sfence_bits_addr[15] = io_imem_sfence_bits_addr[15];
  assign io_ptw_sfence_bits_addr[14] = io_imem_sfence_bits_addr[14];
  assign io_ptw_sfence_bits_addr[13] = io_imem_sfence_bits_addr[13];
  assign io_ptw_sfence_bits_addr[12] = io_imem_sfence_bits_addr[12];
  assign io_ptw_sfence_bits_addr[11] = io_imem_sfence_bits_addr[11];
  assign io_ptw_sfence_bits_addr[10] = io_imem_sfence_bits_addr[10];
  assign io_ptw_sfence_bits_addr[9] = io_imem_sfence_bits_addr[9];
  assign io_ptw_sfence_bits_addr[8] = io_imem_sfence_bits_addr[8];
  assign io_ptw_sfence_bits_addr[7] = io_imem_sfence_bits_addr[7];
  assign io_ptw_sfence_bits_addr[6] = io_imem_sfence_bits_addr[6];
  assign io_ptw_sfence_bits_addr[5] = io_imem_sfence_bits_addr[5];
  assign io_ptw_sfence_bits_addr[4] = io_imem_sfence_bits_addr[4];
  assign io_ptw_sfence_bits_addr[3] = io_imem_sfence_bits_addr[3];
  assign io_ptw_sfence_bits_addr[2] = io_imem_sfence_bits_addr[2];
  assign io_ptw_sfence_bits_addr[1] = io_imem_sfence_bits_addr[1];
  assign io_ptw_sfence_bits_addr[0] = io_imem_sfence_bits_addr[0];
  assign io_imem_bht_update_bits_pc[38] = io_imem_btb_update_bits_br_pc[38];
  assign io_imem_btb_update_bits_pc[38] = io_imem_btb_update_bits_br_pc[38];
  assign io_imem_bht_update_bits_pc[37] = io_imem_btb_update_bits_br_pc[37];
  assign io_imem_btb_update_bits_pc[37] = io_imem_btb_update_bits_br_pc[37];
  assign io_imem_bht_update_bits_pc[36] = io_imem_btb_update_bits_br_pc[36];
  assign io_imem_btb_update_bits_pc[36] = io_imem_btb_update_bits_br_pc[36];
  assign io_imem_bht_update_bits_pc[35] = io_imem_btb_update_bits_br_pc[35];
  assign io_imem_btb_update_bits_pc[35] = io_imem_btb_update_bits_br_pc[35];
  assign io_imem_bht_update_bits_pc[34] = io_imem_btb_update_bits_br_pc[34];
  assign io_imem_btb_update_bits_pc[34] = io_imem_btb_update_bits_br_pc[34];
  assign io_imem_bht_update_bits_pc[33] = io_imem_btb_update_bits_br_pc[33];
  assign io_imem_btb_update_bits_pc[33] = io_imem_btb_update_bits_br_pc[33];
  assign io_imem_bht_update_bits_pc[32] = io_imem_btb_update_bits_br_pc[32];
  assign io_imem_btb_update_bits_pc[32] = io_imem_btb_update_bits_br_pc[32];
  assign io_imem_bht_update_bits_pc[31] = io_imem_btb_update_bits_br_pc[31];
  assign io_imem_btb_update_bits_pc[31] = io_imem_btb_update_bits_br_pc[31];
  assign io_imem_bht_update_bits_pc[30] = io_imem_btb_update_bits_br_pc[30];
  assign io_imem_btb_update_bits_pc[30] = io_imem_btb_update_bits_br_pc[30];
  assign io_imem_bht_update_bits_pc[29] = io_imem_btb_update_bits_br_pc[29];
  assign io_imem_btb_update_bits_pc[29] = io_imem_btb_update_bits_br_pc[29];
  assign io_imem_bht_update_bits_pc[28] = io_imem_btb_update_bits_br_pc[28];
  assign io_imem_btb_update_bits_pc[28] = io_imem_btb_update_bits_br_pc[28];
  assign io_imem_bht_update_bits_pc[27] = io_imem_btb_update_bits_br_pc[27];
  assign io_imem_btb_update_bits_pc[27] = io_imem_btb_update_bits_br_pc[27];
  assign io_imem_bht_update_bits_pc[26] = io_imem_btb_update_bits_br_pc[26];
  assign io_imem_btb_update_bits_pc[26] = io_imem_btb_update_bits_br_pc[26];
  assign io_imem_bht_update_bits_pc[25] = io_imem_btb_update_bits_br_pc[25];
  assign io_imem_btb_update_bits_pc[25] = io_imem_btb_update_bits_br_pc[25];
  assign io_imem_bht_update_bits_pc[24] = io_imem_btb_update_bits_br_pc[24];
  assign io_imem_btb_update_bits_pc[24] = io_imem_btb_update_bits_br_pc[24];
  assign io_imem_bht_update_bits_pc[23] = io_imem_btb_update_bits_br_pc[23];
  assign io_imem_btb_update_bits_pc[23] = io_imem_btb_update_bits_br_pc[23];
  assign io_imem_bht_update_bits_pc[22] = io_imem_btb_update_bits_br_pc[22];
  assign io_imem_btb_update_bits_pc[22] = io_imem_btb_update_bits_br_pc[22];
  assign io_imem_bht_update_bits_pc[21] = io_imem_btb_update_bits_br_pc[21];
  assign io_imem_btb_update_bits_pc[21] = io_imem_btb_update_bits_br_pc[21];
  assign io_imem_bht_update_bits_pc[20] = io_imem_btb_update_bits_br_pc[20];
  assign io_imem_btb_update_bits_pc[20] = io_imem_btb_update_bits_br_pc[20];
  assign io_imem_bht_update_bits_pc[19] = io_imem_btb_update_bits_br_pc[19];
  assign io_imem_btb_update_bits_pc[19] = io_imem_btb_update_bits_br_pc[19];
  assign io_imem_bht_update_bits_pc[18] = io_imem_btb_update_bits_br_pc[18];
  assign io_imem_btb_update_bits_pc[18] = io_imem_btb_update_bits_br_pc[18];
  assign io_imem_bht_update_bits_pc[17] = io_imem_btb_update_bits_br_pc[17];
  assign io_imem_btb_update_bits_pc[17] = io_imem_btb_update_bits_br_pc[17];
  assign io_imem_bht_update_bits_pc[16] = io_imem_btb_update_bits_br_pc[16];
  assign io_imem_btb_update_bits_pc[16] = io_imem_btb_update_bits_br_pc[16];
  assign io_imem_bht_update_bits_pc[15] = io_imem_btb_update_bits_br_pc[15];
  assign io_imem_btb_update_bits_pc[15] = io_imem_btb_update_bits_br_pc[15];
  assign io_imem_bht_update_bits_pc[14] = io_imem_btb_update_bits_br_pc[14];
  assign io_imem_btb_update_bits_pc[14] = io_imem_btb_update_bits_br_pc[14];
  assign io_imem_bht_update_bits_pc[13] = io_imem_btb_update_bits_br_pc[13];
  assign io_imem_btb_update_bits_pc[13] = io_imem_btb_update_bits_br_pc[13];
  assign io_imem_bht_update_bits_pc[12] = io_imem_btb_update_bits_br_pc[12];
  assign io_imem_btb_update_bits_pc[12] = io_imem_btb_update_bits_br_pc[12];
  assign io_imem_bht_update_bits_pc[11] = io_imem_btb_update_bits_br_pc[11];
  assign io_imem_btb_update_bits_pc[11] = io_imem_btb_update_bits_br_pc[11];
  assign io_imem_bht_update_bits_pc[10] = io_imem_btb_update_bits_br_pc[10];
  assign io_imem_btb_update_bits_pc[10] = io_imem_btb_update_bits_br_pc[10];
  assign io_imem_bht_update_bits_pc[9] = io_imem_btb_update_bits_br_pc[9];
  assign io_imem_btb_update_bits_pc[9] = io_imem_btb_update_bits_br_pc[9];
  assign io_imem_bht_update_bits_pc[8] = io_imem_btb_update_bits_br_pc[8];
  assign io_imem_btb_update_bits_pc[8] = io_imem_btb_update_bits_br_pc[8];
  assign io_imem_bht_update_bits_pc[7] = io_imem_btb_update_bits_br_pc[7];
  assign io_imem_btb_update_bits_pc[7] = io_imem_btb_update_bits_br_pc[7];
  assign io_imem_bht_update_bits_pc[6] = io_imem_btb_update_bits_br_pc[6];
  assign io_imem_btb_update_bits_pc[6] = io_imem_btb_update_bits_br_pc[6];
  assign io_imem_bht_update_bits_pc[5] = io_imem_btb_update_bits_br_pc[5];
  assign io_imem_btb_update_bits_pc[5] = io_imem_btb_update_bits_br_pc[5];
  assign io_imem_bht_update_bits_pc[4] = io_imem_btb_update_bits_br_pc[4];
  assign io_imem_btb_update_bits_pc[4] = io_imem_btb_update_bits_br_pc[4];
  assign io_imem_bht_update_bits_pc[3] = io_imem_btb_update_bits_br_pc[3];
  assign io_imem_btb_update_bits_pc[3] = io_imem_btb_update_bits_br_pc[3];
  assign io_imem_bht_update_bits_pc[2] = io_imem_btb_update_bits_br_pc[2];
  assign io_imem_btb_update_bits_pc[2] = io_imem_btb_update_bits_br_pc[2];
  assign io_ptw_status_dprv[1] = io_dmem_req_bits_dprv[1];
  assign io_ptw_status_dprv[0] = io_dmem_req_bits_dprv[0];
  assign io_dmem_req_bits_tag[6] = 1'b0;
  assign io_fpu_dmem_resp_type[2] = 1'b0;
  assign io_imem_btb_update_bits_pc[1] = 1'b0;
  assign io_imem_btb_update_bits_pc[0] = 1'b0;
  assign io_imem_bht_update_bits_pc[1] = 1'b0;
  assign io_imem_bht_update_bits_pc[0] = 1'b0;
  assign io_ptw_ptbr_mode[0] = 1'b0;
  assign io_ptw_ptbr_mode[1] = 1'b0;
  assign io_ptw_ptbr_mode[2] = 1'b0;
  assign io_ptw_ptbr_ppn[20] = 1'b0;
  assign io_ptw_ptbr_ppn[21] = 1'b0;
  assign io_ptw_ptbr_ppn[22] = 1'b0;
  assign io_ptw_ptbr_ppn[23] = 1'b0;
  assign io_ptw_ptbr_ppn[24] = 1'b0;
  assign io_ptw_ptbr_ppn[25] = 1'b0;
  assign io_ptw_ptbr_ppn[26] = 1'b0;
  assign io_ptw_ptbr_ppn[27] = 1'b0;
  assign io_ptw_ptbr_ppn[28] = 1'b0;
  assign io_ptw_ptbr_ppn[29] = 1'b0;
  assign io_ptw_ptbr_ppn[30] = 1'b0;
  assign io_ptw_ptbr_ppn[31] = 1'b0;
  assign io_ptw_ptbr_ppn[32] = 1'b0;
  assign io_ptw_ptbr_ppn[33] = 1'b0;
  assign io_ptw_ptbr_ppn[34] = 1'b0;
  assign io_ptw_ptbr_ppn[35] = 1'b0;
  assign io_ptw_ptbr_ppn[36] = 1'b0;
  assign io_ptw_ptbr_ppn[37] = 1'b0;
  assign io_ptw_ptbr_ppn[38] = 1'b0;
  assign io_ptw_ptbr_ppn[39] = 1'b0;
  assign io_ptw_ptbr_ppn[40] = 1'b0;
  assign io_ptw_ptbr_ppn[41] = 1'b0;
  assign io_ptw_ptbr_ppn[42] = 1'b0;
  assign io_ptw_ptbr_ppn[43] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[0] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[1] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[2] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[4] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[5] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[6] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[7] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[8] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[10] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[11] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[12] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[13] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[14] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[15] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[16] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[17] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[18] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[19] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[20] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[21] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[22] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[23] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[24] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[25] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[26] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[27] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[28] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[29] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[30] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[31] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[32] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[33] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[34] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[35] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[36] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[37] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[38] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[39] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[40] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[41] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[42] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[43] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[44] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[45] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[46] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[47] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[48] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[49] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[50] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[51] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[52] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[53] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[54] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[55] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[56] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[57] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[58] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[59] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[60] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[61] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[62] = 1'b0;
  assign io_ptw_customCSRs_csrs_0_value[63] = 1'b0;
  assign io_ptw_pmp_0_mask[1] = 1'b1;
  assign io_ptw_pmp_0_mask[0] = 1'b1;
  assign io_ptw_pmp_1_mask[1] = 1'b1;
  assign io_ptw_pmp_1_mask[0] = 1'b1;
  assign io_ptw_pmp_2_mask[1] = 1'b1;
  assign io_ptw_pmp_2_mask[0] = 1'b1;
  assign io_ptw_pmp_3_mask[1] = 1'b1;
  assign io_ptw_pmp_3_mask[0] = 1'b1;
  assign io_ptw_pmp_4_mask[1] = 1'b1;
  assign io_ptw_pmp_4_mask[0] = 1'b1;
  assign io_ptw_pmp_5_mask[1] = 1'b1;
  assign io_ptw_pmp_5_mask[0] = 1'b1;
  assign io_ptw_pmp_6_mask[1] = 1'b1;
  assign io_ptw_pmp_6_mask[0] = 1'b1;
  assign io_ptw_pmp_7_mask[1] = 1'b1;
  assign io_ptw_pmp_7_mask[0] = 1'b1;
  assign io_fpu_inst[1] = 1'b1;
  assign io_fpu_inst[0] = 1'b1;
  assign io_fpu_dmem_resp_type[1] = io_dmem_resp_bits_size[1];
  assign io_fpu_dmem_resp_type[0] = io_dmem_resp_bits_size[0];
  assign io_fpu_dmem_resp_tag[4] = io_dmem_resp_bits_tag[5];
  assign io_fpu_dmem_resp_tag[3] = io_dmem_resp_bits_tag[4];
  assign io_fpu_dmem_resp_tag[2] = io_dmem_resp_bits_tag[3];
  assign io_fpu_dmem_resp_tag[1] = io_dmem_resp_bits_tag[2];
  assign io_fpu_dmem_resp_tag[0] = io_dmem_resp_bits_tag[1];
  assign io_fpu_dmem_resp_data[63] = io_dmem_resp_bits_data_word_bypass[63];
  assign io_fpu_dmem_resp_data[62] = io_dmem_resp_bits_data_word_bypass[62];
  assign io_fpu_dmem_resp_data[61] = io_dmem_resp_bits_data_word_bypass[61];
  assign io_fpu_dmem_resp_data[60] = io_dmem_resp_bits_data_word_bypass[60];
  assign io_fpu_dmem_resp_data[59] = io_dmem_resp_bits_data_word_bypass[59];
  assign io_fpu_dmem_resp_data[58] = io_dmem_resp_bits_data_word_bypass[58];
  assign io_fpu_dmem_resp_data[57] = io_dmem_resp_bits_data_word_bypass[57];
  assign io_fpu_dmem_resp_data[56] = io_dmem_resp_bits_data_word_bypass[56];
  assign io_fpu_dmem_resp_data[55] = io_dmem_resp_bits_data_word_bypass[55];
  assign io_fpu_dmem_resp_data[54] = io_dmem_resp_bits_data_word_bypass[54];
  assign io_fpu_dmem_resp_data[53] = io_dmem_resp_bits_data_word_bypass[53];
  assign io_fpu_dmem_resp_data[52] = io_dmem_resp_bits_data_word_bypass[52];
  assign io_fpu_dmem_resp_data[51] = io_dmem_resp_bits_data_word_bypass[51];
  assign io_fpu_dmem_resp_data[50] = io_dmem_resp_bits_data_word_bypass[50];
  assign io_fpu_dmem_resp_data[49] = io_dmem_resp_bits_data_word_bypass[49];
  assign io_fpu_dmem_resp_data[48] = io_dmem_resp_bits_data_word_bypass[48];
  assign io_fpu_dmem_resp_data[47] = io_dmem_resp_bits_data_word_bypass[47];
  assign io_fpu_dmem_resp_data[46] = io_dmem_resp_bits_data_word_bypass[46];
  assign io_fpu_dmem_resp_data[45] = io_dmem_resp_bits_data_word_bypass[45];
  assign io_fpu_dmem_resp_data[44] = io_dmem_resp_bits_data_word_bypass[44];
  assign io_fpu_dmem_resp_data[43] = io_dmem_resp_bits_data_word_bypass[43];
  assign io_fpu_dmem_resp_data[42] = io_dmem_resp_bits_data_word_bypass[42];
  assign io_fpu_dmem_resp_data[41] = io_dmem_resp_bits_data_word_bypass[41];
  assign io_fpu_dmem_resp_data[40] = io_dmem_resp_bits_data_word_bypass[40];
  assign io_fpu_dmem_resp_data[39] = io_dmem_resp_bits_data_word_bypass[39];
  assign io_fpu_dmem_resp_data[38] = io_dmem_resp_bits_data_word_bypass[38];
  assign io_fpu_dmem_resp_data[37] = io_dmem_resp_bits_data_word_bypass[37];
  assign io_fpu_dmem_resp_data[36] = io_dmem_resp_bits_data_word_bypass[36];
  assign io_fpu_dmem_resp_data[35] = io_dmem_resp_bits_data_word_bypass[35];
  assign io_fpu_dmem_resp_data[34] = io_dmem_resp_bits_data_word_bypass[34];
  assign io_fpu_dmem_resp_data[33] = io_dmem_resp_bits_data_word_bypass[33];
  assign io_fpu_dmem_resp_data[32] = io_dmem_resp_bits_data_word_bypass[32];
  assign io_fpu_dmem_resp_data[31] = io_dmem_resp_bits_data_word_bypass[31];
  assign io_fpu_dmem_resp_data[30] = io_dmem_resp_bits_data_word_bypass[30];
  assign io_fpu_dmem_resp_data[29] = io_dmem_resp_bits_data_word_bypass[29];
  assign io_fpu_dmem_resp_data[28] = io_dmem_resp_bits_data_word_bypass[28];
  assign io_fpu_dmem_resp_data[27] = io_dmem_resp_bits_data_word_bypass[27];
  assign io_fpu_dmem_resp_data[26] = io_dmem_resp_bits_data_word_bypass[26];
  assign io_fpu_dmem_resp_data[25] = io_dmem_resp_bits_data_word_bypass[25];
  assign io_fpu_dmem_resp_data[24] = io_dmem_resp_bits_data_word_bypass[24];
  assign io_fpu_dmem_resp_data[23] = io_dmem_resp_bits_data_word_bypass[23];
  assign io_fpu_dmem_resp_data[22] = io_dmem_resp_bits_data_word_bypass[22];
  assign io_fpu_dmem_resp_data[21] = io_dmem_resp_bits_data_word_bypass[21];
  assign io_fpu_dmem_resp_data[20] = io_dmem_resp_bits_data_word_bypass[20];
  assign io_fpu_dmem_resp_data[19] = io_dmem_resp_bits_data_word_bypass[19];
  assign io_fpu_dmem_resp_data[18] = io_dmem_resp_bits_data_word_bypass[18];
  assign io_fpu_dmem_resp_data[17] = io_dmem_resp_bits_data_word_bypass[17];
  assign io_fpu_dmem_resp_data[16] = io_dmem_resp_bits_data_word_bypass[16];
  assign io_fpu_dmem_resp_data[15] = io_dmem_resp_bits_data_word_bypass[15];
  assign io_fpu_dmem_resp_data[14] = io_dmem_resp_bits_data_word_bypass[14];
  assign io_fpu_dmem_resp_data[13] = io_dmem_resp_bits_data_word_bypass[13];
  assign io_fpu_dmem_resp_data[12] = io_dmem_resp_bits_data_word_bypass[12];
  assign io_fpu_dmem_resp_data[11] = io_dmem_resp_bits_data_word_bypass[11];
  assign io_fpu_dmem_resp_data[10] = io_dmem_resp_bits_data_word_bypass[10];
  assign io_fpu_dmem_resp_data[9] = io_dmem_resp_bits_data_word_bypass[9];
  assign io_fpu_dmem_resp_data[8] = io_dmem_resp_bits_data_word_bypass[8];
  assign io_fpu_dmem_resp_data[7] = io_dmem_resp_bits_data_word_bypass[7];
  assign io_fpu_dmem_resp_data[6] = io_dmem_resp_bits_data_word_bypass[6];
  assign io_fpu_dmem_resp_data[5] = io_dmem_resp_bits_data_word_bypass[5];
  assign io_fpu_dmem_resp_data[4] = io_dmem_resp_bits_data_word_bypass[4];
  assign io_fpu_dmem_resp_data[3] = io_dmem_resp_bits_data_word_bypass[3];
  assign io_fpu_dmem_resp_data[2] = io_dmem_resp_bits_data_word_bypass[2];
  assign io_fpu_dmem_resp_data[1] = io_dmem_resp_bits_data_word_bypass[1];
  assign io_fpu_dmem_resp_data[0] = io_dmem_resp_bits_data_word_bypass[0];

  IBuf ibuf ( .clock(n3595), .reset(reset), .io_imem_ready(io_imem_resp_ready), 
        .io_imem_valid(io_imem_resp_valid), .io_imem_bits_btb_taken(
        io_imem_resp_bits_btb_taken), .io_imem_bits_btb_bridx(
        io_imem_resp_bits_btb_bridx), .io_imem_bits_btb_entry(
        io_imem_resp_bits_btb_entry), .io_imem_bits_btb_bht_history(
        io_imem_resp_bits_btb_bht_history), .io_imem_bits_pc(
        io_imem_resp_bits_pc), .io_imem_bits_data(io_imem_resp_bits_data), 
        .io_imem_bits_xcpt_pf_inst(io_imem_resp_bits_xcpt_pf_inst), 
        .io_imem_bits_xcpt_ae_inst(io_imem_resp_bits_xcpt_ae_inst), 
        .io_imem_bits_replay(io_imem_resp_bits_replay), .io_kill(
        io_imem_req_valid), .io_pc(ibuf_io_pc), .io_btb_resp_entry(
        ibuf_io_btb_resp_entry), .io_btb_resp_bht_history(
        ibuf_io_btb_resp_bht_history), .io_inst_0_ready(n1822), 
        .io_inst_0_valid(ibuf_io_inst_0_valid), .io_inst_0_bits_xcpt0_pf_inst(
        n_T_728[1]), .io_inst_0_bits_xcpt0_ae_inst(n_T_728[0]), 
        .io_inst_0_bits_xcpt1_pf_inst(n_T_726[1]), 
        .io_inst_0_bits_xcpt1_ae_inst(n_T_726[0]), .io_inst_0_bits_replay(
        ibuf_io_inst_0_bits_replay), .io_inst_0_bits_inst_bits({n9517, n9518, 
        n9519, n9520, n9521, io_fpu_inst[26], n9522, io_fpu_inst[24:15], n9523, 
        n9524, io_fpu_inst[12:7], n9525, n9526, n9527, n9528, n9529, 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}), 
        .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd), 
        .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1), 
        .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2), 
        .io_inst_0_bits_inst_rs3({n2494, SYNOPSYS_UNCONNECTED_3, n2674, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5}), .io_inst_0_bits_raw(
        {n2576, ibuf_io_inst_0_bits_raw}), .io_inst_0_bits_rvc(
        ibuf_io_inst_0_bits_rvc) );
  CSRFile csr ( .clock(n3785), .reset(reset), .io_ungated_clock(clock), 
        .io_interrupts_debug(io_interrupts_debug), .io_interrupts_mtip(
        io_interrupts_mtip), .io_interrupts_msip(io_interrupts_msip), 
        .io_interrupts_meip(io_interrupts_meip), .io_interrupts_seip(
        io_interrupts_seip), .io_rw_addr(csr_io_rw_addr), .io_rw_cmd({
        csr_io_rw_cmd_2_, wb_ctrl_csr[1:0]}), .io_rw_rdata(csr_io_rw_rdata), 
        .io_rw_wdata({n_T_1165, io_imem_sfence_bits_addr}), .io_decode_0_csr({
        n2576, ibuf_io_inst_0_bits_raw[30], n2674, 
        ibuf_io_inst_0_bits_raw[28:20]}), .io_decode_0_fp_illegal(
        csr_io_decode_0_fp_illegal), .io_decode_0_fp_csr(
        csr_io_decode_0_fp_csr), .io_decode_0_read_illegal(
        csr_io_decode_0_read_illegal), .io_decode_0_write_illegal(
        csr_io_decode_0_write_illegal), .io_decode_0_write_flush(
        csr_io_decode_0_write_flush), .io_decode_0_system_illegal(
        csr_io_decode_0_system_illegal), .io_csr_stall(csr_io_csr_stall), 
        .io_eret(csr_io_eret), .io_singleStep(csr_io_singleStep), 
        .io_status_wfi(io_wfi), .io_status_dprv(io_dmem_req_bits_dprv), 
        .io_status_prv(io_ptw_status_prv), .io_status_zero2({
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32}), .io_status_sxl({
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34}), .io_status_uxl({
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36}), .io_status_zero1({
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44}), .io_status_mxr(
        io_ptw_status_mxr), .io_status_sum(io_ptw_status_sum), .io_status_xs({
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46}), .io_status_fs({
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48}), .io_status_mpp({
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50}), .io_status_vs({
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52}), .io_ptbr_mode({
        io_ptw_ptbr_mode[3], SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55}), .io_ptbr_ppn({SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, io_ptw_ptbr_ppn[19:0]}), .io_evec({
        csr_io_evec, SYNOPSYS_UNCONNECTED_80}), .io_exception(csr_io_exception), .io_retire(csr_io_retire), .io_cause({wb_cause[63], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, wb_cause[3:0]}), .io_pc({
        csr_io_pc[39:1], 1'b0}), .io_tval(csr_io_tval), .io_time({
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, csr_io_time}), 
        .io_fcsr_rm(io_fpu_fcsr_rm), .io_fcsr_flags_valid(
        io_fpu_fcsr_flags_valid), .io_fcsr_flags_bits(io_fpu_fcsr_flags_bits), 
        .io_interrupt(csr_io_interrupt), .io_interrupt_cause({
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, 
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, 
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, 
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, 
        SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        csr_io_interrupt_cause}), .io_bp_0_control_action(
        csr_io_bp_0_control_action), .io_bp_0_control_tmatch(
        csr_io_bp_0_control_tmatch), .io_bp_0_control_m(csr_io_bp_0_control_m), 
        .io_bp_0_control_s(csr_io_bp_0_control_s), .io_bp_0_control_u(
        csr_io_bp_0_control_u), .io_bp_0_control_x(csr_io_bp_0_control_x), 
        .io_bp_0_control_w(csr_io_bp_0_control_w), .io_bp_0_control_r(
        csr_io_bp_0_control_r), .io_bp_0_address(csr_io_bp_0_address), 
        .io_pmp_0_cfg_l(io_ptw_pmp_0_cfg_l), .io_pmp_0_cfg_a(
        io_ptw_pmp_0_cfg_a), .io_pmp_0_cfg_x(io_ptw_pmp_0_cfg_x), 
        .io_pmp_0_cfg_w(io_ptw_pmp_0_cfg_w), .io_pmp_0_cfg_r(
        io_ptw_pmp_0_cfg_r), .io_pmp_0_addr(io_ptw_pmp_0_addr), 
        .io_pmp_0_mask({io_ptw_pmp_0_mask[31:2], SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174}), .io_pmp_1_cfg_l(io_ptw_pmp_1_cfg_l), 
        .io_pmp_1_cfg_a(io_ptw_pmp_1_cfg_a), .io_pmp_1_cfg_x(
        io_ptw_pmp_1_cfg_x), .io_pmp_1_cfg_w(io_ptw_pmp_1_cfg_w), 
        .io_pmp_1_cfg_r(io_ptw_pmp_1_cfg_r), .io_pmp_1_addr(io_ptw_pmp_1_addr), 
        .io_pmp_1_mask({io_ptw_pmp_1_mask[31:2], SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176}), .io_pmp_2_cfg_l(io_ptw_pmp_2_cfg_l), 
        .io_pmp_2_cfg_a(io_ptw_pmp_2_cfg_a), .io_pmp_2_cfg_x(
        io_ptw_pmp_2_cfg_x), .io_pmp_2_cfg_w(io_ptw_pmp_2_cfg_w), 
        .io_pmp_2_cfg_r(io_ptw_pmp_2_cfg_r), .io_pmp_2_addr(io_ptw_pmp_2_addr), 
        .io_pmp_2_mask({io_ptw_pmp_2_mask[31:2], SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178}), .io_pmp_3_cfg_l(io_ptw_pmp_3_cfg_l), 
        .io_pmp_3_cfg_a(io_ptw_pmp_3_cfg_a), .io_pmp_3_cfg_x(
        io_ptw_pmp_3_cfg_x), .io_pmp_3_cfg_w(io_ptw_pmp_3_cfg_w), 
        .io_pmp_3_cfg_r(io_ptw_pmp_3_cfg_r), .io_pmp_3_addr(io_ptw_pmp_3_addr), 
        .io_pmp_3_mask({io_ptw_pmp_3_mask[31:2], SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180}), .io_pmp_4_cfg_l(io_ptw_pmp_4_cfg_l), 
        .io_pmp_4_cfg_a(io_ptw_pmp_4_cfg_a), .io_pmp_4_cfg_x(
        io_ptw_pmp_4_cfg_x), .io_pmp_4_cfg_w(io_ptw_pmp_4_cfg_w), 
        .io_pmp_4_cfg_r(io_ptw_pmp_4_cfg_r), .io_pmp_4_addr(io_ptw_pmp_4_addr), 
        .io_pmp_4_mask({io_ptw_pmp_4_mask[31:2], SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182}), .io_pmp_5_cfg_l(io_ptw_pmp_5_cfg_l), 
        .io_pmp_5_cfg_a(io_ptw_pmp_5_cfg_a), .io_pmp_5_cfg_x(
        io_ptw_pmp_5_cfg_x), .io_pmp_5_cfg_w(io_ptw_pmp_5_cfg_w), 
        .io_pmp_5_cfg_r(io_ptw_pmp_5_cfg_r), .io_pmp_5_addr(io_ptw_pmp_5_addr), 
        .io_pmp_5_mask({io_ptw_pmp_5_mask[31:2], SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184}), .io_pmp_6_cfg_l(io_ptw_pmp_6_cfg_l), 
        .io_pmp_6_cfg_a(io_ptw_pmp_6_cfg_a), .io_pmp_6_cfg_x(
        io_ptw_pmp_6_cfg_x), .io_pmp_6_cfg_w(io_ptw_pmp_6_cfg_w), 
        .io_pmp_6_cfg_r(io_ptw_pmp_6_cfg_r), .io_pmp_6_addr(io_ptw_pmp_6_addr), 
        .io_pmp_6_mask({io_ptw_pmp_6_mask[31:2], SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186}), .io_pmp_7_cfg_l(io_ptw_pmp_7_cfg_l), 
        .io_pmp_7_cfg_a(io_ptw_pmp_7_cfg_a), .io_pmp_7_cfg_x(
        io_ptw_pmp_7_cfg_x), .io_pmp_7_cfg_w(io_ptw_pmp_7_cfg_w), 
        .io_pmp_7_cfg_r(io_ptw_pmp_7_cfg_r), .io_pmp_7_addr(io_ptw_pmp_7_addr), 
        .io_pmp_7_mask({io_ptw_pmp_7_mask[31:2], SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188}), .io_inst_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .io_trace_0_iaddr({SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228}), .io_trace_0_insn({SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260}), .io_customCSRs_0_value({
        SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262, 
        SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, 
        SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, 
        SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, 
        SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, 
        io_ptw_customCSRs_csrs_0_value[9], SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        io_ptw_customCSRs_csrs_0_value[3], SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322}), 
        .io_status_debug_BAR(n9516), .io_status_isa_12__BAR(
        csr_io_status_isa[12]), .io_status_isa_3_(csr_io_status_isa[3]), 
        .io_status_isa_2_(csr_io_status_isa[2]), .io_status_isa_0__BAR(
        csr_io_status_isa[0]) );
  BreakpointUnit bpu ( .io_status_prv(io_ptw_status_prv), 
        .io_bp_0_control_action(csr_io_bp_0_control_action), 
        .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch), 
        .io_bp_0_control_m(csr_io_bp_0_control_m), .io_bp_0_control_s(
        csr_io_bp_0_control_s), .io_bp_0_control_u(csr_io_bp_0_control_u), 
        .io_bp_0_control_x(csr_io_bp_0_control_x), .io_bp_0_control_w(
        csr_io_bp_0_control_w), .io_bp_0_control_r(csr_io_bp_0_control_r), 
        .io_bp_0_address(csr_io_bp_0_address), .io_pc(ibuf_io_pc[38:0]), 
        .io_ea(n_T_918[38:0]), .io_xcpt_if(bpu_io_xcpt_if), .io_xcpt_ld(
        bpu_io_xcpt_ld), .io_xcpt_st(bpu_io_xcpt_st), .io_debug_if(
        bpu_io_debug_if), .io_debug_ld(bpu_io_debug_ld), .io_debug_st(
        bpu_io_debug_st), .io_status_debug_BAR(n9516) );
  ALU alu ( .io_dw(alu_io_dw), .io_fn(alu_io_fn), .io_in2(alu_io_in2), 
        .io_in1(alu_io_in1), .io_out(alu_io_out), .io_adder_out({
        SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, 
        SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, 
        SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, 
        SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, 
        SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        alu_io_adder_out_39_, io_dmem_req_bits_addr[38:0]}), .io_cmp_out(
        alu_io_cmp_out) );
  MulDiv div ( .clock(n3785), .reset(reset), .io_req_ready(div_io_req_ready), 
        .io_req_valid(n9422), .io_req_bits_fn({1'b0, alu_io_fn[2:0]}), 
        .io_req_bits_dw(alu_io_dw), .io_req_bits_in1(io_fpu_fromint_data), 
        .io_req_bits_in2(n_T_702), .io_req_bits_tag(io_dmem_req_bits_tag[5:1]), 
        .io_kill(div_io_kill), .io_resp_ready(div_io_resp_ready), 
        .io_resp_valid(div_io_resp_valid), .io_resp_bits_data(
        div_io_resp_bits_data), .io_resp_bits_tag_4__BAR(
        div_io_resp_bits_tag[4]), .io_resp_bits_tag_2_(div_io_resp_bits_tag[2]), .io_resp_bits_tag_0_(div_io_resp_bits_tag[0]), .io_resp_bits_tag_3__BAR(
        div_io_resp_bits_tag[3]), .io_resp_bits_tag_1__BAR(
        div_io_resp_bits_tag[1]) );
  PlusArgTimeout PlusArgTimeout ( .clock(n3595), .reset(reset), .io_count(
        csr_io_time) );
  SNPS_CLOCK_GATE_HIGH_Rocket_0 clk_gate_ex_reg_rs_bypass_1_reg ( .CLK(n3595), 
        .EN(n406), .ENCLK(net34469), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_39 clk_gate_wb_ctrl_wxd_reg ( .CLK(n4499), .EN(
        mem_pc_valid), .ENCLK(net34475), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_38 clk_gate_mem_ctrl_branch_reg ( .CLK(n4499), 
        .EN(N290), .ENCLK(net34480), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_37 clk_gate__T_427_reg_0_ ( .CLK(n3595), .EN(
        N268), .ENCLK(net34485), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_36 clk_gate__T_427_reg_1_ ( .CLK(n3595), .EN(
        N267), .ENCLK(net34490), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_35 clk_gate__T_427_reg_2_ ( .CLK(n3595), .EN(
        N266), .ENCLK(net34495), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_34 clk_gate__T_427_reg_3_ ( .CLK(n3595), .EN(
        N265), .ENCLK(net34500), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_33 clk_gate__T_427_reg_4_ ( .CLK(n3595), .EN(
        N264), .ENCLK(net34505), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_32 clk_gate__T_427_reg_5_ ( .CLK(n3595), .EN(
        N263), .ENCLK(net34510), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_31 clk_gate__T_427_reg_6_ ( .CLK(n3595), .EN(
        N262), .ENCLK(net34515), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_30 clk_gate__T_427_reg_7_ ( .CLK(n3785), .EN(
        N261), .ENCLK(net34520), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_29 clk_gate__T_427_reg_8_ ( .CLK(n3594), .EN(
        N260), .ENCLK(net34525), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_28 clk_gate__T_427_reg_9_ ( .CLK(n3785), .EN(
        N259), .ENCLK(net34530), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_27 clk_gate__T_427_reg_10_ ( .CLK(n4499), .EN(
        N258), .ENCLK(net34535), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_26 clk_gate__T_427_reg_11_ ( .CLK(n3785), .EN(
        N257), .ENCLK(net34540), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_25 clk_gate__T_427_reg_12_ ( .CLK(n4499), .EN(
        N256), .ENCLK(net34545), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_24 clk_gate__T_427_reg_13_ ( .CLK(n3785), .EN(
        N255), .ENCLK(net34550), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_23 clk_gate__T_427_reg_14_ ( .CLK(n4499), .EN(
        N254), .ENCLK(net34555), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_22 clk_gate__T_427_reg_15_ ( .CLK(n3785), .EN(
        N253), .ENCLK(net34560), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_21 clk_gate__T_427_reg_16_ ( .CLK(n4499), .EN(
        N252), .ENCLK(net34565), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_20 clk_gate__T_427_reg_17_ ( .CLK(n3595), .EN(
        N251), .ENCLK(net34570), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_19 clk_gate__T_427_reg_18_ ( .CLK(n3594), .EN(
        N250), .ENCLK(net34575), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_18 clk_gate__T_427_reg_19_ ( .CLK(n3785), .EN(
        N249), .ENCLK(net34580), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_17 clk_gate__T_427_reg_20_ ( .CLK(n4499), .EN(
        N248), .ENCLK(net34585), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_16 clk_gate__T_427_reg_21_ ( .CLK(n3785), .EN(
        N247), .ENCLK(net34590), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_15 clk_gate__T_427_reg_22_ ( .CLK(n4499), .EN(
        N246), .ENCLK(net34595), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_14 clk_gate__T_427_reg_23_ ( .CLK(n3785), .EN(
        N245), .ENCLK(net34600), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_13 clk_gate__T_427_reg_24_ ( .CLK(n4499), .EN(
        N244), .ENCLK(net34605), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_12 clk_gate__T_427_reg_25_ ( .CLK(n3785), .EN(
        N243), .ENCLK(net34610), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_11 clk_gate__T_427_reg_26_ ( .CLK(n4499), .EN(
        N242), .ENCLK(net34615), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_10 clk_gate__T_427_reg_27_ ( .CLK(n3785), .EN(
        N241), .ENCLK(net34620), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_9 clk_gate__T_427_reg_28_ ( .CLK(n4499), .EN(
        N240), .ENCLK(net34625), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_8 clk_gate__T_427_reg_29_ ( .CLK(n3785), .EN(
        N239), .ENCLK(net34630), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_7 clk_gate__T_427_reg_30_ ( .CLK(n4499), .EN(
        N238), .ENCLK(net34635), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_6 clk_gate_ex_reg_btb_resp_bht_history_reg ( 
        .CLK(n3785), .EN(n_T_760), .ENCLK(net34640), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_5 clk_gate_mem_reg_rs2_reg ( .CLK(n4499), .EN(
        N526), .ENCLK(net34645), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_4 clk_gate_ex_reg_rs_msb_0_reg ( .CLK(n3594), 
        .EN(N744), .ENCLK(net34650), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_3 clk_gate_ex_reg_rs_msb_1_reg ( .CLK(n3785), 
        .EN(N745), .ENCLK(net34655), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_2 clk_gate__T_1185_reg ( .CLK(clock), .EN(N746), 
        .ENCLK(net34660), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Rocket_1 clk_gate__T_1298_reg ( .CLK(n3595), .EN(N778), 
        .ENCLK(net34665), .TE(1'b0) );
  Rocket_DW01_add_J37_0 add_x_94 ( .A(mem_reg_pc[38:0]), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n570, 1'b0}), .CI(1'b0), .SUM(io_imem_btb_update_bits_br_pc) );
  Rocket_DW01_add_J37_1 add_x_5 ( .A(mem_reg_pc), .B({n9427, n9427, n9427, 
        n9427, n9427, n9427, n9427, n9427, n9427, n9427, n9427, n9427, n9427, 
        n9427, n9427, n9427, n9427, n9427, n9427, n9427, n_T_914, 1'b0}), .CI(
        1'b0), .SUM(mem_br_target) );
  DFFX1_LVT mem_reg_inst_reg_7_ ( .D(n592), .CLK(n4286), .Q(n3202), .QN(
        n_T_849[11]) );
  DFFX1_LVT ex_reg_valid_reg ( .D(n2874), .CLK(n3594), .QN(ex_reg_valid) );
  DFFX1_LVT mem_reg_valid_reg ( .D(io_fpu_killx), .CLK(n3594), .Q(n3206), .QN(
        mem_reg_valid) );
  DFFX1_LVT wb_reg_wdata_reg_0_ ( .D(N598), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[0]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_61_ ( .D(id_rs_1[63]), .CLK(n4079), .Q(
        n_T_635[63]) );
  DFFX1_LVT mem_reg_wdata_reg_63_ ( .D(alu_io_out[63]), .CLK(n4293), .Q(
        n_T_918[63]) );
  DFFSSRX1_LVT mem_reg_replay_reg ( .D(n9421), .SETB(n9418), .RSTB(1'b1), 
        .CLK(n3594), .QN(mem_reg_replay) );
  DFFX1_LVT wb_reg_replay_reg ( .D(N530), .CLK(n3594), .Q(wb_reg_replay) );
  DFFX1_LVT ex_ctrl_sel_imm_reg_1_ ( .D(id_ctrl_sel_imm[1]), .CLK(n4312), .QN(
        n546) );
  DFFX1_LVT ex_ctrl_mem_cmd_reg_4_ ( .D(n1891), .CLK(n4315), .Q(
        io_dmem_req_bits_cmd[4]), .QN(n3245) );
  DFFX1_LVT ex_ctrl_jal_reg ( .D(n9428), .CLK(n4315), .Q(ex_ctrl_jal) );
  DFFX1_LVT ex_ctrl_branch_reg ( .D(n9429), .CLK(n4315), .QN(n323) );
  DFFX1_LVT ex_ctrl_sel_imm_reg_0_ ( .D(id_ctrl_sel_imm[0]), .CLK(n4315), .Q(
        ex_ctrl_sel_imm[0]) );
  DFFX1_LVT ex_ctrl_csr_reg_0_ ( .D(N286), .CLK(n4315), .Q(ex_ctrl_csr[0]), 
        .QN(n320) );
  DFFX1_LVT ex_ctrl_csr_reg_1_ ( .D(n1628), .CLK(n4314), .Q(n319), .QN(
        ex_ctrl_csr[1]) );
  DFFX1_LVT ex_ctrl_fence_i_reg ( .D(n1828), .CLK(n4314), .QN(n318) );
  DFFX1_LVT ex_ctrl_sel_imm_reg_2_ ( .D(id_ctrl_sel_imm[2]), .CLK(n4314), .Q(
        ex_ctrl_sel_imm[2]), .QN(n3231) );
  DFFX1_LVT ex_ctrl_jalr_reg ( .D(n1823), .CLK(n4314), .Q(ex_ctrl_jalr), .QN(
        n2495) );
  DFFX1_LVT id_reg_pause_reg ( .D(n1820), .CLK(n3594), .Q(id_reg_pause) );
  DFFX1_LVT ex_ctrl_div_reg ( .D(n9413), .CLK(n4314), .Q(n317), .QN(
        ex_ctrl_div) );
  DFFX1_LVT ex_ctrl_mem_cmd_reg_0_ ( .D(n9431), .CLK(n4314), .Q(
        io_dmem_req_bits_cmd[0]), .QN(n560) );
  DFFSSRX1_LVT ex_ctrl_rxs2_reg ( .D(n1531), .SETB(1'b1), .RSTB(n1532), .CLK(
        n4312), .QN(ex_ctrl_rxs2) );
  DFFX1_LVT ex_ctrl_wfd_reg ( .D(id_ctrl_wfd), .CLK(n4314), .Q(ex_ctrl_wfd), 
        .QN(n315) );
  DFFX1_LVT ex_ctrl_wxd_reg ( .D(id_ctrl_wxd), .CLK(n4314), .Q(ex_ctrl_wxd), 
        .QN(n314) );
  DFFX1_LVT ex_ctrl_mem_cmd_reg_2_ ( .D(id_ctrl_mem_cmd_2_), .CLK(n4314), .Q(
        io_dmem_req_bits_cmd[2]), .QN(n3244) );
  DFFX1_LVT ex_reg_mem_size_reg_0_ ( .D(N369), .CLK(n4314), .Q(
        io_dmem_req_bits_size[0]), .QN(n313) );
  DFFX1_LVT id_reg_fence_reg ( .D(n1821), .CLK(n3595), .Q(id_reg_fence) );
  DFFX1_LVT blocked_reg ( .D(N811), .CLK(n3594), .Q(blocked) );
  DFFSSRX1_LVT ex_ctrl_csr_reg_2_ ( .D(n1628), .SETB(n2569), .RSTB(n2131), 
        .CLK(n4312), .Q(ex_ctrl_csr[2]), .QN(n310) );
  DFFX1_LVT ex_reg_flush_pipe_reg ( .D(n_T_731), .CLK(n4313), .QN(n309) );
  DFFX1_LVT ex_reg_inst_reg_31_ ( .D(n9434), .CLK(n4098), .Q(n172), .QN(
        ex_reg_inst_31_) );
  DFFX1_LVT ex_reg_inst_reg_30_ ( .D(n9435), .CLK(n4098), .Q(n171), .QN(
        n_T_642[10]) );
  DFFX1_LVT ex_reg_inst_reg_29_ ( .D(n9436), .CLK(n4098), .Q(n170), .QN(
        n_T_642[9]) );
  DFFX1_LVT ex_reg_inst_reg_28_ ( .D(n9437), .CLK(n4098), .Q(n169), .QN(
        n_T_642[8]) );
  DFFX1_LVT ex_reg_inst_reg_27_ ( .D(n9438), .CLK(n4098), .Q(n168), .QN(
        n_T_642[7]) );
  DFFX1_LVT ex_reg_inst_reg_26_ ( .D(n9439), .CLK(n4098), .Q(n167), .QN(
        n_T_642[6]) );
  DFFX1_LVT ex_reg_inst_reg_25_ ( .D(n9440), .CLK(n4098), .Q(n166), .QN(
        n_T_642[5]) );
  DFFX1_LVT ex_reg_inst_reg_24_ ( .D(io_fpu_inst[24]), .CLK(n4098), .Q(
        n_T_642[4]), .QN(n165) );
  DFFX1_LVT ex_reg_inst_reg_23_ ( .D(n9441), .CLK(n4098), .Q(n164), .QN(
        n_T_642[3]) );
  DFFX1_LVT ex_reg_inst_reg_22_ ( .D(n9442), .CLK(n4098), .Q(n163), .QN(
        n_T_642[2]) );
  DFFX1_LVT ex_reg_inst_reg_21_ ( .D(n9443), .CLK(n4098), .Q(n162), .QN(
        n_T_642[1]) );
  DFFX1_LVT ex_reg_inst_reg_20_ ( .D(n9444), .CLK(n4097), .Q(n161), .QN(
        n_T_642[0]) );
  DFFX1_LVT ex_reg_inst_reg_19_ ( .D(io_fpu_inst[19]), .CLK(n4097), .Q(
        n_T_648[7]), .QN(n160) );
  DFFX1_LVT ex_reg_inst_reg_18_ ( .D(io_fpu_inst[18]), .CLK(n4097), .Q(
        n_T_648[6]), .QN(n159) );
  DFFX1_LVT ex_reg_inst_reg_17_ ( .D(io_fpu_inst[17]), .CLK(n4097), .Q(
        n_T_648[5]), .QN(n158) );
  DFFX1_LVT ex_reg_inst_reg_16_ ( .D(io_fpu_inst[16]), .CLK(n4097), .Q(
        n_T_648[4]), .QN(n157) );
  DFFX1_LVT ex_reg_inst_reg_15_ ( .D(io_fpu_inst[15]), .CLK(n4097), .Q(
        n_T_648[3]), .QN(n156) );
  DFFX1_LVT ex_reg_inst_reg_14_ ( .D(n9445), .CLK(n4097), .Q(
        io_dmem_req_bits_signed), .QN(n_T_648[2]) );
  DFFX1_LVT ex_reg_inst_reg_13_ ( .D(n9446), .CLK(n4097), .Q(n155), .QN(
        n_T_648[1]) );
  DFFX1_LVT ex_reg_inst_reg_12_ ( .D(n3583), .CLK(n4097), .Q(n154), .QN(
        n_T_648[0]) );
  DFFX1_LVT ex_reg_inst_reg_11_ ( .D(io_fpu_inst[11]), .CLK(n4097), .Q(
        io_dmem_req_bits_tag[5]), .QN(n588) );
  DFFX1_LVT ex_reg_inst_reg_10_ ( .D(n9447), .CLK(n4097), .Q(n589), .QN(
        io_dmem_req_bits_tag[4]) );
  DFFX1_LVT ex_reg_inst_reg_9_ ( .D(io_fpu_inst[9]), .CLK(n4097), .Q(
        io_dmem_req_bits_tag[3]), .QN(n590) );
  DFFX1_LVT ex_reg_inst_reg_8_ ( .D(io_fpu_inst[8]), .CLK(n4096), .Q(
        io_dmem_req_bits_tag[2]), .QN(n591) );
  DFFX1_LVT ex_reg_inst_reg_7_ ( .D(io_fpu_inst[7]), .CLK(n4096), .Q(
        io_dmem_req_bits_tag[1]), .QN(n592) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_0_ ( .D(
        ibuf_io_btb_resp_bht_history[0]), .CLK(n4096), .QN(n152) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_1_ ( .D(
        ibuf_io_btb_resp_bht_history[1]), .CLK(n4096), .QN(n151) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_2_ ( .D(
        ibuf_io_btb_resp_bht_history[2]), .CLK(n4096), .QN(n150) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_3_ ( .D(
        ibuf_io_btb_resp_bht_history[3]), .CLK(n4096), .QN(n149) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_4_ ( .D(
        ibuf_io_btb_resp_bht_history[4]), .CLK(n4096), .QN(n148) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_5_ ( .D(
        ibuf_io_btb_resp_bht_history[5]), .CLK(n4096), .QN(n147) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_6_ ( .D(
        ibuf_io_btb_resp_bht_history[6]), .CLK(n4096), .QN(n146) );
  DFFX1_LVT ex_reg_btb_resp_bht_history_reg_7_ ( .D(
        ibuf_io_btb_resp_bht_history[7]), .CLK(n4096), .QN(n145) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_0_ ( .D(ibuf_io_btb_resp_entry[0]), 
        .CLK(n4096), .QN(n144) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_1_ ( .D(ibuf_io_btb_resp_entry[1]), 
        .CLK(n4096), .QN(n143) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_2_ ( .D(ibuf_io_btb_resp_entry[2]), 
        .CLK(n4095), .QN(n142) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_3_ ( .D(ibuf_io_btb_resp_entry[3]), 
        .CLK(n4095), .QN(n141) );
  DFFX1_LVT ex_reg_btb_resp_entry_reg_4_ ( .D(ibuf_io_btb_resp_entry[4]), 
        .CLK(n4095), .QN(n140) );
  DFFX1_LVT ex_reg_pc_reg_0_ ( .D(ibuf_io_pc[0]), .CLK(n4095), .Q(n_T_698[0]), 
        .QN(n139) );
  DFFX1_LVT ex_reg_pc_reg_1_ ( .D(ibuf_io_pc[1]), .CLK(n4095), .Q(n_T_698[1]), 
        .QN(n138) );
  DFFX1_LVT ex_reg_pc_reg_2_ ( .D(ibuf_io_pc[2]), .CLK(n4095), .Q(n_T_698[2]), 
        .QN(n137) );
  DFFX1_LVT ex_reg_pc_reg_3_ ( .D(ibuf_io_pc[3]), .CLK(n4095), .Q(n_T_698[3]), 
        .QN(n136) );
  DFFX1_LVT ex_reg_pc_reg_4_ ( .D(ibuf_io_pc[4]), .CLK(n4095), .Q(n_T_698[4]), 
        .QN(n135) );
  DFFX1_LVT ex_reg_pc_reg_5_ ( .D(ibuf_io_pc[5]), .CLK(n4095), .Q(n_T_698[5]), 
        .QN(n134) );
  DFFX1_LVT ex_reg_pc_reg_6_ ( .D(ibuf_io_pc[6]), .CLK(n4095), .Q(n_T_698[6]), 
        .QN(n133) );
  DFFX1_LVT ex_reg_pc_reg_7_ ( .D(ibuf_io_pc[7]), .CLK(n4095), .Q(n_T_698[7]), 
        .QN(n132) );
  DFFX1_LVT ex_reg_pc_reg_8_ ( .D(ibuf_io_pc[8]), .CLK(n4095), .Q(n_T_698[8]), 
        .QN(n131) );
  DFFX1_LVT ex_reg_pc_reg_9_ ( .D(ibuf_io_pc[9]), .CLK(n4094), .Q(n_T_698[9]), 
        .QN(n130) );
  DFFX1_LVT ex_reg_pc_reg_10_ ( .D(ibuf_io_pc[10]), .CLK(n4094), .Q(
        n_T_698[10]), .QN(n129) );
  DFFX1_LVT ex_reg_pc_reg_11_ ( .D(ibuf_io_pc[11]), .CLK(n4094), .Q(
        n_T_698[11]), .QN(n128) );
  DFFX1_LVT ex_reg_pc_reg_12_ ( .D(ibuf_io_pc[12]), .CLK(n4094), .Q(
        n_T_698[12]), .QN(n127) );
  DFFX1_LVT ex_reg_pc_reg_13_ ( .D(ibuf_io_pc[13]), .CLK(n4094), .Q(
        n_T_698[13]), .QN(n126) );
  DFFX1_LVT ex_reg_pc_reg_14_ ( .D(ibuf_io_pc[14]), .CLK(n4094), .Q(
        n_T_698[14]), .QN(n125) );
  DFFX1_LVT ex_reg_pc_reg_15_ ( .D(ibuf_io_pc[15]), .CLK(n4094), .Q(
        n_T_698[15]), .QN(n124) );
  DFFX1_LVT ex_reg_pc_reg_16_ ( .D(ibuf_io_pc[16]), .CLK(n4094), .Q(
        n_T_698[16]), .QN(n123) );
  DFFX1_LVT ex_reg_pc_reg_17_ ( .D(ibuf_io_pc[17]), .CLK(n4094), .Q(
        n_T_698[17]), .QN(n122) );
  DFFX1_LVT ex_reg_pc_reg_18_ ( .D(ibuf_io_pc[18]), .CLK(n4094), .Q(
        n_T_698[18]), .QN(n121) );
  DFFX1_LVT ex_reg_pc_reg_19_ ( .D(ibuf_io_pc[19]), .CLK(n4094), .Q(
        n_T_698[19]), .QN(n120) );
  DFFX1_LVT ex_reg_pc_reg_20_ ( .D(ibuf_io_pc[20]), .CLK(n4094), .Q(
        n_T_698[20]), .QN(n119) );
  DFFX1_LVT ex_reg_pc_reg_21_ ( .D(ibuf_io_pc[21]), .CLK(n4093), .Q(
        n_T_698[21]), .QN(n118) );
  DFFX1_LVT ex_reg_pc_reg_22_ ( .D(ibuf_io_pc[22]), .CLK(n4093), .Q(
        n_T_698[22]), .QN(n117) );
  DFFX1_LVT ex_reg_pc_reg_23_ ( .D(ibuf_io_pc[23]), .CLK(n4093), .Q(
        n_T_698[23]), .QN(n116) );
  DFFX1_LVT ex_reg_pc_reg_24_ ( .D(ibuf_io_pc[24]), .CLK(n4093), .Q(
        n_T_698[24]), .QN(n115) );
  DFFX1_LVT ex_reg_pc_reg_25_ ( .D(ibuf_io_pc[25]), .CLK(n4093), .Q(
        n_T_698[25]), .QN(n114) );
  DFFX1_LVT ex_reg_pc_reg_26_ ( .D(ibuf_io_pc[26]), .CLK(n4093), .Q(
        n_T_698[26]), .QN(n113) );
  DFFX1_LVT ex_reg_pc_reg_27_ ( .D(ibuf_io_pc[27]), .CLK(n4093), .Q(
        n_T_698[27]), .QN(n112) );
  DFFX1_LVT ex_reg_pc_reg_28_ ( .D(ibuf_io_pc[28]), .CLK(n4093), .Q(
        n_T_698[28]), .QN(n111) );
  DFFX1_LVT ex_reg_pc_reg_29_ ( .D(ibuf_io_pc[29]), .CLK(n4093), .Q(
        n_T_698[29]), .QN(n110) );
  DFFX1_LVT ex_reg_pc_reg_30_ ( .D(ibuf_io_pc[30]), .CLK(n4093), .Q(
        n_T_698[30]), .QN(n109) );
  DFFX1_LVT ex_reg_pc_reg_31_ ( .D(ibuf_io_pc[31]), .CLK(n4093), .Q(
        n_T_698[31]), .QN(n108) );
  DFFX1_LVT ex_reg_pc_reg_32_ ( .D(ibuf_io_pc[32]), .CLK(n4093), .Q(
        n_T_698[32]), .QN(n107) );
  DFFX1_LVT ex_reg_pc_reg_33_ ( .D(ibuf_io_pc[33]), .CLK(n4092), .Q(
        n_T_698[33]), .QN(n106) );
  DFFX1_LVT ex_reg_pc_reg_34_ ( .D(ibuf_io_pc[34]), .CLK(n4092), .Q(
        n_T_698[34]), .QN(n105) );
  DFFX1_LVT ex_reg_pc_reg_35_ ( .D(ibuf_io_pc[35]), .CLK(n4092), .Q(
        n_T_698[35]), .QN(n104) );
  DFFX1_LVT ex_reg_pc_reg_36_ ( .D(ibuf_io_pc[36]), .CLK(n4092), .Q(
        n_T_698[36]), .QN(n103) );
  DFFX1_LVT ex_reg_pc_reg_37_ ( .D(ibuf_io_pc[37]), .CLK(n4092), .Q(
        n_T_698[37]), .QN(n102) );
  DFFX1_LVT ex_reg_pc_reg_38_ ( .D(ibuf_io_pc[38]), .CLK(n4092), .Q(
        n_T_698[38]), .QN(n101) );
  DFFX1_LVT ex_reg_pc_reg_39_ ( .D(ibuf_io_pc[39]), .CLK(n4092), .Q(
        n_T_698[39]), .QN(n100) );
  DFFSSRX1_LVT ex_reg_replay_reg ( .D(n9433), .SETB(n9417), .RSTB(1'b1), .CLK(
        n3594), .Q(n3233), .QN(ex_reg_replay) );
  DFFSSRX1_LVT ex_reg_xcpt_interrupt_reg ( .D(n9448), .SETB(n9417), .RSTB(1'b1), .CLK(n3594), .Q(n98), .QN(ex_reg_xcpt_interrupt) );
  DFFX1_LVT mem_ctrl_branch_reg ( .D(n323), .CLK(n4286), .QN(
        io_imem_bht_update_bits_branch) );
  DFFX1_LVT mem_ctrl_fp_reg ( .D(n322), .CLK(n4286), .Q(n3246), .QN(n2492) );
  DFFX1_LVT mem_ctrl_jalr_reg ( .D(ex_ctrl_jalr), .CLK(n4286), .Q(
        mem_ctrl_jalr), .QN(n3104) );
  DFFX1_LVT mem_reg_wdata_reg_62_ ( .D(alu_io_out[62]), .CLK(n4286), .Q(
        n_T_918[62]) );
  DFFX1_LVT mem_reg_wdata_reg_61_ ( .D(alu_io_out[61]), .CLK(n4286), .Q(
        n_T_918[61]) );
  DFFX1_LVT mem_reg_wdata_reg_60_ ( .D(alu_io_out[60]), .CLK(n4286), .Q(
        n_T_918[60]) );
  DFFX1_LVT mem_reg_wdata_reg_59_ ( .D(alu_io_out[59]), .CLK(n4287), .Q(
        n_T_918[59]) );
  DFFX1_LVT mem_reg_wdata_reg_58_ ( .D(alu_io_out[58]), .CLK(n4287), .Q(
        n_T_918[58]) );
  DFFX1_LVT mem_reg_wdata_reg_57_ ( .D(alu_io_out[57]), .CLK(n4287), .Q(
        n_T_918[57]) );
  DFFX1_LVT mem_reg_wdata_reg_56_ ( .D(alu_io_out[56]), .CLK(n4287), .Q(
        n_T_918[56]) );
  DFFX1_LVT mem_reg_wdata_reg_55_ ( .D(alu_io_out[55]), .CLK(n4287), .Q(
        n_T_918[55]) );
  DFFX1_LVT mem_reg_wdata_reg_54_ ( .D(alu_io_out[54]), .CLK(n4287), .Q(
        n_T_918[54]) );
  DFFX1_LVT mem_reg_wdata_reg_53_ ( .D(alu_io_out[53]), .CLK(n4287), .Q(
        n_T_918[53]) );
  DFFX1_LVT mem_reg_wdata_reg_52_ ( .D(alu_io_out[52]), .CLK(n4287), .Q(
        n_T_918[52]) );
  DFFX1_LVT mem_reg_wdata_reg_51_ ( .D(alu_io_out[51]), .CLK(n4288), .Q(
        n_T_918[51]), .QN(n3249) );
  DFFX1_LVT mem_reg_wdata_reg_50_ ( .D(alu_io_out[50]), .CLK(n4287), .Q(
        n_T_918[50]) );
  DFFX1_LVT mem_reg_wdata_reg_49_ ( .D(alu_io_out[49]), .CLK(n4287), .Q(
        n_T_918[49]) );
  DFFX1_LVT mem_reg_wdata_reg_48_ ( .D(alu_io_out[48]), .CLK(n4287), .Q(
        n_T_918[48]) );
  DFFX1_LVT mem_reg_wdata_reg_47_ ( .D(alu_io_out[47]), .CLK(n4288), .Q(
        n_T_918[47]) );
  DFFX1_LVT mem_reg_wdata_reg_46_ ( .D(alu_io_out[46]), .CLK(n4287), .Q(
        n_T_918[46]) );
  DFFX1_LVT mem_reg_wdata_reg_45_ ( .D(alu_io_out[45]), .CLK(n4288), .Q(
        n_T_918[45]) );
  DFFX1_LVT mem_reg_wdata_reg_44_ ( .D(alu_io_out[44]), .CLK(n4288), .Q(
        n_T_918[44]) );
  DFFX1_LVT mem_reg_wdata_reg_43_ ( .D(alu_io_out[43]), .CLK(n4288), .Q(
        n_T_918[43]) );
  DFFX1_LVT mem_reg_wdata_reg_42_ ( .D(alu_io_out[42]), .CLK(n4288), .Q(
        n_T_918[42]) );
  DFFX1_LVT mem_reg_wdata_reg_41_ ( .D(alu_io_out[41]), .CLK(n4288), .Q(
        n_T_918[41]) );
  DFFX1_LVT mem_reg_wdata_reg_40_ ( .D(alu_io_out[40]), .CLK(n4288), .Q(
        n_T_918[40]) );
  DFFX1_LVT mem_reg_wdata_reg_39_ ( .D(alu_io_out[39]), .CLK(n4288), .Q(
        n_T_918[39]) );
  DFFX1_LVT mem_reg_wdata_reg_38_ ( .D(alu_io_out[38]), .CLK(n4288), .Q(
        n_T_918[38]), .QN(n3205) );
  DFFX1_LVT mem_reg_wdata_reg_37_ ( .D(alu_io_out[37]), .CLK(n4289), .Q(
        n_T_918[37]), .QN(n3528) );
  DFFX1_LVT mem_reg_wdata_reg_36_ ( .D(alu_io_out[36]), .CLK(n4288), .Q(
        n_T_918[36]), .QN(n3227) );
  DFFX1_LVT mem_reg_wdata_reg_35_ ( .D(alu_io_out[35]), .CLK(n4289), .Q(
        n_T_918[35]) );
  DFFX1_LVT mem_reg_wdata_reg_34_ ( .D(alu_io_out[34]), .CLK(n4288), .Q(
        n_T_918[34]) );
  DFFX1_LVT mem_reg_wdata_reg_33_ ( .D(alu_io_out[33]), .CLK(n4289), .Q(
        n_T_918[33]), .QN(n3210) );
  DFFX1_LVT mem_reg_wdata_reg_32_ ( .D(alu_io_out[32]), .CLK(n4289), .Q(
        n_T_918[32]), .QN(n3226) );
  DFFX1_LVT mem_reg_wdata_reg_31_ ( .D(alu_io_out[31]), .CLK(n4289), .Q(
        n_T_918[31]), .QN(n3105) );
  DFFX1_LVT mem_reg_wdata_reg_30_ ( .D(alu_io_out[30]), .CLK(n4290), .Q(
        n_T_918[30]), .QN(n3219) );
  DFFX1_LVT mem_reg_wdata_reg_29_ ( .D(alu_io_out[29]), .CLK(n4289), .Q(
        n_T_918[29]), .QN(n3111) );
  DFFX1_LVT mem_reg_wdata_reg_28_ ( .D(alu_io_out[28]), .CLK(n4289), .Q(
        n_T_918[28]) );
  DFFX1_LVT mem_reg_wdata_reg_27_ ( .D(alu_io_out[27]), .CLK(n4289), .Q(
        n_T_918[27]), .QN(n3209) );
  DFFX1_LVT mem_reg_wdata_reg_26_ ( .D(alu_io_out[26]), .CLK(n4289), .Q(
        n_T_918[26]), .QN(n3218) );
  DFFX1_LVT mem_reg_wdata_reg_25_ ( .D(alu_io_out[25]), .CLK(n4289), .Q(
        n_T_918[25]), .QN(n3110) );
  DFFX1_LVT mem_reg_wdata_reg_24_ ( .D(alu_io_out[24]), .CLK(n4289), .Q(
        n_T_918[24]) );
  DFFX1_LVT mem_reg_wdata_reg_23_ ( .D(alu_io_out[23]), .CLK(n4290), .Q(
        n_T_918[23]), .QN(n3213) );
  DFFX1_LVT mem_reg_wdata_reg_22_ ( .D(alu_io_out[22]), .CLK(n4289), .Q(
        n_T_918[22]), .QN(n3216) );
  DFFX1_LVT mem_reg_wdata_reg_21_ ( .D(alu_io_out[21]), .CLK(n4290), .Q(
        n_T_918[21]) );
  DFFX1_LVT mem_reg_wdata_reg_20_ ( .D(alu_io_out[20]), .CLK(n4290), .Q(
        n_T_918[20]), .QN(n3224) );
  DFFX1_LVT mem_reg_wdata_reg_19_ ( .D(alu_io_out[19]), .CLK(n4290), .Q(
        n_T_918[19]), .QN(n3212) );
  DFFX1_LVT mem_reg_wdata_reg_18_ ( .D(alu_io_out[18]), .CLK(n4290), .Q(
        n_T_918[18]), .QN(n3220) );
  DFFX1_LVT mem_reg_wdata_reg_17_ ( .D(alu_io_out[17]), .CLK(n4290), .Q(
        n_T_918[17]), .QN(n3107) );
  DFFX1_LVT mem_reg_wdata_reg_16_ ( .D(alu_io_out[16]), .CLK(n4291), .Q(
        n_T_918[16]) );
  DFFX1_LVT mem_reg_wdata_reg_15_ ( .D(alu_io_out[15]), .CLK(n4290), .Q(
        n_T_918[15]) );
  DFFX1_LVT mem_reg_wdata_reg_14_ ( .D(alu_io_out[14]), .CLK(n4290), .Q(
        n_T_918[14]), .QN(n3223) );
  DFFX1_LVT mem_reg_wdata_reg_13_ ( .D(alu_io_out[13]), .CLK(n4290), .Q(
        n_T_918[13]), .QN(n3106) );
  DFFX1_LVT mem_reg_wdata_reg_12_ ( .D(alu_io_out[12]), .CLK(n4290), .Q(
        n_T_918[12]), .QN(n3221) );
  DFFX1_LVT mem_reg_wdata_reg_11_ ( .D(alu_io_out[11]), .CLK(n4291), .Q(
        n_T_918[11]), .QN(n3211) );
  DFFX1_LVT mem_reg_wdata_reg_10_ ( .D(alu_io_out[10]), .CLK(n4290), .Q(
        n_T_918[10]), .QN(n3225) );
  DFFX1_LVT mem_reg_wdata_reg_9_ ( .D(alu_io_out[9]), .CLK(n4291), .Q(
        n_T_918[9]), .QN(n3108) );
  DFFX1_LVT mem_reg_wdata_reg_8_ ( .D(alu_io_out[8]), .CLK(n4291), .Q(
        n_T_918[8]), .QN(n3222) );
  DFFX1_LVT mem_reg_wdata_reg_7_ ( .D(alu_io_out[7]), .CLK(n4291), .Q(
        n_T_918[7]), .QN(n3214) );
  DFFX1_LVT mem_reg_wdata_reg_6_ ( .D(alu_io_out[6]), .CLK(n4291), .Q(
        n_T_918[6]), .QN(n3217) );
  DFFX1_LVT mem_reg_wdata_reg_5_ ( .D(alu_io_out[5]), .CLK(n4291), .Q(
        n_T_918[5]), .QN(n3109) );
  DFFX1_LVT mem_reg_wdata_reg_4_ ( .D(alu_io_out[4]), .CLK(n4291), .Q(
        n_T_918[4]), .QN(n3112) );
  DFFX1_LVT mem_reg_wdata_reg_3_ ( .D(alu_io_out[3]), .CLK(n4291), .Q(
        n_T_918[3]), .QN(n3208) );
  DFFX1_LVT mem_reg_wdata_reg_2_ ( .D(alu_io_out[2]), .CLK(n4292), .Q(
        n_T_918[2]) );
  DFFX1_LVT mem_reg_wdata_reg_1_ ( .D(alu_io_out[1]), .CLK(n4291), .Q(
        n_T_918[1]), .QN(n3207) );
  DFFX1_LVT mem_reg_wdata_reg_0_ ( .D(alu_io_out[0]), .CLK(n4291), .Q(
        n_T_918[0]) );
  DFFX1_LVT ex_reg_cause_reg_0_ ( .D(N303), .CLK(n4092), .QN(n80) );
  DFFX1_LVT ex_ctrl_sel_alu2_reg_1_ ( .D(N275), .CLK(n4313), .Q(
        ex_ctrl_sel_alu2[1]), .QN(n3278) );
  DFFX1_LVT ex_ctrl_sel_alu1_reg_0_ ( .D(N279), .CLK(n4313), .Q(
        ex_ctrl_sel_alu1_0_) );
  DFFSSRX1_LVT ex_ctrl_alu_fn_reg_0_ ( .D(n3583), .SETB(n1589), .RSTB(1'b1), 
        .CLK(n4312), .QN(alu_io_fn[0]) );
  DFFX1_LVT ex_ctrl_alu_fn_reg_1_ ( .D(N282), .CLK(n4313), .Q(alu_io_fn[1]) );
  DFFX1_LVT ex_ctrl_alu_fn_reg_3_ ( .D(N284), .CLK(n4313), .Q(alu_io_fn[3]) );
  DFFX1_LVT ex_ctrl_alu_dw_reg ( .D(n_GEN_9), .CLK(n4313), .Q(alu_io_dw) );
  DFFX1_LVT ex_ctrl_sel_alu2_reg_0_ ( .D(N274), .CLK(n4313), .Q(
        ex_ctrl_sel_alu2[0]) );
  DFFX1_LVT ex_reg_cause_reg_1_ ( .D(N304), .CLK(n4092), .QN(n76) );
  DFFSSRX1_LVT ex_reg_cause_reg_2_ ( .D(n9448), .SETB(
        csr_io_interrupt_cause[2]), .RSTB(n74), .CLK(n4092), .Q(n73) );
  DFFX1_LVT mem_reg_mem_size_reg_1_ ( .D(n586), .CLK(n4292), .Q(n72) );
  DFFX1_LVT mem_reg_mem_size_reg_0_ ( .D(n313), .CLK(n4291), .Q(n71) );
  DFFX1_LVT mem_ctrl_jal_reg ( .D(ex_ctrl_jal), .CLK(n4292), .Q(n3230), .QN(
        n555) );
  DFFX1_LVT mem_reg_rvc_reg ( .D(ex_reg_rvc), .CLK(n4292), .Q(mem_reg_rvc), 
        .QN(n570) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_4_ ( .D(n140), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[4]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_3_ ( .D(n141), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[3]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_2_ ( .D(n142), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[2]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_1_ ( .D(n143), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[1]) );
  DFFX1_LVT mem_reg_btb_resp_entry_reg_0_ ( .D(n144), .CLK(n4292), .QN(
        io_imem_btb_update_bits_prediction_entry[0]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_7_ ( .D(n145), .CLK(n4292), .QN(
        io_imem_bht_update_bits_prediction_history[7]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_6_ ( .D(n146), .CLK(n4292), .QN(
        io_imem_bht_update_bits_prediction_history[6]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_5_ ( .D(n147), .CLK(n4292), .QN(
        io_imem_bht_update_bits_prediction_history[5]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_4_ ( .D(n148), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[4]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_3_ ( .D(n149), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[3]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_2_ ( .D(n150), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[2]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_1_ ( .D(n151), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[1]) );
  DFFX1_LVT mem_reg_btb_resp_bht_history_reg_0_ ( .D(n152), .CLK(n4293), .QN(
        io_imem_bht_update_bits_prediction_history[0]) );
  DFFSSRX1_LVT mem_reg_load_reg ( .D(n312), .SETB(n997), .RSTB(n882), .CLK(
        n4286), .QN(mem_reg_load) );
  DFFSSRX1_LVT mem_reg_store_reg ( .D(n312), .SETB(n997), .RSTB(n996), .CLK(
        n4286), .QN(mem_reg_store) );
  DFFX1_LVT mem_ctrl_mem_reg ( .D(n312), .CLK(n4293), .Q(n572), .QN(
        mem_ctrl_mem) );
  DFFX1_LVT mem_br_taken_reg ( .D(alu_io_cmp_out), .CLK(n4293), .Q(
        io_imem_bht_update_bits_taken), .QN(n3310) );
  DFFX1_LVT mem_ctrl_wfd_reg ( .D(n315), .CLK(n4293), .Q(n69), .QN(
        mem_ctrl_wfd) );
  DFFX1_LVT mem_ctrl_div_reg ( .D(n317), .CLK(n4293), .Q(n370) );
  DFFX1_LVT mem_ctrl_wxd_reg ( .D(n314), .CLK(n4293), .QN(mem_ctrl_wxd) );
  DFFX1_LVT mem_ctrl_csr_reg_2_ ( .D(n310), .CLK(n4293), .Q(n68), .QN(
        mem_ctrl_csr[2]) );
  DFFX1_LVT mem_ctrl_csr_reg_1_ ( .D(n319), .CLK(n4294), .Q(n369), .QN(n3279)
         );
  DFFX1_LVT mem_ctrl_csr_reg_0_ ( .D(n320), .CLK(n4294), .Q(n67), .QN(
        mem_ctrl_csr[0]) );
  DFFSSRX1_LVT mem_ctrl_fence_i_reg ( .D(n9516), .SETB(ex_ctrl_jalr), .RSTB(
        n318), .CLK(n4286), .Q(n66) );
  DFFX1_LVT mem_reg_cause_reg_3_ ( .D(n75), .CLK(n4294), .QN(mem_reg_cause[3])
         );
  DFFX1_LVT mem_reg_cause_reg_2_ ( .D(n73), .CLK(n4294), .QN(mem_reg_cause[2])
         );
  DFFX1_LVT mem_reg_cause_reg_1_ ( .D(n76), .CLK(n4294), .Q(n63) );
  DFFX1_LVT mem_reg_cause_reg_0_ ( .D(n80), .CLK(n4294), .QN(mem_reg_cause[0])
         );
  DFFX1_LVT mem_reg_pc_reg_39_ ( .D(n100), .CLK(n4294), .Q(n62), .QN(
        mem_reg_pc[39]) );
  DFFX1_LVT mem_reg_pc_reg_38_ ( .D(n101), .CLK(n4294), .Q(n61), .QN(
        mem_reg_pc[38]) );
  DFFX1_LVT mem_reg_pc_reg_37_ ( .D(n102), .CLK(n4294), .Q(n60), .QN(
        mem_reg_pc[37]) );
  DFFX1_LVT mem_reg_pc_reg_36_ ( .D(n103), .CLK(n4294), .Q(n59), .QN(
        mem_reg_pc[36]) );
  DFFX1_LVT mem_reg_pc_reg_35_ ( .D(n104), .CLK(n4295), .Q(n58), .QN(
        mem_reg_pc[35]) );
  DFFX1_LVT mem_reg_pc_reg_34_ ( .D(n105), .CLK(n4295), .Q(n57), .QN(
        mem_reg_pc[34]) );
  DFFX1_LVT mem_reg_pc_reg_33_ ( .D(n106), .CLK(n4295), .Q(n56), .QN(
        mem_reg_pc[33]) );
  DFFX1_LVT mem_reg_pc_reg_32_ ( .D(n107), .CLK(n4295), .Q(n55), .QN(
        mem_reg_pc[32]) );
  DFFX1_LVT mem_reg_pc_reg_31_ ( .D(n108), .CLK(n4295), .Q(n54), .QN(
        mem_reg_pc[31]) );
  DFFX1_LVT mem_reg_pc_reg_30_ ( .D(n109), .CLK(n4295), .Q(n53), .QN(
        mem_reg_pc[30]) );
  DFFX1_LVT mem_reg_pc_reg_29_ ( .D(n110), .CLK(n4295), .Q(n52), .QN(
        mem_reg_pc[29]) );
  DFFX1_LVT mem_reg_pc_reg_28_ ( .D(n111), .CLK(n4295), .Q(n51), .QN(
        mem_reg_pc[28]) );
  DFFX1_LVT mem_reg_pc_reg_27_ ( .D(n112), .CLK(n4295), .Q(n50), .QN(
        mem_reg_pc[27]) );
  DFFX1_LVT mem_reg_pc_reg_26_ ( .D(n113), .CLK(n4295), .Q(n49), .QN(
        mem_reg_pc[26]) );
  DFFX1_LVT mem_reg_pc_reg_25_ ( .D(n114), .CLK(n4295), .Q(n48), .QN(
        mem_reg_pc[25]) );
  DFFX1_LVT mem_reg_pc_reg_24_ ( .D(n115), .CLK(n4295), .Q(n47), .QN(
        mem_reg_pc[24]) );
  DFFX1_LVT mem_reg_pc_reg_23_ ( .D(n116), .CLK(n4296), .Q(n46), .QN(
        mem_reg_pc[23]) );
  DFFX1_LVT mem_reg_pc_reg_22_ ( .D(n117), .CLK(n4296), .Q(n45), .QN(
        mem_reg_pc[22]) );
  DFFX1_LVT mem_reg_pc_reg_21_ ( .D(n118), .CLK(n4296), .Q(n44), .QN(
        mem_reg_pc[21]) );
  DFFX1_LVT mem_reg_pc_reg_20_ ( .D(n119), .CLK(n4296), .Q(n43), .QN(
        mem_reg_pc[20]) );
  DFFX1_LVT mem_reg_pc_reg_19_ ( .D(n120), .CLK(n4296), .Q(n42), .QN(
        mem_reg_pc[19]) );
  DFFX1_LVT mem_reg_pc_reg_18_ ( .D(n121), .CLK(n4296), .Q(n41), .QN(
        mem_reg_pc[18]) );
  DFFX1_LVT mem_reg_pc_reg_17_ ( .D(n122), .CLK(n4296), .Q(n40), .QN(
        mem_reg_pc[17]) );
  DFFX1_LVT mem_reg_pc_reg_16_ ( .D(n123), .CLK(n4296), .Q(n39), .QN(
        mem_reg_pc[16]) );
  DFFX1_LVT mem_reg_pc_reg_15_ ( .D(n124), .CLK(n4296), .Q(n38), .QN(
        mem_reg_pc[15]) );
  DFFX1_LVT mem_reg_pc_reg_14_ ( .D(n125), .CLK(n4296), .Q(n37), .QN(
        mem_reg_pc[14]) );
  DFFX1_LVT mem_reg_pc_reg_13_ ( .D(n126), .CLK(n4296), .Q(n36), .QN(
        mem_reg_pc[13]) );
  DFFX1_LVT mem_reg_pc_reg_12_ ( .D(n127), .CLK(n4296), .Q(n35), .QN(
        mem_reg_pc[12]) );
  DFFX1_LVT mem_reg_pc_reg_11_ ( .D(n128), .CLK(n4297), .Q(n34), .QN(
        mem_reg_pc[11]) );
  DFFX1_LVT mem_reg_pc_reg_10_ ( .D(n129), .CLK(n4297), .Q(n33), .QN(
        mem_reg_pc[10]) );
  DFFX1_LVT mem_reg_pc_reg_9_ ( .D(n130), .CLK(n4297), .Q(n32), .QN(
        mem_reg_pc[9]) );
  DFFX1_LVT mem_reg_pc_reg_8_ ( .D(n131), .CLK(n4297), .Q(n31), .QN(
        mem_reg_pc[8]) );
  DFFX1_LVT mem_reg_pc_reg_7_ ( .D(n132), .CLK(n4297), .Q(n30), .QN(
        mem_reg_pc[7]) );
  DFFX1_LVT mem_reg_pc_reg_6_ ( .D(n133), .CLK(n4297), .Q(n29), .QN(
        mem_reg_pc[6]) );
  DFFX1_LVT mem_reg_pc_reg_5_ ( .D(n134), .CLK(n4297), .Q(n28), .QN(
        mem_reg_pc[5]) );
  DFFX1_LVT mem_reg_pc_reg_4_ ( .D(n135), .CLK(n4297), .Q(n27), .QN(
        mem_reg_pc[4]) );
  DFFX1_LVT mem_reg_pc_reg_3_ ( .D(n136), .CLK(n4297), .Q(n26), .QN(
        mem_reg_pc[3]) );
  DFFX1_LVT mem_reg_pc_reg_2_ ( .D(n137), .CLK(n4297), .Q(n25), .QN(
        mem_reg_pc[2]) );
  DFFX1_LVT mem_reg_pc_reg_1_ ( .D(n138), .CLK(n4297), .Q(n24), .QN(
        mem_reg_pc[1]) );
  DFFX1_LVT mem_reg_pc_reg_0_ ( .D(n139), .CLK(n4297), .Q(n23), .QN(
        mem_reg_pc[0]) );
  DFFX1_LVT mem_reg_inst_reg_31_ ( .D(n172), .CLK(n4298), .Q(n22), .QN(
        n_T_844_10_) );
  DFFX1_LVT mem_reg_inst_reg_30_ ( .D(n171), .CLK(n4298), .Q(n21), .QN(
        n_T_849[10]) );
  DFFX1_LVT mem_reg_inst_reg_29_ ( .D(n170), .CLK(n4298), .Q(n20), .QN(
        n_T_849[9]) );
  DFFX1_LVT mem_reg_inst_reg_28_ ( .D(n169), .CLK(n4298), .Q(n19), .QN(
        n_T_849[8]) );
  DFFX1_LVT mem_reg_inst_reg_27_ ( .D(n168), .CLK(n4298), .Q(n18), .QN(
        n_T_849[7]) );
  DFFX1_LVT mem_reg_inst_reg_26_ ( .D(n167), .CLK(n4298), .Q(n17), .QN(
        n_T_849[6]) );
  DFFX1_LVT mem_reg_inst_reg_25_ ( .D(n166), .CLK(n4298), .Q(n16), .QN(
        n_T_849[5]) );
  DFFX1_LVT mem_reg_inst_reg_24_ ( .D(n165), .CLK(n4298), .Q(n15), .QN(
        n_T_911[4]) );
  DFFX1_LVT mem_reg_inst_reg_23_ ( .D(n164), .CLK(n4298), .Q(n14), .QN(
        n_T_911[3]) );
  DFFX1_LVT mem_reg_inst_reg_22_ ( .D(n163), .CLK(n4298), .Q(n13), .QN(
        n_T_911[2]) );
  DFFX1_LVT mem_reg_inst_reg_21_ ( .D(n162), .CLK(n4298), .Q(n12), .QN(
        n_T_911[1]) );
  DFFX1_LVT mem_reg_inst_reg_20_ ( .D(n161), .CLK(n4298), .Q(n11), .QN(
        n_T_911_11) );
  DFFX1_LVT mem_reg_inst_reg_19_ ( .D(n160), .CLK(n4299), .QN(n_T_904[7]) );
  DFFX1_LVT mem_reg_inst_reg_18_ ( .D(n159), .CLK(n4299), .QN(n_T_904[6]) );
  DFFX1_LVT mem_reg_inst_reg_17_ ( .D(n158), .CLK(n4299), .QN(n_T_904[5]) );
  DFFX1_LVT mem_reg_inst_reg_16_ ( .D(n157), .CLK(n4299), .QN(n_T_904[4]) );
  DFFX1_LVT mem_reg_inst_reg_15_ ( .D(n156), .CLK(n4299), .QN(n_T_904[3]) );
  DFFX1_LVT mem_reg_inst_reg_14_ ( .D(io_dmem_req_bits_signed), .CLK(n4299), 
        .QN(n_T_904[2]) );
  DFFX1_LVT mem_reg_inst_reg_13_ ( .D(n155), .CLK(n4299), .QN(n_T_904[1]) );
  DFFX1_LVT mem_reg_inst_reg_12_ ( .D(n154), .CLK(n4299), .QN(n_T_904[0]) );
  DFFX1_LVT mem_reg_inst_reg_11_ ( .D(n588), .CLK(n4299), .Q(n595), .QN(
        n_T_849[4]) );
  DFFX1_LVT mem_reg_inst_reg_10_ ( .D(n589), .CLK(n4299), .Q(n596), .QN(n2566)
         );
  DFFX1_LVT mem_reg_inst_reg_9_ ( .D(n590), .CLK(n4299), .Q(n3200), .QN(
        n_T_849[2]) );
  DFFX1_LVT mem_reg_inst_reg_8_ ( .D(n591), .CLK(n4299), .Q(n598), .QN(
        n_T_849[1]) );
  DFFX1_LVT ex_reg_rs_bypass_1_reg ( .D(do_bypass_1), .CLK(n4313), .Q(
        ex_reg_rs_bypass_1), .QN(n3243) );
  DFFX1_LVT ex_reg_load_use_reg ( .D(n9424), .CLK(n4312), .Q(ex_reg_load_use)
         );
  DFFSSRX1_LVT mem_reg_xcpt_interrupt_reg ( .D(n98), .SETB(n9418), .RSTB(1'b1), 
        .CLK(n3594), .QN(mem_reg_xcpt_interrupt) );
  DFFX1_LVT wb_ctrl_wxd_reg ( .D(mem_ctrl_wxd), .CLK(n4300), .Q(wb_ctrl_wxd)
         );
  DFFX1_LVT wb_ctrl_csr_reg_2_ ( .D(n68), .CLK(n4300), .QN(wb_ctrl_csr[2]) );
  DFFX1_LVT wb_ctrl_csr_reg_1_ ( .D(n369), .CLK(n4300), .QN(wb_ctrl_csr[1]) );
  DFFX1_LVT wb_ctrl_csr_reg_0_ ( .D(n67), .CLK(n4300), .QN(wb_ctrl_csr[0]) );
  DFFX1_LVT wb_ctrl_wfd_reg ( .D(n69), .CLK(n4300), .Q(n3229), .QN(wb_ctrl_wfd) );
  DFFX1_LVT wb_ctrl_div_reg ( .D(n370), .CLK(n4300), .QN(wb_ctrl_div) );
  DFFX1_LVT wb_ctrl_mem_reg ( .D(n572), .CLK(n4300), .QN(wb_ctrl_mem) );
  DFFX1_LVT wb_reg_wdata_reg_63_ ( .D(N661), .CLK(n4300), .Q(n_T_1165[63]) );
  DFFX1_LVT wb_reg_wdata_reg_62_ ( .D(N660), .CLK(n4300), .Q(n_T_1165[62]) );
  DFFX1_LVT wb_reg_wdata_reg_61_ ( .D(N659), .CLK(n4300), .Q(n_T_1165[61]) );
  DFFX1_LVT wb_reg_wdata_reg_60_ ( .D(N658), .CLK(n4301), .Q(n_T_1165[60]) );
  DFFX1_LVT wb_reg_wdata_reg_59_ ( .D(N657), .CLK(n4301), .Q(n_T_1165[59]) );
  DFFX1_LVT wb_reg_wdata_reg_58_ ( .D(N656), .CLK(n4301), .Q(n_T_1165[58]) );
  DFFX1_LVT wb_reg_wdata_reg_57_ ( .D(N655), .CLK(n4301), .Q(n_T_1165[57]) );
  DFFX1_LVT wb_reg_wdata_reg_56_ ( .D(N654), .CLK(n4301), .Q(n_T_1165[56]) );
  DFFX1_LVT wb_reg_wdata_reg_55_ ( .D(N653), .CLK(n4301), .Q(n_T_1165[55]) );
  DFFX1_LVT wb_reg_wdata_reg_54_ ( .D(N652), .CLK(n4301), .Q(n_T_1165[54]) );
  DFFX1_LVT wb_reg_wdata_reg_53_ ( .D(N651), .CLK(n4301), .Q(n_T_1165[53]) );
  DFFX1_LVT wb_reg_wdata_reg_52_ ( .D(N650), .CLK(n4301), .Q(n_T_1165[52]) );
  DFFX1_LVT wb_reg_wdata_reg_51_ ( .D(N649), .CLK(n4301), .Q(n_T_1165[51]) );
  DFFX1_LVT wb_reg_wdata_reg_50_ ( .D(N648), .CLK(n4301), .Q(n_T_1165[50]) );
  DFFX1_LVT wb_reg_wdata_reg_49_ ( .D(N647), .CLK(n4301), .Q(n_T_1165[49]) );
  DFFX1_LVT wb_reg_wdata_reg_48_ ( .D(N646), .CLK(n4302), .Q(n_T_1165[48]) );
  DFFX1_LVT wb_reg_wdata_reg_47_ ( .D(N645), .CLK(n4302), .Q(n_T_1165[47]) );
  DFFX1_LVT wb_reg_wdata_reg_46_ ( .D(N644), .CLK(n4302), .Q(n_T_1165[46]) );
  DFFX1_LVT wb_reg_wdata_reg_45_ ( .D(N643), .CLK(n4302), .Q(n_T_1165[45]) );
  DFFX1_LVT wb_reg_wdata_reg_44_ ( .D(N642), .CLK(n4302), .Q(n_T_1165[44]) );
  DFFX1_LVT wb_reg_wdata_reg_43_ ( .D(N641), .CLK(n4302), .Q(n_T_1165[43]) );
  DFFX1_LVT wb_reg_wdata_reg_42_ ( .D(N640), .CLK(n4302), .Q(n_T_1165[42]) );
  DFFX1_LVT wb_reg_wdata_reg_41_ ( .D(N639), .CLK(n4302), .Q(n_T_1165[41]) );
  DFFX1_LVT wb_reg_wdata_reg_40_ ( .D(N638), .CLK(n4302), .Q(n_T_1165[40]) );
  DFFX1_LVT wb_reg_wdata_reg_39_ ( .D(N637), .CLK(n4302), .Q(n_T_1165[39]) );
  DFFX1_LVT wb_reg_wdata_reg_38_ ( .D(N636), .CLK(n4302), .Q(
        io_imem_sfence_bits_addr[38]), .QN(n3228) );
  DFFX1_LVT wb_reg_wdata_reg_37_ ( .D(N635), .CLK(n4302), .Q(
        io_imem_sfence_bits_addr[37]) );
  DFFX1_LVT wb_reg_wdata_reg_36_ ( .D(N634), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[36]) );
  DFFX1_LVT wb_reg_wdata_reg_35_ ( .D(N633), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[35]) );
  DFFX1_LVT wb_reg_wdata_reg_34_ ( .D(N632), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[34]) );
  DFFX1_LVT wb_reg_wdata_reg_33_ ( .D(N631), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[33]) );
  DFFX1_LVT wb_reg_wdata_reg_32_ ( .D(N630), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[32]) );
  DFFX1_LVT wb_reg_wdata_reg_31_ ( .D(N629), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[31]) );
  DFFX1_LVT wb_reg_wdata_reg_30_ ( .D(N628), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[30]) );
  DFFX1_LVT wb_reg_wdata_reg_29_ ( .D(N627), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[29]) );
  DFFX1_LVT wb_reg_wdata_reg_28_ ( .D(N626), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[28]) );
  DFFX1_LVT wb_reg_wdata_reg_27_ ( .D(N625), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[27]) );
  DFFX1_LVT wb_reg_wdata_reg_26_ ( .D(N624), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[26]) );
  DFFX1_LVT wb_reg_wdata_reg_25_ ( .D(N623), .CLK(n4303), .Q(
        io_imem_sfence_bits_addr[25]) );
  DFFX1_LVT wb_reg_wdata_reg_24_ ( .D(N622), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[24]) );
  DFFX1_LVT wb_reg_wdata_reg_23_ ( .D(N621), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[23]) );
  DFFX1_LVT wb_reg_wdata_reg_22_ ( .D(N620), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[22]) );
  DFFX1_LVT wb_reg_wdata_reg_21_ ( .D(N619), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[21]) );
  DFFX1_LVT wb_reg_wdata_reg_20_ ( .D(N618), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[20]) );
  DFFX1_LVT wb_reg_wdata_reg_19_ ( .D(N617), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[19]) );
  DFFX1_LVT wb_reg_wdata_reg_18_ ( .D(N616), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[18]) );
  DFFX1_LVT wb_reg_wdata_reg_17_ ( .D(N615), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[17]) );
  DFFX1_LVT wb_reg_wdata_reg_16_ ( .D(N614), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[16]) );
  DFFX1_LVT wb_reg_wdata_reg_15_ ( .D(N613), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[15]) );
  DFFX1_LVT wb_reg_wdata_reg_14_ ( .D(N612), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[14]) );
  DFFX1_LVT wb_reg_wdata_reg_13_ ( .D(N611), .CLK(n4304), .Q(
        io_imem_sfence_bits_addr[13]) );
  DFFX1_LVT wb_reg_wdata_reg_12_ ( .D(N610), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[12]) );
  DFFX1_LVT wb_reg_wdata_reg_11_ ( .D(N609), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[11]) );
  DFFX1_LVT wb_reg_wdata_reg_10_ ( .D(N608), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[10]) );
  DFFX1_LVT wb_reg_wdata_reg_9_ ( .D(N607), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[9]) );
  DFFX1_LVT wb_reg_wdata_reg_8_ ( .D(N606), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[8]) );
  DFFX1_LVT wb_reg_wdata_reg_7_ ( .D(N605), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[7]) );
  DFFX1_LVT wb_reg_wdata_reg_6_ ( .D(N604), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[6]) );
  DFFX1_LVT wb_reg_wdata_reg_5_ ( .D(N603), .CLK(n4300), .Q(
        io_imem_sfence_bits_addr[5]) );
  DFFX1_LVT wb_reg_wdata_reg_4_ ( .D(N602), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[4]) );
  DFFX1_LVT wb_reg_wdata_reg_3_ ( .D(N601), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[3]) );
  DFFX1_LVT wb_reg_wdata_reg_2_ ( .D(N600), .CLK(n4305), .Q(
        io_imem_sfence_bits_addr[2]) );
  DFFX1_LVT wb_reg_wdata_reg_1_ ( .D(N599), .CLK(n4306), .Q(
        io_imem_sfence_bits_addr[1]) );
  DFFX1_LVT wb_ctrl_fence_i_reg ( .D(n66), .CLK(n4306), .QN(wb_ctrl_fence_i)
         );
  DFFX1_LVT wb_reg_sfence_reg ( .D(n326), .CLK(n4306), .QN(wb_reg_sfence) );
  DFFX1_LVT wb_reg_pc_reg_39_ ( .D(n62), .CLK(n4306), .QN(csr_io_pc[39]) );
  DFFX1_LVT wb_reg_pc_reg_38_ ( .D(n61), .CLK(n4306), .QN(csr_io_pc[38]) );
  DFFX1_LVT wb_reg_pc_reg_37_ ( .D(n60), .CLK(n4306), .QN(csr_io_pc[37]) );
  DFFX1_LVT wb_reg_pc_reg_36_ ( .D(n59), .CLK(n4306), .QN(csr_io_pc[36]) );
  DFFX1_LVT wb_reg_pc_reg_35_ ( .D(n58), .CLK(n4306), .QN(csr_io_pc[35]) );
  DFFX1_LVT wb_reg_pc_reg_34_ ( .D(n57), .CLK(n4306), .QN(csr_io_pc[34]) );
  DFFX1_LVT wb_reg_pc_reg_33_ ( .D(n56), .CLK(n4306), .QN(csr_io_pc[33]) );
  DFFX1_LVT wb_reg_pc_reg_32_ ( .D(n55), .CLK(n4306), .QN(csr_io_pc[32]) );
  DFFX1_LVT wb_reg_pc_reg_31_ ( .D(n54), .CLK(n4306), .QN(csr_io_pc[31]) );
  DFFX1_LVT wb_reg_pc_reg_30_ ( .D(n53), .CLK(n4307), .QN(csr_io_pc[30]) );
  DFFX1_LVT wb_reg_pc_reg_29_ ( .D(n52), .CLK(n4307), .QN(csr_io_pc[29]) );
  DFFX1_LVT wb_reg_pc_reg_28_ ( .D(n51), .CLK(n4307), .QN(csr_io_pc[28]) );
  DFFX1_LVT wb_reg_pc_reg_27_ ( .D(n50), .CLK(n4307), .QN(csr_io_pc[27]) );
  DFFX1_LVT wb_reg_pc_reg_26_ ( .D(n49), .CLK(n4307), .QN(csr_io_pc[26]) );
  DFFX1_LVT wb_reg_pc_reg_25_ ( .D(n48), .CLK(n4307), .QN(csr_io_pc[25]) );
  DFFX1_LVT wb_reg_pc_reg_24_ ( .D(n47), .CLK(n4307), .QN(csr_io_pc[24]) );
  DFFX1_LVT wb_reg_pc_reg_23_ ( .D(n46), .CLK(n4307), .QN(csr_io_pc[23]) );
  DFFX1_LVT wb_reg_pc_reg_22_ ( .D(n45), .CLK(n4307), .QN(csr_io_pc[22]) );
  DFFX1_LVT wb_reg_pc_reg_21_ ( .D(n44), .CLK(n4307), .QN(csr_io_pc[21]) );
  DFFX1_LVT wb_reg_pc_reg_20_ ( .D(n43), .CLK(n4307), .QN(csr_io_pc[20]) );
  DFFX1_LVT wb_reg_pc_reg_19_ ( .D(n42), .CLK(n4307), .QN(csr_io_pc[19]) );
  DFFX1_LVT wb_reg_pc_reg_18_ ( .D(n41), .CLK(n4308), .QN(csr_io_pc[18]) );
  DFFX1_LVT wb_reg_pc_reg_17_ ( .D(n40), .CLK(n4308), .QN(csr_io_pc[17]) );
  DFFX1_LVT wb_reg_pc_reg_16_ ( .D(n39), .CLK(n4308), .QN(csr_io_pc[16]) );
  DFFX1_LVT wb_reg_pc_reg_15_ ( .D(n38), .CLK(n4308), .QN(csr_io_pc[15]) );
  DFFX1_LVT wb_reg_pc_reg_14_ ( .D(n37), .CLK(n4308), .QN(csr_io_pc[14]) );
  DFFX1_LVT wb_reg_pc_reg_13_ ( .D(n36), .CLK(n4308), .QN(csr_io_pc[13]) );
  DFFX1_LVT wb_reg_pc_reg_12_ ( .D(n35), .CLK(n4308), .QN(csr_io_pc[12]) );
  DFFX1_LVT wb_reg_pc_reg_11_ ( .D(n34), .CLK(n4308), .QN(csr_io_pc[11]) );
  DFFX1_LVT wb_reg_pc_reg_10_ ( .D(n33), .CLK(n4308), .QN(csr_io_pc[10]) );
  DFFX1_LVT wb_reg_pc_reg_9_ ( .D(n32), .CLK(n4308), .QN(csr_io_pc[9]) );
  DFFX1_LVT wb_reg_pc_reg_8_ ( .D(n31), .CLK(n4308), .QN(csr_io_pc[8]) );
  DFFX1_LVT wb_reg_pc_reg_7_ ( .D(n30), .CLK(n4308), .QN(csr_io_pc[7]) );
  DFFX1_LVT wb_reg_pc_reg_6_ ( .D(n29), .CLK(n4309), .QN(csr_io_pc[6]) );
  DFFX1_LVT wb_reg_pc_reg_5_ ( .D(n28), .CLK(n4309), .QN(csr_io_pc[5]) );
  DFFX1_LVT wb_reg_pc_reg_4_ ( .D(n27), .CLK(n4309), .QN(csr_io_pc[4]) );
  DFFX1_LVT wb_reg_pc_reg_3_ ( .D(n26), .CLK(n4309), .QN(csr_io_pc[3]) );
  DFFX1_LVT wb_reg_pc_reg_2_ ( .D(n25), .CLK(n4309), .QN(csr_io_pc[2]) );
  DFFX1_LVT wb_reg_pc_reg_1_ ( .D(n24), .CLK(n4309), .QN(csr_io_pc[1]) );
  DFFX1_LVT wb_reg_pc_reg_0_ ( .D(n23), .CLK(n4309), .QN(csr_io_pc[0]) );
  DFFX1_LVT wb_reg_mem_size_reg_1_ ( .D(n72), .CLK(n4309), .QN(
        io_imem_sfence_bits_rs2) );
  DFFX1_LVT wb_reg_mem_size_reg_0_ ( .D(n71), .CLK(n4309), .QN(
        io_imem_sfence_bits_rs1) );
  DFFX1_LVT wb_reg_inst_reg_31_ ( .D(n22), .CLK(n4309), .QN(csr_io_rw_addr[11]) );
  DFFX1_LVT wb_reg_inst_reg_30_ ( .D(n21), .CLK(n4309), .QN(csr_io_rw_addr[10]) );
  DFFX1_LVT wb_reg_inst_reg_29_ ( .D(n20), .CLK(n4309), .QN(csr_io_rw_addr[9])
         );
  DFFX1_LVT wb_reg_inst_reg_28_ ( .D(n19), .CLK(n4310), .QN(csr_io_rw_addr[8])
         );
  DFFX1_LVT wb_reg_inst_reg_27_ ( .D(n18), .CLK(n4310), .QN(csr_io_rw_addr[7])
         );
  DFFX1_LVT wb_reg_inst_reg_26_ ( .D(n17), .CLK(n4310), .QN(csr_io_rw_addr[6])
         );
  DFFX1_LVT wb_reg_inst_reg_25_ ( .D(n16), .CLK(n4310), .QN(csr_io_rw_addr[5])
         );
  DFFX1_LVT wb_reg_inst_reg_24_ ( .D(n15), .CLK(n4310), .QN(csr_io_rw_addr[4])
         );
  DFFX1_LVT wb_reg_inst_reg_23_ ( .D(n14), .CLK(n4310), .QN(csr_io_rw_addr[3])
         );
  DFFX1_LVT wb_reg_inst_reg_22_ ( .D(n13), .CLK(n4310), .QN(csr_io_rw_addr[2])
         );
  DFFX1_LVT wb_reg_inst_reg_21_ ( .D(n12), .CLK(n4310), .QN(csr_io_rw_addr[1])
         );
  DFFX1_LVT wb_reg_inst_reg_20_ ( .D(n11), .CLK(n4310), .QN(csr_io_rw_addr[0])
         );
  DFFX1_LVT wb_reg_inst_reg_11_ ( .D(n_T_849[4]), .CLK(n4310), .Q(wb_waddr[4]), 
        .QN(n3198) );
  DFFX1_LVT wb_reg_inst_reg_10_ ( .D(n2566), .CLK(n4310), .Q(wb_waddr[3]), 
        .QN(n3199) );
  DFFX1_LVT wb_reg_inst_reg_9_ ( .D(n_T_849[2]), .CLK(n4310), .Q(n3043), .QN(
        n3102) );
  DFFX1_LVT wb_reg_inst_reg_7_ ( .D(n_T_849[11]), .CLK(n4311), .Q(n3041), .QN(
        n3201) );
  DFFX1_LVT wb_reg_cause_reg_0_ ( .D(N533), .CLK(n4311), .Q(wb_reg_cause[0])
         );
  DFFX1_LVT wb_reg_cause_reg_2_ ( .D(N535), .CLK(n4311), .Q(wb_reg_cause[2])
         );
  DFFX1_LVT wb_reg_cause_reg_3_ ( .D(N536), .CLK(n4305), .QN(n3565) );
  DFFX1_LVT wb_reg_xcpt_reg ( .D(N529), .CLK(n3594), .Q(n3262), .QN(n576) );
  DFFX1_LVT ex_reg_rs_lsb_1_reg_0_ ( .D(N678), .CLK(n4312), .Q(n5481), .QN(
        n594) );
  DFFX1_LVT ex_reg_rs_lsb_1_reg_1_ ( .D(N679), .CLK(n4313), .Q(n_T_635[1]) );
  DFFX1_LVT mem_reg_rs2_reg_0_ ( .D(n_T_702[0]), .CLK(n4091), .Q(
        mem_reg_rs2[0]) );
  DFFX1_LVT mem_reg_rs2_reg_1_ ( .D(n_T_702[1]), .CLK(n4091), .Q(
        mem_reg_rs2[1]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_8_ ( .D(id_rs_1[10]), .CLK(n4079), .Q(
        n_T_635[10]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_9_ ( .D(id_rs_1[11]), .CLK(n4078), .Q(
        n_T_635[11]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_10_ ( .D(id_rs_1[12]), .CLK(n4078), .Q(
        n_T_635[12]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_11_ ( .D(id_rs_1[13]), .CLK(n4078), .Q(
        n_T_635[13]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_12_ ( .D(id_rs_1[14]), .CLK(n4078), .Q(
        n_T_635[14]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_13_ ( .D(id_rs_1[15]), .CLK(n4078), .Q(
        n_T_635[15]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_14_ ( .D(id_rs_1[16]), .CLK(n4078), .Q(
        n_T_635[16]) );
  DFFX1_LVT mem_reg_rs2_reg_16_ ( .D(N477), .CLK(n4091), .Q(mem_reg_rs2[16])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_15_ ( .D(id_rs_1[17]), .CLK(n4078), .Q(
        n_T_635[17]) );
  DFFX1_LVT mem_reg_rs2_reg_17_ ( .D(N478), .CLK(n4091), .Q(mem_reg_rs2[17])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_16_ ( .D(id_rs_1[18]), .CLK(n4078), .Q(
        n_T_635[18]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_17_ ( .D(id_rs_1[19]), .CLK(n4078), .Q(
        n_T_635[19]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_18_ ( .D(id_rs_1[20]), .CLK(n4078), .Q(
        n_T_635[20]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_19_ ( .D(id_rs_1[21]), .CLK(n4078), .Q(
        n_T_635[21]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_20_ ( .D(id_rs_1[22]), .CLK(n4078), .Q(
        n_T_635[22]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_21_ ( .D(id_rs_1[23]), .CLK(n4077), .Q(
        n_T_635[23]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_22_ ( .D(id_rs_1[24]), .CLK(n4077), .Q(
        n_T_635[24]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_23_ ( .D(id_rs_1[25]), .CLK(n4077), .Q(
        n_T_635[25]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_24_ ( .D(id_rs_1[26]), .CLK(n4077), .Q(
        n_T_635[26]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_25_ ( .D(id_rs_1[27]), .CLK(n4077), .Q(
        n_T_635[27]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_26_ ( .D(id_rs_1[28]), .CLK(n4077), .Q(
        n_T_635[28]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_27_ ( .D(id_rs_1[29]), .CLK(n4077), .Q(
        n_T_635[29]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_0_ ( .D(id_rs_1[2]), .CLK(n4077), .Q(
        n_T_635[2]) );
  DFFX1_LVT mem_reg_rs2_reg_26_ ( .D(N487), .CLK(n4090), .Q(mem_reg_rs2[26])
         );
  DFFX1_LVT mem_reg_rs2_reg_18_ ( .D(N479), .CLK(n4090), .Q(mem_reg_rs2[18])
         );
  DFFX1_LVT mem_reg_rs2_reg_10_ ( .D(N471), .CLK(n4090), .Q(mem_reg_rs2[10])
         );
  DFFX1_LVT mem_reg_rs2_reg_2_ ( .D(n_T_702[2]), .CLK(n4090), .Q(
        mem_reg_rs2[2]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_28_ ( .D(id_rs_1[30]), .CLK(n4077), .Q(
        n_T_635[30]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_29_ ( .D(id_rs_1[31]), .CLK(n4077), .Q(
        n_T_635[31]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_30_ ( .D(id_rs_1[32]), .CLK(n4077), .Q(
        n_T_635[32]) );
  DFFX1_LVT mem_reg_rs2_reg_32_ ( .D(N493), .CLK(n4090), .Q(mem_reg_rs2[32])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_31_ ( .D(id_rs_1[33]), .CLK(n4077), .Q(
        n_T_635[33]) );
  DFFX1_LVT mem_reg_rs2_reg_33_ ( .D(N494), .CLK(n4090), .Q(mem_reg_rs2[33])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_32_ ( .D(id_rs_1[34]), .CLK(n4076), .Q(
        n_T_635[34]) );
  DFFX1_LVT mem_reg_rs2_reg_34_ ( .D(N495), .CLK(n4090), .Q(mem_reg_rs2[34])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_33_ ( .D(id_rs_1[35]), .CLK(n4076), .Q(
        n_T_635[35]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_34_ ( .D(id_rs_1[36]), .CLK(n4076), .Q(
        n_T_635[36]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_35_ ( .D(id_rs_1[37]), .CLK(n4076), .Q(
        n_T_635[37]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_36_ ( .D(id_rs_1[38]), .CLK(n4076), .Q(
        n_T_635[38]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_37_ ( .D(id_rs_1[39]), .CLK(n4076), .Q(
        n_T_635[39]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_1_ ( .D(id_rs_1[3]), .CLK(n4076), .Q(
        n_T_635[3]) );
  DFFX1_LVT mem_reg_rs2_reg_35_ ( .D(N496), .CLK(n4090), .Q(mem_reg_rs2[35])
         );
  DFFX1_LVT mem_reg_rs2_reg_27_ ( .D(N488), .CLK(n4090), .Q(mem_reg_rs2[27])
         );
  DFFX1_LVT mem_reg_rs2_reg_19_ ( .D(N480), .CLK(n4090), .Q(mem_reg_rs2[19])
         );
  DFFX1_LVT mem_reg_rs2_reg_11_ ( .D(N472), .CLK(n4090), .Q(mem_reg_rs2[11])
         );
  DFFX1_LVT mem_reg_rs2_reg_3_ ( .D(n_T_702[3]), .CLK(n4090), .Q(
        mem_reg_rs2[3]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_38_ ( .D(id_rs_1[40]), .CLK(n4076), .Q(
        n_T_635[40]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_39_ ( .D(id_rs_1[41]), .CLK(n4076), .Q(
        n_T_635[41]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_40_ ( .D(id_rs_1[42]), .CLK(n4076), .Q(
        n_T_635[42]) );
  DFFX1_LVT mem_reg_rs2_reg_42_ ( .D(N503), .CLK(n4089), .Q(mem_reg_rs2[42])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_41_ ( .D(id_rs_1[43]), .CLK(n4076), .Q(
        n_T_635[43]) );
  DFFX1_LVT mem_reg_rs2_reg_43_ ( .D(N504), .CLK(n4089), .Q(mem_reg_rs2[43])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_42_ ( .D(id_rs_1[44]), .CLK(n4076), .Q(
        n_T_635[44]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_43_ ( .D(id_rs_1[45]), .CLK(n4075), .Q(
        n_T_635[45]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_44_ ( .D(id_rs_1[46]), .CLK(n4075), .Q(
        n_T_635[46]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_45_ ( .D(id_rs_1[47]), .CLK(n4075), .Q(
        n_T_635[47]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_46_ ( .D(id_rs_1[48]), .CLK(n4075), .Q(
        n_T_635[48]) );
  DFFX1_LVT mem_reg_rs2_reg_48_ ( .D(N509), .CLK(n4089), .Q(mem_reg_rs2[48])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_47_ ( .D(id_rs_1[49]), .CLK(n4075), .Q(
        n_T_635[49]) );
  DFFX1_LVT mem_reg_rs2_reg_49_ ( .D(N510), .CLK(n4089), .Q(mem_reg_rs2[49])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_2_ ( .D(id_rs_1[4]), .CLK(n4075), .Q(
        n_T_635[4]) );
  DFFX1_LVT mem_reg_rs2_reg_36_ ( .D(N497), .CLK(n4089), .Q(mem_reg_rs2[36])
         );
  DFFX1_LVT mem_reg_rs2_reg_28_ ( .D(N489), .CLK(n4089), .Q(mem_reg_rs2[28])
         );
  DFFX1_LVT mem_reg_rs2_reg_20_ ( .D(N481), .CLK(n4089), .Q(mem_reg_rs2[20])
         );
  DFFX1_LVT mem_reg_rs2_reg_44_ ( .D(N505), .CLK(n4089), .Q(mem_reg_rs2[44])
         );
  DFFX1_LVT mem_reg_rs2_reg_12_ ( .D(N473), .CLK(n4089), .Q(mem_reg_rs2[12])
         );
  DFFX1_LVT mem_reg_rs2_reg_4_ ( .D(n_T_702[4]), .CLK(n4089), .Q(
        mem_reg_rs2[4]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_48_ ( .D(id_rs_1[50]), .CLK(n4075), .Q(
        n_T_635[50]) );
  DFFX1_LVT mem_reg_rs2_reg_50_ ( .D(N511), .CLK(n4089), .Q(mem_reg_rs2[50])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_49_ ( .D(id_rs_1[51]), .CLK(n4075), .Q(
        n_T_635[51]) );
  DFFX1_LVT mem_reg_rs2_reg_51_ ( .D(N512), .CLK(n4089), .Q(mem_reg_rs2[51])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_50_ ( .D(id_rs_1[52]), .CLK(n4075), .Q(
        n_T_635[52]) );
  DFFX1_LVT mem_reg_rs2_reg_52_ ( .D(N513), .CLK(n4088), .Q(mem_reg_rs2[52])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_51_ ( .D(id_rs_1[53]), .CLK(n4075), .Q(
        n_T_635[53]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_52_ ( .D(id_rs_1[54]), .CLK(n4075), .Q(
        n_T_635[54]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_53_ ( .D(id_rs_1[55]), .CLK(n4075), .Q(
        n_T_635[55]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_54_ ( .D(id_rs_1[56]), .CLK(n4074), .Q(
        n_T_635[56]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_55_ ( .D(id_rs_1[57]), .CLK(n4074), .Q(
        n_T_635[57]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_56_ ( .D(id_rs_1[58]), .CLK(n4074), .Q(
        n_T_635[58]) );
  DFFX1_LVT mem_reg_rs2_reg_58_ ( .D(N519), .CLK(n4088), .Q(mem_reg_rs2[58])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_57_ ( .D(id_rs_1[59]), .CLK(n4074), .Q(
        n_T_635[59]) );
  DFFX1_LVT mem_reg_rs2_reg_59_ ( .D(N520), .CLK(n4088), .Q(mem_reg_rs2[59])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_3_ ( .D(id_rs_1[5]), .CLK(n4074), .Q(
        n_T_635[5]) );
  DFFX1_LVT mem_reg_rs2_reg_37_ ( .D(N498), .CLK(n4088), .Q(mem_reg_rs2[37])
         );
  DFFX1_LVT mem_reg_rs2_reg_29_ ( .D(N490), .CLK(n4088), .Q(mem_reg_rs2[29])
         );
  DFFX1_LVT mem_reg_rs2_reg_53_ ( .D(N514), .CLK(n4088), .Q(mem_reg_rs2[53])
         );
  DFFX1_LVT mem_reg_rs2_reg_21_ ( .D(N482), .CLK(n4088), .Q(mem_reg_rs2[21])
         );
  DFFX1_LVT mem_reg_rs2_reg_45_ ( .D(N506), .CLK(n4088), .Q(mem_reg_rs2[45])
         );
  DFFX1_LVT mem_reg_rs2_reg_13_ ( .D(N474), .CLK(n4088), .Q(mem_reg_rs2[13])
         );
  DFFX1_LVT mem_reg_rs2_reg_5_ ( .D(n_T_702[5]), .CLK(n4088), .Q(
        mem_reg_rs2[5]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_58_ ( .D(id_rs_1[60]), .CLK(n4074), .Q(
        n_T_635[60]) );
  DFFX1_LVT mem_reg_rs2_reg_60_ ( .D(N521), .CLK(n4088), .Q(mem_reg_rs2[60])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_59_ ( .D(id_rs_1[61]), .CLK(n4074), .Q(
        n_T_635[61]) );
  DFFX1_LVT mem_reg_rs2_reg_61_ ( .D(N522), .CLK(n4088), .Q(mem_reg_rs2[61])
         );
  DFFX1_LVT ex_reg_rs_msb_1_reg_60_ ( .D(id_rs_1[62]), .CLK(n4074), .Q(
        n_T_635[62]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_4_ ( .D(id_rs_1[6]), .CLK(n4074), .Q(
        n_T_635[6]) );
  DFFX1_LVT mem_reg_rs2_reg_38_ ( .D(N499), .CLK(n4087), .Q(mem_reg_rs2[38])
         );
  DFFX1_LVT mem_reg_rs2_reg_62_ ( .D(N523), .CLK(n4087), .Q(mem_reg_rs2[62])
         );
  DFFX1_LVT mem_reg_rs2_reg_30_ ( .D(N491), .CLK(n4087), .Q(mem_reg_rs2[30])
         );
  DFFX1_LVT mem_reg_rs2_reg_54_ ( .D(N515), .CLK(n4087), .Q(mem_reg_rs2[54])
         );
  DFFX1_LVT mem_reg_rs2_reg_22_ ( .D(N483), .CLK(n4087), .Q(mem_reg_rs2[22])
         );
  DFFX1_LVT mem_reg_rs2_reg_46_ ( .D(N507), .CLK(n4087), .Q(mem_reg_rs2[46])
         );
  DFFX1_LVT mem_reg_rs2_reg_14_ ( .D(N475), .CLK(n4087), .Q(mem_reg_rs2[14])
         );
  DFFX1_LVT mem_reg_rs2_reg_6_ ( .D(n_T_702[6]), .CLK(n4087), .Q(
        mem_reg_rs2[6]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_5_ ( .D(id_rs_1[7]), .CLK(n4074), .Q(
        n_T_635[7]) );
  DFFX1_LVT mem_reg_rs2_reg_39_ ( .D(N500), .CLK(n4087), .Q(mem_reg_rs2[39])
         );
  DFFX1_LVT mem_reg_rs2_reg_63_ ( .D(N524), .CLK(n4087), .Q(mem_reg_rs2[63])
         );
  DFFX1_LVT mem_reg_rs2_reg_31_ ( .D(N492), .CLK(n4087), .Q(mem_reg_rs2[31])
         );
  DFFX1_LVT mem_reg_rs2_reg_55_ ( .D(N516), .CLK(n4087), .Q(mem_reg_rs2[55])
         );
  DFFX1_LVT mem_reg_rs2_reg_23_ ( .D(N484), .CLK(n4086), .Q(mem_reg_rs2[23])
         );
  DFFX1_LVT mem_reg_rs2_reg_47_ ( .D(N508), .CLK(n4086), .Q(mem_reg_rs2[47])
         );
  DFFX1_LVT mem_reg_rs2_reg_15_ ( .D(N476), .CLK(n4086), .Q(mem_reg_rs2[15])
         );
  DFFX1_LVT mem_reg_rs2_reg_7_ ( .D(n_T_702[7]), .CLK(n4086), .Q(
        mem_reg_rs2[7]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_6_ ( .D(id_rs_1[8]), .CLK(n4074), .Q(
        n_T_635[8]) );
  DFFX1_LVT mem_reg_rs2_reg_40_ ( .D(N501), .CLK(n4086), .Q(mem_reg_rs2[40])
         );
  DFFX1_LVT mem_reg_rs2_reg_56_ ( .D(N517), .CLK(n4086), .Q(mem_reg_rs2[56])
         );
  DFFX1_LVT mem_reg_rs2_reg_24_ ( .D(N485), .CLK(n4086), .Q(mem_reg_rs2[24])
         );
  DFFX1_LVT mem_reg_rs2_reg_8_ ( .D(N469), .CLK(n4086), .Q(mem_reg_rs2[8]) );
  DFFX1_LVT ex_reg_rs_msb_1_reg_7_ ( .D(id_rs_1[9]), .CLK(n4074), .Q(
        n_T_635[9]) );
  DFFX1_LVT mem_reg_rs2_reg_41_ ( .D(N502), .CLK(n4086), .Q(mem_reg_rs2[41])
         );
  DFFX1_LVT mem_reg_rs2_reg_57_ ( .D(N518), .CLK(n4086), .Q(mem_reg_rs2[57])
         );
  DFFX1_LVT mem_reg_rs2_reg_25_ ( .D(N486), .CLK(n4086), .Q(mem_reg_rs2[25])
         );
  DFFX1_LVT mem_reg_rs2_reg_9_ ( .D(N470), .CLK(n4086), .Q(mem_reg_rs2[9]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_60_ ( .D(N742), .CLK(n4085), .Q(n_T_628[62])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_58_ ( .D(N740), .CLK(n4084), .Q(n_T_628[60])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_57_ ( .D(N739), .CLK(n4084), .Q(n_T_628[59])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_55_ ( .D(N737), .CLK(n4084), .Q(n_T_628[57])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_54_ ( .D(N736), .CLK(n4084), .Q(n_T_628[56])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_52_ ( .D(N734), .CLK(n4084), .Q(n_T_628[54])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_51_ ( .D(N733), .CLK(n4084), .Q(n_T_628[53])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_49_ ( .D(N731), .CLK(n4084), .Q(n_T_628[51])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_48_ ( .D(N730), .CLK(n4084), .Q(n_T_628[50])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_47_ ( .D(N729), .CLK(n4083), .Q(n_T_628[49])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_46_ ( .D(N728), .CLK(n4083), .Q(n_T_628[48])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_45_ ( .D(N727), .CLK(n4083), .Q(n_T_628[47])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_44_ ( .D(N726), .CLK(n4083), .Q(n_T_628[46])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_43_ ( .D(N725), .CLK(n4083), .Q(n_T_628[45])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_42_ ( .D(N724), .CLK(n4083), .Q(n_T_628[44])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_41_ ( .D(N723), .CLK(n4083), .Q(n_T_628[43])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_40_ ( .D(N722), .CLK(n4083), .Q(n_T_628[42])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_37_ ( .D(N719), .CLK(n4083), .Q(n_T_628[39])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_36_ ( .D(N718), .CLK(n4083), .Q(n_T_628[38])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_35_ ( .D(N717), .CLK(n4082), .Q(n_T_628[37])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_34_ ( .D(N716), .CLK(n4082), .Q(n_T_628[36])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_31_ ( .D(N713), .CLK(n4082), .Q(n_T_628[33])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_30_ ( .D(N712), .CLK(n4082), .Q(n_T_628[32])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_29_ ( .D(N711), .CLK(n4082), .Q(n_T_628[31])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_28_ ( .D(N710), .CLK(n4082), .Q(n_T_628[30])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_27_ ( .D(N709), .CLK(n4082), .Q(n_T_628[29])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_26_ ( .D(N708), .CLK(n4082), .Q(n_T_628[28])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_25_ ( .D(N707), .CLK(n4082), .Q(n_T_628[27])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_24_ ( .D(N706), .CLK(n4082), .Q(n_T_628[26])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_23_ ( .D(N705), .CLK(n4081), .Q(n_T_628[25])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_22_ ( .D(N704), .CLK(n4081), .Q(n_T_628[24])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_21_ ( .D(N703), .CLK(n4081), .Q(n_T_628[23])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_20_ ( .D(N702), .CLK(n4081), .Q(n_T_628[22])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_19_ ( .D(N701), .CLK(n4081), .Q(n_T_628[21])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_18_ ( .D(N700), .CLK(n4081), .Q(n_T_628[20])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_17_ ( .D(N699), .CLK(n4081), .Q(n_T_628[19])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_16_ ( .D(N698), .CLK(n4081), .Q(n_T_628[18])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_15_ ( .D(N697), .CLK(n4081), .Q(n_T_628[17])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_14_ ( .D(N696), .CLK(n4081), .Q(n_T_628[16])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_13_ ( .D(N695), .CLK(n4081), .Q(n_T_628[15])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_12_ ( .D(N694), .CLK(n4081), .Q(n_T_628[14])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_11_ ( .D(N693), .CLK(n4080), .Q(n_T_628[13])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_10_ ( .D(N692), .CLK(n4080), .Q(n_T_628[12])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_9_ ( .D(N691), .CLK(n4080), .Q(n_T_628[11]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_8_ ( .D(N690), .CLK(n4080), .Q(n_T_628[10]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_7_ ( .D(N689), .CLK(n4080), .Q(n_T_628[9]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_6_ ( .D(N688), .CLK(n4080), .Q(n_T_628[8]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_5_ ( .D(N687), .CLK(n4080), .Q(n_T_628[7]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_4_ ( .D(N686), .CLK(n4080), .Q(n_T_628[6]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_3_ ( .D(N685), .CLK(n4080), .Q(n_T_628[5]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_2_ ( .D(N684), .CLK(n4080), .Q(n_T_628[4]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_1_ ( .D(N683), .CLK(n4080), .Q(n_T_628[3]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_0_ ( .D(N682), .CLK(n4080), .Q(n_T_628[2]) );
  DFFX1_LVT ex_reg_rs_lsb_0_reg_1_ ( .D(N673), .CLK(n4312), .Q(n_T_628[1]), 
        .QN(n3255) );
  DFFX1_LVT ex_reg_rs_lsb_0_reg_0_ ( .D(N672), .CLK(n4313), .Q(n7019), .QN(
        n569) );
  DFFX1_LVT u_T_427_reg_0__63_ ( .D(n4494), .CLK(n4284), .Q(n_T_427[1942]), 
        .QN(n3529) );
  DFFX1_LVT u_T_427_reg_0__62_ ( .D(n4491), .CLK(n4284), .Q(n_T_427[1941]), 
        .QN(n3484) );
  DFFX1_LVT u_T_427_reg_0__61_ ( .D(n4488), .CLK(n4284), .Q(n_T_427[1940]), 
        .QN(n3483) );
  DFFX1_LVT u_T_427_reg_0__60_ ( .D(n4485), .CLK(n4284), .Q(n_T_427[1939]) );
  DFFX1_LVT u_T_427_reg_0__58_ ( .D(n4479), .CLK(n4283), .Q(n_T_427[1937]), 
        .QN(n3492) );
  DFFX1_LVT u_T_427_reg_0__56_ ( .D(n4473), .CLK(n4283), .Q(n_T_427[1935]), 
        .QN(n3564) );
  DFFX1_LVT u_T_427_reg_0__54_ ( .D(n4467), .CLK(n4283), .Q(n_T_427[1933]), 
        .QN(n3562) );
  DFFX1_LVT u_T_427_reg_0__52_ ( .D(n4461), .CLK(n4283), .Q(n_T_427[1931]), 
        .QN(n3560) );
  DFFX1_LVT u_T_427_reg_0__51_ ( .D(n4458), .CLK(n4283), .Q(n_T_427[1930]), 
        .QN(n3559) );
  DFFX1_LVT u_T_427_reg_0__49_ ( .D(n4452), .CLK(n4283), .Q(n_T_427[1929]), 
        .QN(n3558) );
  DFFX1_LVT u_T_427_reg_0__46_ ( .D(n4443), .CLK(n4282), .Q(n_T_427[1926]) );
  DFFX1_LVT u_T_427_reg_0__45_ ( .D(n4440), .CLK(n4282), .Q(n_T_427[1925]), 
        .QN(n3555) );
  DFFX1_LVT u_T_427_reg_0__44_ ( .D(n4437), .CLK(n4282), .Q(n_T_427[1924]), 
        .QN(n2496) );
  DFFX1_LVT u_T_427_reg_0__43_ ( .D(n4434), .CLK(n4282), .Q(n_T_427[1923]), 
        .QN(n3554) );
  DFFX1_LVT u_T_427_reg_0__42_ ( .D(n4431), .CLK(n4282), .Q(n_T_427[1922]), 
        .QN(n3553) );
  DFFX1_LVT u_T_427_reg_0__41_ ( .D(n4428), .CLK(n4282), .Q(n_T_427[1921]), 
        .QN(n3552) );
  DFFX1_LVT u_T_427_reg_0__39_ ( .D(n4422), .CLK(n4282), .Q(n_T_427[1919]) );
  DFFX1_LVT u_T_427_reg_0__38_ ( .D(n4420), .CLK(n4282), .Q(n_T_427[1918]) );
  DFFX1_LVT u_T_427_reg_0__36_ ( .D(n4414), .CLK(n4282), .Q(n_T_427[1916]), 
        .QN(n3549) );
  DFFX1_LVT u_T_427_reg_0__35_ ( .D(n4412), .CLK(n4281), .Q(n_T_427[1915]) );
  DFFX1_LVT u_T_427_reg_0__34_ ( .D(n4409), .CLK(n4281), .Q(n_T_427[1914]) );
  DFFX1_LVT u_T_427_reg_0__33_ ( .D(n4407), .CLK(n4281), .Q(n_T_427[1913]) );
  DFFX1_LVT u_T_427_reg_0__31_ ( .D(n4402), .CLK(n4281), .Q(n_T_427[1912]) );
  DFFX1_LVT u_T_427_reg_0__30_ ( .D(n4399), .CLK(n4281), .Q(n_T_427[1911]), 
        .QN(n3547) );
  DFFX1_LVT u_T_427_reg_0__29_ ( .D(n4396), .CLK(n4281), .Q(n_T_427[1910]) );
  DFFX1_LVT u_T_427_reg_0__28_ ( .D(n4394), .CLK(n4281), .Q(n_T_427[1909]) );
  DFFX1_LVT u_T_427_reg_0__27_ ( .D(n4391), .CLK(n4281), .Q(n_T_427[1908]) );
  DFFX1_LVT u_T_427_reg_0__26_ ( .D(n4389), .CLK(n4281), .Q(n_T_427[1907]) );
  DFFX1_LVT u_T_427_reg_0__25_ ( .D(n4387), .CLK(n4281), .Q(n_T_427[1906]) );
  DFFX1_LVT u_T_427_reg_0__24_ ( .D(n4384), .CLK(n4281), .Q(n_T_427[1905]), 
        .QN(n3545) );
  DFFX1_LVT u_T_427_reg_0__23_ ( .D(n4381), .CLK(n4280), .Q(n_T_427[1904]) );
  DFFX1_LVT u_T_427_reg_0__22_ ( .D(n4379), .CLK(n4280), .Q(n_T_427[1903]), 
        .QN(n2684) );
  DFFX1_LVT u_T_427_reg_0__21_ ( .D(n4377), .CLK(n4280), .Q(n_T_427[1902]) );
  DFFX1_LVT u_T_427_reg_0__20_ ( .D(n4374), .CLK(n4280), .Q(n_T_427[1901]), 
        .QN(n3544) );
  DFFX1_LVT u_T_427_reg_0__19_ ( .D(n4371), .CLK(n4280), .Q(n_T_427[1900]), 
        .QN(n3543) );
  DFFX1_LVT u_T_427_reg_0__18_ ( .D(n4368), .CLK(n4280), .Q(n_T_427[1899]), 
        .QN(n3542) );
  DFFX1_LVT u_T_427_reg_0__14_ ( .D(n4357), .CLK(n4280), .Q(n_T_427[1895]) );
  DFFX1_LVT u_T_427_reg_0__11_ ( .D(n4351), .CLK(n4279), .Q(n_T_427[1892]) );
  DFFX1_LVT u_T_427_reg_0__5_ ( .D(n4331), .CLK(n4279), .Q(n_T_427[1886]) );
  DFFX1_LVT u_T_427_reg_0__4_ ( .D(n4328), .CLK(n4279), .Q(n_T_427[1885]) );
  DFFX1_LVT u_T_427_reg_0__2_ ( .D(n4322), .CLK(n4279), .Q(n_T_427[1884]) );
  DFFX1_LVT u_T_427_reg_0__0_ ( .D(n4316), .CLK(n4279), .Q(n_T_427[1882]), 
        .QN(n3490) );
  DFFX1_LVT u_T_427_reg_1__63_ ( .D(n4494), .CLK(n4278), .QN(n3170) );
  DFFX1_LVT u_T_427_reg_1__62_ ( .D(n4491), .CLK(n4278), .QN(n3169) );
  DFFX1_LVT u_T_427_reg_1__61_ ( .D(n4488), .CLK(n4278), .QN(n3167) );
  DFFX1_LVT u_T_427_reg_1__60_ ( .D(n4485), .CLK(n4278), .Q(n_T_427[1881]), 
        .QN(n3409) );
  DFFX1_LVT u_T_427_reg_1__59_ ( .D(n4482), .CLK(n4277), .QN(n3165) );
  DFFX1_LVT u_T_427_reg_1__58_ ( .D(n4481), .CLK(n4277), .QN(n3164) );
  DFFX1_LVT u_T_427_reg_1__57_ ( .D(n4476), .CLK(n4277), .QN(n3163) );
  DFFX1_LVT u_T_427_reg_1__56_ ( .D(n4475), .CLK(n4277), .QN(n3162) );
  DFFX1_LVT u_T_427_reg_1__55_ ( .D(n4470), .CLK(n4277), .QN(n3160) );
  DFFX1_LVT u_T_427_reg_1__54_ ( .D(n4469), .CLK(n4277), .QN(n3159) );
  DFFX1_LVT u_T_427_reg_1__53_ ( .D(n4464), .CLK(n4277), .QN(n3158) );
  DFFX1_LVT u_T_427_reg_1__52_ ( .D(n4463), .CLK(n4277), .QN(n3157) );
  DFFX1_LVT u_T_427_reg_1__51_ ( .D(n4460), .CLK(n4277), .QN(n3156) );
  DFFX1_LVT u_T_427_reg_1__50_ ( .D(n4455), .CLK(n4277), .QN(n3155) );
  DFFX1_LVT u_T_427_reg_1__49_ ( .D(n4454), .CLK(n4277), .QN(n3154) );
  DFFX1_LVT u_T_427_reg_1__48_ ( .D(n4449), .CLK(n4277), .QN(n3153) );
  DFFX1_LVT u_T_427_reg_1__47_ ( .D(n4446), .CLK(n4276), .QN(n3152) );
  DFFX1_LVT u_T_427_reg_1__45_ ( .D(n4442), .CLK(n4276), .QN(n3151) );
  DFFX1_LVT u_T_427_reg_1__43_ ( .D(n4436), .CLK(n4276), .QN(n3150) );
  DFFX1_LVT u_T_427_reg_1__42_ ( .D(n4433), .CLK(n4276), .QN(n3149) );
  DFFX1_LVT u_T_427_reg_1__41_ ( .D(n4430), .CLK(n4276), .QN(n3148) );
  DFFX1_LVT u_T_427_reg_1__40_ ( .D(n4425), .CLK(n4276), .QN(n3147) );
  DFFX1_LVT u_T_427_reg_1__37_ ( .D(n4417), .CLK(n4276), .QN(n3146) );
  DFFX1_LVT u_T_427_reg_1__36_ ( .D(n4416), .CLK(n4276), .QN(n3145) );
  DFFX1_LVT u_T_427_reg_1__32_ ( .D(n4404), .CLK(n4275), .QN(n3144) );
  DFFX1_LVT u_T_427_reg_1__30_ ( .D(n4401), .CLK(n4275), .QN(n3140) );
  DFFX1_LVT u_T_427_reg_1__29_ ( .D(n4398), .CLK(n4275), .Q(n_T_427[1872]), 
        .QN(n3375) );
  DFFX1_LVT u_T_427_reg_1__27_ ( .D(n4391), .CLK(n4275), .Q(n_T_427[1870]), 
        .QN(n3330) );
  DFFX1_LVT u_T_427_reg_1__24_ ( .D(n4386), .CLK(n4275), .QN(n3137) );
  DFFX1_LVT u_T_427_reg_1__20_ ( .D(n4376), .CLK(n4274), .Q(n_T_427[1865]), 
        .QN(n3322) );
  DFFX1_LVT u_T_427_reg_1__19_ ( .D(n4373), .CLK(n4274), .Q(n_T_427[1864]), 
        .QN(n3319) );
  DFFX1_LVT u_T_427_reg_1__18_ ( .D(n4370), .CLK(n4274), .Q(n_T_427[1863]), 
        .QN(n3316) );
  DFFX1_LVT u_T_427_reg_1__17_ ( .D(n4365), .CLK(n4274), .QN(n3139) );
  DFFX1_LVT u_T_427_reg_1__16_ ( .D(n4362), .CLK(n4274), .Q(n_T_427[1862]), 
        .QN(n3178) );
  DFFX1_LVT u_T_427_reg_1__15_ ( .D(n4360), .CLK(n4274), .Q(n_T_427[1861]) );
  DFFX1_LVT u_T_427_reg_1__14_ ( .D(n4357), .CLK(n4274), .Q(n_T_427[1860]) );
  DFFX1_LVT u_T_427_reg_1__13_ ( .D(n4355), .CLK(n4274), .Q(n_T_427[1859]) );
  DFFX1_LVT u_T_427_reg_1__12_ ( .D(n4352), .CLK(n4274), .Q(n_T_427[1858]) );
  DFFX1_LVT u_T_427_reg_1__11_ ( .D(n4351), .CLK(n4273), .Q(n_T_427[1857]) );
  DFFX1_LVT u_T_427_reg_1__10_ ( .D(n4346), .CLK(n4273), .Q(n_T_427[1856]) );
  DFFX1_LVT u_T_427_reg_1__9_ ( .D(n4343), .CLK(n4273), .Q(n_T_427[1855]) );
  DFFX1_LVT u_T_427_reg_1__8_ ( .D(n4340), .CLK(n4273), .Q(n_T_427[1854]) );
  DFFX1_LVT u_T_427_reg_1__7_ ( .D(n4337), .CLK(n4273), .Q(n_T_427[1853]) );
  DFFX1_LVT u_T_427_reg_1__6_ ( .D(n4334), .CLK(n4273), .Q(n_T_427[1852]) );
  DFFX1_LVT u_T_427_reg_1__5_ ( .D(n4331), .CLK(n4273), .Q(n_T_427[1851]) );
  DFFX1_LVT u_T_427_reg_1__4_ ( .D(n4328), .CLK(n4273), .Q(n_T_427[1850]) );
  DFFX1_LVT u_T_427_reg_1__3_ ( .D(n4325), .CLK(n4273), .Q(n_T_427[1849]) );
  DFFX1_LVT u_T_427_reg_1__2_ ( .D(n4322), .CLK(n4273), .Q(n_T_427[1848]) );
  DFFX1_LVT u_T_427_reg_1__1_ ( .D(n4321), .CLK(n4273), .QN(n3654) );
  DFFX1_LVT u_T_427_reg_1__0_ ( .D(n4318), .CLK(n4273), .QN(n3633) );
  DFFX1_LVT u_T_427_reg_2__63_ ( .D(n4494), .CLK(n4272), .QN(n3171) );
  DFFX1_LVT u_T_427_reg_2__62_ ( .D(n4491), .CLK(n4272), .Q(n_T_427[1847]), 
        .QN(n3411) );
  DFFX1_LVT u_T_427_reg_2__61_ ( .D(n4488), .CLK(n4272), .QN(n3168) );
  DFFX1_LVT u_T_427_reg_2__60_ ( .D(n4485), .CLK(n4272), .Q(n_T_427[1846]), 
        .QN(n3410) );
  DFFX1_LVT u_T_427_reg_2__59_ ( .D(n4482), .CLK(n4271), .QN(n3166) );
  DFFX1_LVT u_T_427_reg_2__58_ ( .D(n4481), .CLK(n4271), .Q(n_T_427[1845]), 
        .QN(n3474) );
  DFFX1_LVT u_T_427_reg_2__56_ ( .D(n4475), .CLK(n4271), .Q(n_T_427[1843]), 
        .QN(n3472) );
  DFFX1_LVT u_T_427_reg_2__55_ ( .D(n4470), .CLK(n4271), .QN(n3161) );
  DFFX1_LVT u_T_427_reg_2__54_ ( .D(n4469), .CLK(n4271), .Q(n_T_427[1842]), 
        .QN(n3471) );
  DFFX1_LVT u_T_427_reg_2__52_ ( .D(n4463), .CLK(n4271), .Q(n_T_427[1840]), 
        .QN(n3469) );
  DFFX1_LVT u_T_427_reg_2__51_ ( .D(n4460), .CLK(n4271), .Q(n_T_427[1839]), 
        .QN(n3412) );
  DFFX1_LVT u_T_427_reg_2__49_ ( .D(n4454), .CLK(n4271), .Q(n_T_427[1837]), 
        .QN(n3468) );
  DFFX1_LVT u_T_427_reg_2__45_ ( .D(n4442), .CLK(n4270), .Q(n_T_427[1833]), 
        .QN(n3413) );
  DFFX1_LVT u_T_427_reg_2__43_ ( .D(n4436), .CLK(n4270), .Q(n_T_427[1831]), 
        .QN(n3464) );
  DFFX1_LVT u_T_427_reg_2__42_ ( .D(n4433), .CLK(n4270), .Q(n_T_427[1830]), 
        .QN(n3462) );
  DFFX1_LVT u_T_427_reg_2__41_ ( .D(n4430), .CLK(n4270), .Q(n_T_427[1829]), 
        .QN(n3475) );
  DFFX1_LVT u_T_427_reg_2__36_ ( .D(n4416), .CLK(n4270), .Q(n_T_427[1824]), 
        .QN(n3454) );
  DFFX1_LVT u_T_427_reg_2__32_ ( .D(n4404), .CLK(n4269), .QN(n3143) );
  DFFX1_LVT u_T_427_reg_2__30_ ( .D(n4401), .CLK(n4269), .Q(n_T_427[1819]), 
        .QN(n3451) );
  DFFX1_LVT u_T_427_reg_2__29_ ( .D(n4398), .CLK(n4269), .Q(n_T_427[1818]), 
        .QN(n3396) );
  DFFX1_LVT u_T_427_reg_2__27_ ( .D(n4391), .CLK(n4269), .Q(n_T_427[1816]), 
        .QN(n3450) );
  DFFX1_LVT u_T_427_reg_2__24_ ( .D(n4386), .CLK(n4269), .Q(n_T_427[1813]), 
        .QN(n3449) );
  DFFX1_LVT u_T_427_reg_2__20_ ( .D(n4376), .CLK(n4268), .Q(n_T_427[1809]), 
        .QN(n3447) );
  DFFX1_LVT u_T_427_reg_2__19_ ( .D(n4373), .CLK(n4268), .Q(n_T_427[1808]), 
        .QN(n3446) );
  DFFX1_LVT u_T_427_reg_2__18_ ( .D(n4370), .CLK(n4268), .Q(n_T_427[1807]), 
        .QN(n3445) );
  DFFX1_LVT u_T_427_reg_2__17_ ( .D(n4365), .CLK(n4268), .QN(n3142) );
  DFFX1_LVT u_T_427_reg_2__15_ ( .D(n4360), .CLK(n4268), .Q(n_T_427[1805]) );
  DFFX1_LVT u_T_427_reg_2__14_ ( .D(n4357), .CLK(n4268), .Q(n_T_427[1804]) );
  DFFX1_LVT u_T_427_reg_2__13_ ( .D(n4355), .CLK(n4268), .Q(n_T_427[1803]) );
  DFFX1_LVT u_T_427_reg_2__12_ ( .D(n4352), .CLK(n4268), .Q(n_T_427[1802]) );
  DFFX1_LVT u_T_427_reg_2__11_ ( .D(n4351), .CLK(n4267), .Q(n_T_427[1801]) );
  DFFX1_LVT u_T_427_reg_2__10_ ( .D(n4346), .CLK(n4267), .Q(n_T_427[1800]) );
  DFFX1_LVT u_T_427_reg_2__9_ ( .D(n4343), .CLK(n4267), .Q(n_T_427[1799]) );
  DFFX1_LVT u_T_427_reg_2__8_ ( .D(n4340), .CLK(n4267), .Q(n_T_427[1798]) );
  DFFX1_LVT u_T_427_reg_2__7_ ( .D(n4337), .CLK(n4267), .Q(n_T_427[1797]) );
  DFFX1_LVT u_T_427_reg_2__6_ ( .D(n4334), .CLK(n4267), .Q(n_T_427[1796]) );
  DFFX1_LVT u_T_427_reg_2__5_ ( .D(n4331), .CLK(n4267), .Q(n_T_427[1795]) );
  DFFX1_LVT u_T_427_reg_2__4_ ( .D(n4328), .CLK(n4267), .Q(n_T_427[1794]) );
  DFFX1_LVT u_T_427_reg_2__3_ ( .D(n4325), .CLK(n4267), .Q(n_T_427[1793]) );
  DFFX1_LVT u_T_427_reg_2__2_ ( .D(n4322), .CLK(n4267), .Q(n_T_427[1792]) );
  DFFX1_LVT u_T_427_reg_2__1_ ( .D(n4321), .CLK(n4267), .QN(n3138) );
  DFFX1_LVT u_T_427_reg_2__0_ ( .D(n4318), .CLK(n4267), .Q(n_T_427[1791]), 
        .QN(n3311) );
  DFFX1_LVT u_T_427_reg_3__63_ ( .D(n4494), .CLK(n4266), .Q(n_T_427[1790]), 
        .QN(n3488) );
  DFFX1_LVT u_T_427_reg_3__62_ ( .D(n4491), .CLK(n4266), .Q(n_T_427[1789]), 
        .QN(n3487) );
  DFFX1_LVT u_T_427_reg_3__61_ ( .D(n4488), .CLK(n4266), .Q(n_T_427[1788]), 
        .QN(n3485) );
  DFFX1_LVT u_T_427_reg_3__60_ ( .D(n4485), .CLK(n4266), .Q(n_T_427[1787]) );
  DFFX1_LVT u_T_427_reg_3__58_ ( .D(n4481), .CLK(n4265), .Q(n_T_427[1785]), 
        .QN(n3516) );
  DFFX1_LVT u_T_427_reg_3__56_ ( .D(n4475), .CLK(n4265), .Q(n_T_427[1783]), 
        .QN(n3514) );
  DFFX1_LVT u_T_427_reg_3__54_ ( .D(n4469), .CLK(n4265), .Q(n_T_427[1781]), 
        .QN(n3511) );
  DFFX1_LVT u_T_427_reg_3__52_ ( .D(n4463), .CLK(n4265), .Q(n_T_427[1779]), 
        .QN(n3509) );
  DFFX1_LVT u_T_427_reg_3__51_ ( .D(n4460), .CLK(n4265), .Q(n_T_427[1778]), 
        .QN(n3508) );
  DFFX1_LVT u_T_427_reg_3__49_ ( .D(n4454), .CLK(n4265), .Q(n_T_427[1776]), 
        .QN(n3506) );
  DFFX1_LVT u_T_427_reg_3__46_ ( .D(n4443), .CLK(n4264), .Q(n_T_427[1773]) );
  DFFX1_LVT u_T_427_reg_3__45_ ( .D(n4442), .CLK(n4264), .Q(n_T_427[1772]), 
        .QN(n3503) );
  DFFX1_LVT u_T_427_reg_3__44_ ( .D(n4437), .CLK(n4264), .Q(n_T_427[1771]) );
  DFFX1_LVT u_T_427_reg_3__43_ ( .D(n4436), .CLK(n4264), .Q(n_T_427[1770]), 
        .QN(n3502) );
  DFFX1_LVT u_T_427_reg_3__42_ ( .D(n4433), .CLK(n4264), .Q(n_T_427[1769]), 
        .QN(n3501) );
  DFFX1_LVT u_T_427_reg_3__41_ ( .D(n4430), .CLK(n4264), .Q(n_T_427[1768]), 
        .QN(n3500) );
  DFFX1_LVT u_T_427_reg_3__39_ ( .D(n4422), .CLK(n4264), .Q(n_T_427[1766]) );
  DFFX1_LVT u_T_427_reg_3__38_ ( .D(n4420), .CLK(n4264), .Q(n_T_427[1765]) );
  DFFX1_LVT u_T_427_reg_3__36_ ( .D(n4416), .CLK(n4264), .Q(n_T_427[1763]), 
        .QN(n3497) );
  DFFX1_LVT u_T_427_reg_3__35_ ( .D(n4412), .CLK(n4263), .Q(n_T_427[1762]) );
  DFFX1_LVT u_T_427_reg_3__34_ ( .D(n4409), .CLK(n4263), .Q(n_T_427[1761]) );
  DFFX1_LVT u_T_427_reg_3__33_ ( .D(n4407), .CLK(n4263), .Q(n_T_427[1760]) );
  DFFX1_LVT u_T_427_reg_3__31_ ( .D(n4402), .CLK(n4263), .Q(n_T_427[1758]) );
  DFFX1_LVT u_T_427_reg_3__30_ ( .D(n4401), .CLK(n4263), .Q(n_T_427[1757]), 
        .QN(n3548) );
  DFFX1_LVT u_T_427_reg_3__29_ ( .D(n4398), .CLK(n4263), .Q(n_T_427[1756]) );
  DFFX1_LVT u_T_427_reg_3__28_ ( .D(n4394), .CLK(n4263), .Q(n_T_427[1755]) );
  DFFX1_LVT u_T_427_reg_3__27_ ( .D(n4391), .CLK(n4263), .Q(n_T_427[1754]) );
  DFFX1_LVT u_T_427_reg_3__26_ ( .D(n4389), .CLK(n4263), .Q(n_T_427[1753]) );
  DFFX1_LVT u_T_427_reg_3__25_ ( .D(n4387), .CLK(n4263), .Q(n_T_427[1752]) );
  DFFX1_LVT u_T_427_reg_3__24_ ( .D(n4386), .CLK(n4263), .Q(n_T_427[1751]), 
        .QN(n3546) );
  DFFX1_LVT u_T_427_reg_3__23_ ( .D(n4381), .CLK(n4262), .Q(n_T_427[1750]) );
  DFFX1_LVT u_T_427_reg_3__22_ ( .D(n4379), .CLK(n4262), .Q(n_T_427[1749]) );
  DFFX1_LVT u_T_427_reg_3__21_ ( .D(n4377), .CLK(n4262), .Q(n_T_427[1748]) );
  DFFX1_LVT u_T_427_reg_3__20_ ( .D(n4376), .CLK(n4262), .Q(n_T_427[1747]) );
  DFFX1_LVT u_T_427_reg_3__19_ ( .D(n4373), .CLK(n4262), .Q(n_T_427[1746]) );
  DFFX1_LVT u_T_427_reg_3__18_ ( .D(n4370), .CLK(n4262), .Q(n_T_427[1745]) );
  DFFX1_LVT u_T_427_reg_3__16_ ( .D(n4362), .CLK(n4262), .Q(n_T_427[1743]) );
  DFFX1_LVT u_T_427_reg_3__15_ ( .D(n4360), .CLK(n4262), .Q(n_T_427[1742]) );
  DFFX1_LVT u_T_427_reg_3__14_ ( .D(n4357), .CLK(n4262), .Q(n_T_427[1741]) );
  DFFX1_LVT u_T_427_reg_3__13_ ( .D(n4355), .CLK(n4262), .Q(n_T_427[1740]) );
  DFFX1_LVT u_T_427_reg_3__12_ ( .D(n4352), .CLK(n4262), .Q(n_T_427[1739]) );
  DFFX1_LVT u_T_427_reg_3__11_ ( .D(n4351), .CLK(n4261), .Q(n_T_427[1738]) );
  DFFX1_LVT u_T_427_reg_3__10_ ( .D(n4346), .CLK(n4261), .Q(n_T_427[1737]) );
  DFFX1_LVT u_T_427_reg_3__9_ ( .D(n4343), .CLK(n4261), .Q(n_T_427[1736]) );
  DFFX1_LVT u_T_427_reg_3__8_ ( .D(n4340), .CLK(n4261), .Q(n_T_427[1735]) );
  DFFX1_LVT u_T_427_reg_3__7_ ( .D(n4337), .CLK(n4261), .Q(n_T_427[1734]) );
  DFFX1_LVT u_T_427_reg_3__6_ ( .D(n4334), .CLK(n4261), .Q(n_T_427[1733]) );
  DFFX1_LVT u_T_427_reg_3__5_ ( .D(n4331), .CLK(n4261), .Q(n_T_427[1732]) );
  DFFX1_LVT u_T_427_reg_3__4_ ( .D(n4328), .CLK(n4261), .Q(n_T_427[1731]) );
  DFFX1_LVT u_T_427_reg_3__3_ ( .D(n4325), .CLK(n4261), .Q(n_T_427[1730]) );
  DFFX1_LVT u_T_427_reg_3__2_ ( .D(n4322), .CLK(n4261), .Q(n_T_427[1729]) );
  DFFX1_LVT u_T_427_reg_3__1_ ( .D(n4321), .CLK(n4261), .Q(n_T_427[1728]), 
        .QN(n3257) );
  DFFX1_LVT u_T_427_reg_3__0_ ( .D(n4318), .CLK(n4261), .Q(n_T_427[1727]), 
        .QN(n3256) );
  DFFX1_LVT u_T_427_reg_4__63_ ( .D(n4494), .CLK(n4260), .Q(n_T_427[1726]), 
        .QN(n3489) );
  DFFX1_LVT u_T_427_reg_4__62_ ( .D(n4491), .CLK(n4260), .Q(n_T_427[1725]) );
  DFFX1_LVT u_T_427_reg_4__61_ ( .D(n4488), .CLK(n4260), .Q(n_T_427[1724]), 
        .QN(n3486) );
  DFFX1_LVT u_T_427_reg_4__60_ ( .D(n4485), .CLK(n4260), .Q(n_T_427[1723]) );
  DFFX1_LVT u_T_427_reg_4__58_ ( .D(n4481), .CLK(n4259), .Q(n_T_427[1721]) );
  DFFX1_LVT u_T_427_reg_4__57_ ( .D(n4476), .CLK(n4259), .Q(n_T_427[1720]) );
  DFFX1_LVT u_T_427_reg_4__56_ ( .D(n4475), .CLK(n4259), .Q(n_T_427[1719]) );
  DFFX1_LVT u_T_427_reg_4__54_ ( .D(n4469), .CLK(n4259), .Q(n_T_427[1717]) );
  DFFX1_LVT u_T_427_reg_4__53_ ( .D(n4464), .CLK(n4259), .Q(n_T_427[1716]) );
  DFFX1_LVT u_T_427_reg_4__52_ ( .D(n4463), .CLK(n4259), .Q(n_T_427[1715]) );
  DFFX1_LVT u_T_427_reg_4__51_ ( .D(n4460), .CLK(n4259), .Q(n_T_427[1714]) );
  DFFX1_LVT u_T_427_reg_4__50_ ( .D(n4455), .CLK(n4259), .Q(n_T_427[1713]) );
  DFFX1_LVT u_T_427_reg_4__49_ ( .D(n4454), .CLK(n4259), .Q(n_T_427[1712]) );
  DFFX1_LVT u_T_427_reg_4__48_ ( .D(n4449), .CLK(n4259), .Q(n_T_427[1711]) );
  DFFX1_LVT u_T_427_reg_4__47_ ( .D(n4446), .CLK(n4258), .Q(n_T_427[1710]) );
  DFFX1_LVT u_T_427_reg_4__46_ ( .D(n4443), .CLK(n4258), .Q(n_T_427[1709]) );
  DFFX1_LVT u_T_427_reg_4__45_ ( .D(n4442), .CLK(n4258), .Q(n_T_427[1708]) );
  DFFX1_LVT u_T_427_reg_4__44_ ( .D(n4437), .CLK(n4258), .Q(n_T_427[1707]) );
  DFFX1_LVT u_T_427_reg_4__43_ ( .D(n4436), .CLK(n4258), .Q(n_T_427[1706]) );
  DFFX1_LVT u_T_427_reg_4__42_ ( .D(n4433), .CLK(n4258), .Q(n_T_427[1705]) );
  DFFX1_LVT u_T_427_reg_4__41_ ( .D(n4430), .CLK(n4258), .Q(n_T_427[1704]), 
        .QN(n2980) );
  DFFX1_LVT u_T_427_reg_4__40_ ( .D(n4425), .CLK(n4258), .Q(n_T_427[1703]) );
  DFFX1_LVT u_T_427_reg_4__39_ ( .D(n4422), .CLK(n4258), .Q(n_T_427[1702]) );
  DFFX1_LVT u_T_427_reg_4__37_ ( .D(n4417), .CLK(n4258), .Q(n_T_427[1700]) );
  DFFX1_LVT u_T_427_reg_4__36_ ( .D(n4416), .CLK(n4258), .Q(n_T_427[1699]) );
  DFFX1_LVT u_T_427_reg_4__35_ ( .D(n4412), .CLK(n4257), .Q(n_T_427[1698]) );
  DFFX1_LVT u_T_427_reg_4__34_ ( .D(n4409), .CLK(n4257), .Q(n_T_427[1697]) );
  DFFX1_LVT u_T_427_reg_4__31_ ( .D(n4402), .CLK(n4257), .Q(n_T_427[1694]) );
  DFFX1_LVT u_T_427_reg_4__30_ ( .D(n4401), .CLK(n4257), .Q(n_T_427[1693]) );
  DFFX1_LVT u_T_427_reg_4__29_ ( .D(n4398), .CLK(n4257), .Q(n_T_427[1692]) );
  DFFX1_LVT u_T_427_reg_4__28_ ( .D(n4394), .CLK(n4257), .Q(n_T_427[1691]) );
  DFFX1_LVT u_T_427_reg_4__27_ ( .D(n4391), .CLK(n4257), .Q(n_T_427[1690]) );
  DFFX1_LVT u_T_427_reg_4__26_ ( .D(n4389), .CLK(n4257), .Q(n_T_427[1689]) );
  DFFX1_LVT u_T_427_reg_4__25_ ( .D(n4387), .CLK(n4257), .Q(n_T_427[1688]) );
  DFFX1_LVT u_T_427_reg_4__24_ ( .D(n4386), .CLK(n4257), .Q(n_T_427[1687]) );
  DFFX1_LVT u_T_427_reg_4__23_ ( .D(n4381), .CLK(n4256), .Q(n_T_427[1686]) );
  DFFX1_LVT u_T_427_reg_4__22_ ( .D(n4379), .CLK(n4256), .Q(n_T_427[1685]) );
  DFFX1_LVT u_T_427_reg_4__21_ ( .D(n4377), .CLK(n4256), .Q(n_T_427[1684]) );
  DFFX1_LVT u_T_427_reg_4__20_ ( .D(n4376), .CLK(n4256), .Q(n_T_427[1683]) );
  DFFX1_LVT u_T_427_reg_4__19_ ( .D(n4373), .CLK(n4256), .Q(n_T_427[1682]) );
  DFFX1_LVT u_T_427_reg_4__18_ ( .D(n4370), .CLK(n4256), .Q(n_T_427[1681]) );
  DFFX1_LVT u_T_427_reg_4__16_ ( .D(n4362), .CLK(n4256), .Q(n_T_427[1679]) );
  DFFX1_LVT u_T_427_reg_4__11_ ( .D(n4351), .CLK(n4255), .Q(n_T_427[1674]), 
        .QN(n3435) );
  DFFX1_LVT u_T_427_reg_4__1_ ( .D(n4321), .CLK(n4255), .Q(n_T_427[1664]) );
  DFFX1_LVT u_T_427_reg_4__0_ ( .D(n4318), .CLK(n4255), .Q(n_T_427[1663]) );
  DFFX1_LVT u_T_427_reg_5__63_ ( .D(n4494), .CLK(n4254), .Q(n_T_427[1662]) );
  DFFX1_LVT u_T_427_reg_5__62_ ( .D(n4491), .CLK(n4254), .Q(n_T_427[1661]) );
  DFFX1_LVT u_T_427_reg_5__61_ ( .D(n4488), .CLK(n4254), .Q(n_T_427[1660]) );
  DFFX1_LVT u_T_427_reg_5__60_ ( .D(n4485), .CLK(n4254), .Q(n_T_427[1659]) );
  DFFX1_LVT u_T_427_reg_5__59_ ( .D(n4482), .CLK(n4253), .Q(n_T_427[1658]) );
  DFFX1_LVT u_T_427_reg_5__58_ ( .D(n4481), .CLK(n4253), .Q(n_T_427[1657]) );
  DFFX1_LVT u_T_427_reg_5__57_ ( .D(n4476), .CLK(n4253), .Q(n_T_427[1656]) );
  DFFX1_LVT u_T_427_reg_5__56_ ( .D(n4475), .CLK(n4253), .Q(n_T_427[1655]) );
  DFFX1_LVT u_T_427_reg_5__55_ ( .D(n4470), .CLK(n4253), .Q(n_T_427[1654]) );
  DFFX1_LVT u_T_427_reg_5__54_ ( .D(n4469), .CLK(n4253), .Q(n_T_427[1653]) );
  DFFX1_LVT u_T_427_reg_5__53_ ( .D(n4464), .CLK(n4253), .Q(n_T_427[1652]) );
  DFFX1_LVT u_T_427_reg_5__52_ ( .D(n4463), .CLK(n4253), .Q(n_T_427[1651]) );
  DFFX1_LVT u_T_427_reg_5__51_ ( .D(n4460), .CLK(n4253), .Q(n_T_427[1650]) );
  DFFX1_LVT u_T_427_reg_5__50_ ( .D(n4455), .CLK(n4253), .Q(n_T_427[1649]) );
  DFFX1_LVT u_T_427_reg_5__49_ ( .D(n4454), .CLK(n4253), .Q(n_T_427[1648]) );
  DFFX1_LVT u_T_427_reg_5__48_ ( .D(n4449), .CLK(n4253), .Q(n_T_427[1647]) );
  DFFX1_LVT u_T_427_reg_5__47_ ( .D(n4446), .CLK(n4252), .Q(n_T_427[1646]) );
  DFFX1_LVT u_T_427_reg_5__46_ ( .D(n4443), .CLK(n4252), .Q(n_T_427[1645]) );
  DFFX1_LVT u_T_427_reg_5__45_ ( .D(n4442), .CLK(n4252), .Q(n_T_427[1644]) );
  DFFX1_LVT u_T_427_reg_5__44_ ( .D(n4437), .CLK(n4252), .Q(n_T_427[1643]) );
  DFFX1_LVT u_T_427_reg_5__43_ ( .D(n4436), .CLK(n4252), .Q(n_T_427[1642]) );
  DFFX1_LVT u_T_427_reg_5__42_ ( .D(n4433), .CLK(n4252), .Q(n_T_427[1641]) );
  DFFX1_LVT u_T_427_reg_5__41_ ( .D(n4430), .CLK(n4252), .Q(n_T_427[1640]) );
  DFFX1_LVT u_T_427_reg_5__40_ ( .D(n4425), .CLK(n4252), .Q(n_T_427[1639]) );
  DFFX1_LVT u_T_427_reg_5__39_ ( .D(n4422), .CLK(n4252), .Q(n_T_427[1638]) );
  DFFX1_LVT u_T_427_reg_5__38_ ( .D(n4420), .CLK(n4252), .Q(n_T_427[1637]) );
  DFFX1_LVT u_T_427_reg_5__37_ ( .D(n4417), .CLK(n4252), .Q(n_T_427[1636]) );
  DFFX1_LVT u_T_427_reg_5__36_ ( .D(n4416), .CLK(n4252), .Q(n_T_427[1635]) );
  DFFX1_LVT u_T_427_reg_5__35_ ( .D(n4412), .CLK(n4251), .Q(n_T_427[1634]) );
  DFFX1_LVT u_T_427_reg_5__34_ ( .D(n4409), .CLK(n4251), .Q(n_T_427[1633]) );
  DFFX1_LVT u_T_427_reg_5__33_ ( .D(n4407), .CLK(n4251), .Q(n_T_427[1632]) );
  DFFX1_LVT u_T_427_reg_5__32_ ( .D(n4404), .CLK(n4251), .Q(n_T_427[1631]) );
  DFFX1_LVT u_T_427_reg_5__31_ ( .D(n4402), .CLK(n4251), .Q(n_T_427[1630]) );
  DFFX1_LVT u_T_427_reg_5__30_ ( .D(n4401), .CLK(n4251), .Q(n_T_427[1629]) );
  DFFX1_LVT u_T_427_reg_5__29_ ( .D(n4398), .CLK(n4251), .Q(n_T_427[1628]) );
  DFFX1_LVT u_T_427_reg_5__28_ ( .D(n4394), .CLK(n4251), .Q(n_T_427[1627]) );
  DFFX1_LVT u_T_427_reg_5__27_ ( .D(n4391), .CLK(n4251), .Q(n_T_427[1626]) );
  DFFX1_LVT u_T_427_reg_5__26_ ( .D(n4389), .CLK(n4251), .Q(n_T_427[1625]) );
  DFFX1_LVT u_T_427_reg_5__25_ ( .D(n4387), .CLK(n4251), .Q(n_T_427[1624]) );
  DFFX1_LVT u_T_427_reg_5__24_ ( .D(n4386), .CLK(n4251), .Q(n_T_427[1623]) );
  DFFX1_LVT u_T_427_reg_5__23_ ( .D(n4381), .CLK(n4250), .Q(n_T_427[1622]) );
  DFFX1_LVT u_T_427_reg_5__22_ ( .D(n4379), .CLK(n4250), .Q(n_T_427[1621]) );
  DFFX1_LVT u_T_427_reg_5__21_ ( .D(n4377), .CLK(n4250), .Q(n_T_427[1620]) );
  DFFX1_LVT u_T_427_reg_5__20_ ( .D(n4376), .CLK(n4250), .Q(n_T_427[1619]) );
  DFFX1_LVT u_T_427_reg_5__19_ ( .D(n4373), .CLK(n4250), .Q(n_T_427[1618]) );
  DFFX1_LVT u_T_427_reg_5__18_ ( .D(n4370), .CLK(n4250), .Q(n_T_427[1617]) );
  DFFX1_LVT u_T_427_reg_5__17_ ( .D(n4365), .CLK(n4250), .Q(n_T_427[1616]) );
  DFFX1_LVT u_T_427_reg_5__16_ ( .D(n4362), .CLK(n4250), .Q(n_T_427[1615]) );
  DFFX1_LVT u_T_427_reg_5__15_ ( .D(n4360), .CLK(n4250), .Q(n_T_427[1614]) );
  DFFX1_LVT u_T_427_reg_5__14_ ( .D(n4357), .CLK(n4250), .Q(n_T_427[1613]) );
  DFFX1_LVT u_T_427_reg_5__13_ ( .D(n4355), .CLK(n4250), .Q(n_T_427[1612]) );
  DFFX1_LVT u_T_427_reg_5__12_ ( .D(n4352), .CLK(n4250), .Q(n_T_427[1611]) );
  DFFX1_LVT u_T_427_reg_5__11_ ( .D(n4351), .CLK(n4249), .Q(n_T_427[1610]) );
  DFFX1_LVT u_T_427_reg_5__10_ ( .D(n4346), .CLK(n4249), .Q(n_T_427[1609]) );
  DFFX1_LVT u_T_427_reg_5__9_ ( .D(n4343), .CLK(n4249), .Q(n_T_427[1608]) );
  DFFX1_LVT u_T_427_reg_5__8_ ( .D(n4340), .CLK(n4249), .Q(n_T_427[1607]) );
  DFFX1_LVT u_T_427_reg_5__7_ ( .D(n4337), .CLK(n4249), .Q(n_T_427[1606]) );
  DFFX1_LVT u_T_427_reg_5__6_ ( .D(n4334), .CLK(n4249), .Q(n_T_427[1605]) );
  DFFX1_LVT u_T_427_reg_5__5_ ( .D(n4331), .CLK(n4249), .Q(n_T_427[1604]) );
  DFFX1_LVT u_T_427_reg_5__4_ ( .D(n4328), .CLK(n4249), .Q(n_T_427[1603]) );
  DFFX1_LVT u_T_427_reg_5__3_ ( .D(n4325), .CLK(n4249), .Q(n_T_427[1602]) );
  DFFX1_LVT u_T_427_reg_5__2_ ( .D(n4322), .CLK(n4249), .Q(n_T_427[1601]) );
  DFFX1_LVT u_T_427_reg_5__1_ ( .D(n4321), .CLK(n4249), .Q(n_T_427[1600]) );
  DFFX1_LVT u_T_427_reg_5__0_ ( .D(n4318), .CLK(n4249), .Q(n_T_427[1599]) );
  DFFX1_LVT u_T_427_reg_6__63_ ( .D(n4494), .CLK(n4248), .Q(n_T_427[1598]) );
  DFFX1_LVT u_T_427_reg_6__62_ ( .D(n4491), .CLK(n4248), .Q(n_T_427[1597]) );
  DFFX1_LVT u_T_427_reg_6__61_ ( .D(n4488), .CLK(n4248), .Q(n_T_427[1596]) );
  DFFX1_LVT u_T_427_reg_6__60_ ( .D(n4485), .CLK(n4248), .Q(n_T_427[1595]) );
  DFFX1_LVT u_T_427_reg_6__59_ ( .D(n4482), .CLK(n4247), .Q(n_T_427[1594]) );
  DFFX1_LVT u_T_427_reg_6__58_ ( .D(n4481), .CLK(n4247), .Q(n_T_427[1593]) );
  DFFX1_LVT u_T_427_reg_6__57_ ( .D(n4476), .CLK(n4247), .Q(n_T_427[1592]) );
  DFFX1_LVT u_T_427_reg_6__56_ ( .D(n4475), .CLK(n4247), .Q(n_T_427[1591]) );
  DFFX1_LVT u_T_427_reg_6__55_ ( .D(n4470), .CLK(n4247), .Q(n_T_427[1590]) );
  DFFX1_LVT u_T_427_reg_6__54_ ( .D(n4469), .CLK(n4247), .Q(n_T_427[1589]) );
  DFFX1_LVT u_T_427_reg_6__53_ ( .D(n4464), .CLK(n4247), .Q(n_T_427[1588]) );
  DFFX1_LVT u_T_427_reg_6__52_ ( .D(n4463), .CLK(n4247), .Q(n_T_427[1587]) );
  DFFX1_LVT u_T_427_reg_6__51_ ( .D(n4460), .CLK(n4247), .Q(n_T_427[1586]) );
  DFFX1_LVT u_T_427_reg_6__50_ ( .D(n4455), .CLK(n4247), .Q(n_T_427[1585]) );
  DFFX1_LVT u_T_427_reg_6__49_ ( .D(n4454), .CLK(n4247), .Q(n_T_427[1584]) );
  DFFX1_LVT u_T_427_reg_6__48_ ( .D(n4449), .CLK(n4247), .Q(n_T_427[1583]) );
  DFFX1_LVT u_T_427_reg_6__47_ ( .D(n4446), .CLK(n4246), .Q(n_T_427[1582]) );
  DFFX1_LVT u_T_427_reg_6__46_ ( .D(n4443), .CLK(n4246), .Q(n_T_427[1581]) );
  DFFX1_LVT u_T_427_reg_6__45_ ( .D(n4442), .CLK(n4246), .Q(n_T_427[1580]) );
  DFFX1_LVT u_T_427_reg_6__44_ ( .D(n4437), .CLK(n4246), .Q(n_T_427[1579]) );
  DFFX1_LVT u_T_427_reg_6__43_ ( .D(n4436), .CLK(n4246), .Q(n_T_427[1578]) );
  DFFX1_LVT u_T_427_reg_6__42_ ( .D(n4433), .CLK(n4246), .Q(n_T_427[1577]) );
  DFFX1_LVT u_T_427_reg_6__41_ ( .D(n4430), .CLK(n4246), .Q(n_T_427[1576]) );
  DFFX1_LVT u_T_427_reg_6__40_ ( .D(n4425), .CLK(n4246), .Q(n_T_427[1575]) );
  DFFX1_LVT u_T_427_reg_6__39_ ( .D(n4422), .CLK(n4246), .Q(n_T_427[1574]) );
  DFFX1_LVT u_T_427_reg_6__38_ ( .D(n4420), .CLK(n4246), .Q(n_T_427[1573]) );
  DFFX1_LVT u_T_427_reg_6__37_ ( .D(n4417), .CLK(n4246), .Q(n_T_427[1572]) );
  DFFX1_LVT u_T_427_reg_6__36_ ( .D(n4416), .CLK(n4246), .Q(n_T_427[1571]) );
  DFFX1_LVT u_T_427_reg_6__35_ ( .D(n4412), .CLK(n4245), .Q(n_T_427[1570]) );
  DFFX1_LVT u_T_427_reg_6__34_ ( .D(n4409), .CLK(n4245), .Q(n_T_427[1569]) );
  DFFX1_LVT u_T_427_reg_6__33_ ( .D(n4407), .CLK(n4245), .Q(n_T_427[1568]) );
  DFFX1_LVT u_T_427_reg_6__32_ ( .D(n4404), .CLK(n4245), .Q(n_T_427[1567]) );
  DFFX1_LVT u_T_427_reg_6__31_ ( .D(n4402), .CLK(n4245), .Q(n_T_427[1566]) );
  DFFX1_LVT u_T_427_reg_6__30_ ( .D(n4401), .CLK(n4245), .Q(n_T_427[1565]) );
  DFFX1_LVT u_T_427_reg_6__29_ ( .D(n4398), .CLK(n4245), .Q(n_T_427[1564]) );
  DFFX1_LVT u_T_427_reg_6__28_ ( .D(n4394), .CLK(n4245), .Q(n_T_427[1563]) );
  DFFX1_LVT u_T_427_reg_6__27_ ( .D(n4391), .CLK(n4245), .Q(n_T_427[1562]) );
  DFFX1_LVT u_T_427_reg_6__26_ ( .D(n4389), .CLK(n4245), .Q(n_T_427[1561]) );
  DFFX1_LVT u_T_427_reg_6__25_ ( .D(n4387), .CLK(n4245), .Q(n_T_427[1560]) );
  DFFX1_LVT u_T_427_reg_6__24_ ( .D(n4386), .CLK(n4245), .Q(n_T_427[1559]) );
  DFFX1_LVT u_T_427_reg_6__23_ ( .D(n4381), .CLK(n4244), .Q(n_T_427[1558]) );
  DFFX1_LVT u_T_427_reg_6__22_ ( .D(n4379), .CLK(n4244), .Q(n_T_427[1557]) );
  DFFX1_LVT u_T_427_reg_6__21_ ( .D(n4377), .CLK(n4244), .Q(n_T_427[1556]) );
  DFFX1_LVT u_T_427_reg_6__20_ ( .D(n4376), .CLK(n4244), .Q(n_T_427[1555]) );
  DFFX1_LVT u_T_427_reg_6__19_ ( .D(n4373), .CLK(n4244), .Q(n_T_427[1554]) );
  DFFX1_LVT u_T_427_reg_6__18_ ( .D(n4370), .CLK(n4244), .Q(n_T_427[1553]) );
  DFFX1_LVT u_T_427_reg_6__17_ ( .D(n4365), .CLK(n4244), .Q(n_T_427[1552]) );
  DFFX1_LVT u_T_427_reg_6__16_ ( .D(n4362), .CLK(n4244), .Q(n_T_427[1551]) );
  DFFX1_LVT u_T_427_reg_6__15_ ( .D(n4360), .CLK(n4244), .Q(n_T_427[1550]) );
  DFFX1_LVT u_T_427_reg_6__14_ ( .D(n4357), .CLK(n4244), .Q(n_T_427[1549]) );
  DFFX1_LVT u_T_427_reg_6__13_ ( .D(n4355), .CLK(n4244), .Q(n_T_427[1548]) );
  DFFX1_LVT u_T_427_reg_6__12_ ( .D(n4352), .CLK(n4244), .Q(n_T_427[1547]) );
  DFFX1_LVT u_T_427_reg_6__11_ ( .D(n4351), .CLK(n4243), .Q(n_T_427[1546]) );
  DFFX1_LVT u_T_427_reg_6__10_ ( .D(n4346), .CLK(n4243), .Q(n_T_427[1545]) );
  DFFX1_LVT u_T_427_reg_6__9_ ( .D(n4343), .CLK(n4243), .Q(n_T_427[1544]) );
  DFFX1_LVT u_T_427_reg_6__8_ ( .D(n4340), .CLK(n4243), .Q(n_T_427[1543]) );
  DFFX1_LVT u_T_427_reg_6__7_ ( .D(n4337), .CLK(n4243), .Q(n_T_427[1542]) );
  DFFX1_LVT u_T_427_reg_6__6_ ( .D(n4334), .CLK(n4243), .Q(n_T_427[1541]) );
  DFFX1_LVT u_T_427_reg_6__5_ ( .D(n4331), .CLK(n4243), .Q(n_T_427[1540]) );
  DFFX1_LVT u_T_427_reg_6__4_ ( .D(n4328), .CLK(n4243), .Q(n_T_427[1539]) );
  DFFX1_LVT u_T_427_reg_6__3_ ( .D(n4325), .CLK(n4243), .Q(n_T_427[1538]) );
  DFFX1_LVT u_T_427_reg_6__2_ ( .D(n4322), .CLK(n4243), .Q(n_T_427[1537]) );
  DFFX1_LVT u_T_427_reg_6__1_ ( .D(n4321), .CLK(n4243), .Q(n_T_427[1536]) );
  DFFX1_LVT u_T_427_reg_6__0_ ( .D(n4318), .CLK(n4243), .Q(n_T_427[1535]) );
  DFFX1_LVT u_T_427_reg_7__63_ ( .D(n4494), .CLK(n4242), .Q(n_T_427[1534]) );
  DFFX1_LVT u_T_427_reg_7__62_ ( .D(n4491), .CLK(n4242), .Q(n_T_427[1533]) );
  DFFX1_LVT u_T_427_reg_7__61_ ( .D(n4488), .CLK(n4242), .Q(n_T_427[1532]) );
  DFFX1_LVT u_T_427_reg_7__60_ ( .D(n4485), .CLK(n4242), .Q(n_T_427[1531]) );
  DFFX1_LVT u_T_427_reg_7__59_ ( .D(n4482), .CLK(n4241), .Q(n_T_427[1530]) );
  DFFX1_LVT u_T_427_reg_7__58_ ( .D(n4481), .CLK(n4241), .Q(n_T_427[1529]) );
  DFFX1_LVT u_T_427_reg_7__57_ ( .D(n4476), .CLK(n4241), .Q(n_T_427[1528]) );
  DFFX1_LVT u_T_427_reg_7__56_ ( .D(n4475), .CLK(n4241), .Q(n_T_427[1527]) );
  DFFX1_LVT u_T_427_reg_7__55_ ( .D(n4470), .CLK(n4241), .Q(n_T_427[1526]) );
  DFFX1_LVT u_T_427_reg_7__54_ ( .D(n4469), .CLK(n4241), .Q(n_T_427[1525]) );
  DFFX1_LVT u_T_427_reg_7__53_ ( .D(n4464), .CLK(n4241), .Q(n_T_427[1524]) );
  DFFX1_LVT u_T_427_reg_7__52_ ( .D(n4463), .CLK(n4241), .Q(n_T_427[1523]) );
  DFFX1_LVT u_T_427_reg_7__51_ ( .D(n4460), .CLK(n4241), .Q(n_T_427[1522]) );
  DFFX1_LVT u_T_427_reg_7__50_ ( .D(n4455), .CLK(n4241), .Q(n_T_427[1521]) );
  DFFX1_LVT u_T_427_reg_7__49_ ( .D(n4454), .CLK(n4241), .Q(n_T_427[1520]) );
  DFFX1_LVT u_T_427_reg_7__48_ ( .D(n4449), .CLK(n4241), .Q(n_T_427[1519]), 
        .QN(n3774) );
  DFFX1_LVT u_T_427_reg_7__47_ ( .D(n4446), .CLK(n4240), .Q(n_T_427[1518]) );
  DFFX1_LVT u_T_427_reg_7__46_ ( .D(n4443), .CLK(n4240), .Q(n_T_427[1517]) );
  DFFX1_LVT u_T_427_reg_7__45_ ( .D(n4442), .CLK(n4240), .Q(n_T_427[1516]) );
  DFFX1_LVT u_T_427_reg_7__44_ ( .D(n4437), .CLK(n4240), .Q(n_T_427[1515]) );
  DFFX1_LVT u_T_427_reg_7__43_ ( .D(n4436), .CLK(n4240), .Q(n_T_427[1514]) );
  DFFX1_LVT u_T_427_reg_7__42_ ( .D(n4433), .CLK(n4240), .Q(n_T_427[1513]), 
        .QN(n3463) );
  DFFX1_LVT u_T_427_reg_7__41_ ( .D(n4430), .CLK(n4240), .Q(n_T_427[1512]) );
  DFFX1_LVT u_T_427_reg_7__40_ ( .D(n4425), .CLK(n4240), .Q(n_T_427[1511]) );
  DFFX1_LVT u_T_427_reg_7__37_ ( .D(n4417), .CLK(n4240), .Q(n_T_427[1508]) );
  DFFX1_LVT u_T_427_reg_7__36_ ( .D(n4416), .CLK(n4240), .Q(n_T_427[1507]), 
        .QN(n3455) );
  DFFX1_LVT u_T_427_reg_7__35_ ( .D(n4412), .CLK(n4239), .Q(n_T_427[1506]) );
  DFFX1_LVT u_T_427_reg_7__34_ ( .D(n4409), .CLK(n4239), .Q(n_T_427[1505]) );
  DFFX1_LVT u_T_427_reg_7__33_ ( .D(n4407), .CLK(n4239), .Q(n_T_427[1504]) );
  DFFX1_LVT u_T_427_reg_7__32_ ( .D(n4404), .CLK(n4239), .Q(n_T_427[1503]) );
  DFFX1_LVT u_T_427_reg_7__31_ ( .D(n4402), .CLK(n4239), .Q(n_T_427[1502]) );
  DFFX1_LVT u_T_427_reg_7__30_ ( .D(n4401), .CLK(n4239), .Q(n_T_427[1501]) );
  DFFX1_LVT u_T_427_reg_7__29_ ( .D(n4398), .CLK(n4239), .Q(n_T_427[1500]) );
  DFFX1_LVT u_T_427_reg_7__28_ ( .D(n4394), .CLK(n4239), .Q(n_T_427[1499]) );
  DFFX1_LVT u_T_427_reg_7__27_ ( .D(n4391), .CLK(n4239), .Q(n_T_427[1498]) );
  DFFX1_LVT u_T_427_reg_7__26_ ( .D(n4389), .CLK(n4239), .Q(n_T_427[1497]) );
  DFFX1_LVT u_T_427_reg_7__25_ ( .D(n4387), .CLK(n4239), .Q(n_T_427[1496]) );
  DFFX1_LVT u_T_427_reg_7__24_ ( .D(n4386), .CLK(n4239), .Q(n_T_427[1495]) );
  DFFX1_LVT u_T_427_reg_7__23_ ( .D(n4381), .CLK(n4238), .Q(n_T_427[1494]) );
  DFFX1_LVT u_T_427_reg_7__22_ ( .D(n4379), .CLK(n4238), .Q(n_T_427[1493]) );
  DFFX1_LVT u_T_427_reg_7__21_ ( .D(n4377), .CLK(n4238), .Q(n_T_427[1492]) );
  DFFX1_LVT u_T_427_reg_7__20_ ( .D(n4376), .CLK(n4238), .Q(n_T_427[1491]) );
  DFFX1_LVT u_T_427_reg_7__19_ ( .D(n4373), .CLK(n4238), .Q(n_T_427[1490]) );
  DFFX1_LVT u_T_427_reg_7__18_ ( .D(n4370), .CLK(n4238), .Q(n_T_427[1489]) );
  DFFX1_LVT u_T_427_reg_7__17_ ( .D(n4365), .CLK(n4238), .Q(n_T_427[1488]) );
  DFFX1_LVT u_T_427_reg_7__16_ ( .D(n4362), .CLK(n4238), .Q(n_T_427[1487]) );
  DFFX1_LVT u_T_427_reg_7__1_ ( .D(n4321), .CLK(n4237), .Q(n_T_427[1472]), 
        .QN(n3416) );
  DFFX1_LVT u_T_427_reg_7__0_ ( .D(n4318), .CLK(n4237), .Q(n_T_427[1471]), 
        .QN(n3417) );
  DFFX1_LVT u_T_427_reg_8__63_ ( .D(n4494), .CLK(n4236), .Q(n_T_427[1470]) );
  DFFX1_LVT u_T_427_reg_8__62_ ( .D(n4491), .CLK(n4236), .Q(n_T_427[1469]) );
  DFFX1_LVT u_T_427_reg_8__61_ ( .D(n4488), .CLK(n4236), .Q(n_T_427[1468]) );
  DFFX1_LVT u_T_427_reg_8__60_ ( .D(n4485), .CLK(n4236), .Q(n_T_427[1467]) );
  DFFX1_LVT u_T_427_reg_8__59_ ( .D(n4482), .CLK(n4235), .Q(n_T_427[1466]) );
  DFFX1_LVT u_T_427_reg_8__58_ ( .D(n4480), .CLK(n4235), .Q(n_T_427[1465]) );
  DFFX1_LVT u_T_427_reg_8__57_ ( .D(n4476), .CLK(n4235), .Q(n_T_427[1464]) );
  DFFX1_LVT u_T_427_reg_8__56_ ( .D(n4474), .CLK(n4235), .Q(n_T_427[1463]) );
  DFFX1_LVT u_T_427_reg_8__55_ ( .D(n4470), .CLK(n4235), .Q(n_T_427[1462]) );
  DFFX1_LVT u_T_427_reg_8__54_ ( .D(n4468), .CLK(n4235), .Q(n_T_427[1461]) );
  DFFX1_LVT u_T_427_reg_8__53_ ( .D(n4464), .CLK(n4235), .Q(n_T_427[1460]) );
  DFFX1_LVT u_T_427_reg_8__52_ ( .D(n4462), .CLK(n4235), .Q(n_T_427[1459]) );
  DFFX1_LVT u_T_427_reg_8__51_ ( .D(n4459), .CLK(n4235), .Q(n_T_427[1458]) );
  DFFX1_LVT u_T_427_reg_8__50_ ( .D(n4455), .CLK(n4235), .Q(n_T_427[1457]) );
  DFFX1_LVT u_T_427_reg_8__49_ ( .D(n4453), .CLK(n4235), .Q(n_T_427[1456]) );
  DFFX1_LVT u_T_427_reg_8__48_ ( .D(n4449), .CLK(n4235), .Q(n_T_427[1455]) );
  DFFX1_LVT u_T_427_reg_8__47_ ( .D(n4446), .CLK(n4234), .Q(n_T_427[1454]) );
  DFFX1_LVT u_T_427_reg_8__46_ ( .D(n4443), .CLK(n4234), .Q(n_T_427[1453]) );
  DFFX1_LVT u_T_427_reg_8__45_ ( .D(n4441), .CLK(n4234), .Q(n_T_427[1452]) );
  DFFX1_LVT u_T_427_reg_8__44_ ( .D(n4437), .CLK(n4234), .Q(n_T_427[1451]) );
  DFFX1_LVT u_T_427_reg_8__43_ ( .D(n4435), .CLK(n4234), .Q(n_T_427[1450]) );
  DFFX1_LVT u_T_427_reg_8__42_ ( .D(n4432), .CLK(n4234), .Q(n_T_427[1449]) );
  DFFX1_LVT u_T_427_reg_8__41_ ( .D(n4429), .CLK(n4234), .Q(n_T_427[1448]) );
  DFFX1_LVT u_T_427_reg_8__40_ ( .D(n4425), .CLK(n4234), .Q(n_T_427[1447]) );
  DFFX1_LVT u_T_427_reg_8__39_ ( .D(n4422), .CLK(n4234), .Q(n_T_427[1446]) );
  DFFX1_LVT u_T_427_reg_8__38_ ( .D(n4420), .CLK(n4234), .Q(n_T_427[1445]) );
  DFFX1_LVT u_T_427_reg_8__37_ ( .D(n4417), .CLK(n4234), .Q(n_T_427[1444]) );
  DFFX1_LVT u_T_427_reg_8__36_ ( .D(n4415), .CLK(n4234), .Q(n_T_427[1443]) );
  DFFX1_LVT u_T_427_reg_8__35_ ( .D(n4412), .CLK(n4233), .Q(n_T_427[1442]) );
  DFFX1_LVT u_T_427_reg_8__34_ ( .D(n4409), .CLK(n4233), .Q(n_T_427[1441]) );
  DFFX1_LVT u_T_427_reg_8__33_ ( .D(n4407), .CLK(n4233), .Q(n_T_427[1440]) );
  DFFX1_LVT u_T_427_reg_8__32_ ( .D(n4404), .CLK(n4233), .Q(n_T_427[1439]) );
  DFFX1_LVT u_T_427_reg_8__31_ ( .D(n4402), .CLK(n4233), .Q(n_T_427[1438]) );
  DFFX1_LVT u_T_427_reg_8__30_ ( .D(n4400), .CLK(n4233), .Q(n_T_427[1437]) );
  DFFX1_LVT u_T_427_reg_8__29_ ( .D(n4397), .CLK(n4233), .Q(n_T_427[1436]) );
  DFFX1_LVT u_T_427_reg_8__28_ ( .D(n4394), .CLK(n4233), .Q(n_T_427[1435]) );
  DFFX1_LVT u_T_427_reg_8__27_ ( .D(n4391), .CLK(n4233), .Q(n_T_427[1434]) );
  DFFX1_LVT u_T_427_reg_8__26_ ( .D(n4389), .CLK(n4233), .Q(n_T_427[1433]) );
  DFFX1_LVT u_T_427_reg_8__25_ ( .D(n4387), .CLK(n4233), .Q(n_T_427[1432]) );
  DFFX1_LVT u_T_427_reg_8__24_ ( .D(n4385), .CLK(n4233), .Q(n_T_427[1431]) );
  DFFX1_LVT u_T_427_reg_8__23_ ( .D(n4381), .CLK(n4232), .Q(n_T_427[1430]) );
  DFFX1_LVT u_T_427_reg_8__22_ ( .D(n4379), .CLK(n4232), .Q(n_T_427[1429]) );
  DFFX1_LVT u_T_427_reg_8__21_ ( .D(n4377), .CLK(n4232), .Q(n_T_427[1428]) );
  DFFX1_LVT u_T_427_reg_8__20_ ( .D(n4375), .CLK(n4232), .Q(n_T_427[1427]) );
  DFFX1_LVT u_T_427_reg_8__19_ ( .D(n4372), .CLK(n4232), .Q(n_T_427[1426]) );
  DFFX1_LVT u_T_427_reg_8__18_ ( .D(n4369), .CLK(n4232), .Q(n_T_427[1425]) );
  DFFX1_LVT u_T_427_reg_8__17_ ( .D(n4365), .CLK(n4232), .Q(n_T_427[1424]) );
  DFFX1_LVT u_T_427_reg_8__16_ ( .D(n4362), .CLK(n4232), .Q(n_T_427[1423]) );
  DFFX1_LVT u_T_427_reg_8__15_ ( .D(n4360), .CLK(n4232), .Q(n_T_427[1422]) );
  DFFX1_LVT u_T_427_reg_8__14_ ( .D(n4357), .CLK(n4232), .Q(n_T_427[1421]) );
  DFFX1_LVT u_T_427_reg_8__13_ ( .D(n4355), .CLK(n4232), .Q(n_T_427[1420]) );
  DFFX1_LVT u_T_427_reg_8__12_ ( .D(n4352), .CLK(n4232), .Q(n_T_427[1419]) );
  DFFX1_LVT u_T_427_reg_8__11_ ( .D(n4350), .CLK(n4231), .Q(n_T_427[1418]) );
  DFFX1_LVT u_T_427_reg_8__10_ ( .D(n4346), .CLK(n4231), .Q(n_T_427[1417]) );
  DFFX1_LVT u_T_427_reg_8__9_ ( .D(n4343), .CLK(n4231), .Q(n_T_427[1416]) );
  DFFX1_LVT u_T_427_reg_8__8_ ( .D(n4340), .CLK(n4231), .Q(n_T_427[1415]) );
  DFFX1_LVT u_T_427_reg_8__7_ ( .D(n4337), .CLK(n4231), .Q(n_T_427[1414]) );
  DFFX1_LVT u_T_427_reg_8__6_ ( .D(n4334), .CLK(n4231), .Q(n_T_427[1413]) );
  DFFX1_LVT u_T_427_reg_8__5_ ( .D(n4331), .CLK(n4231), .Q(n_T_427[1412]) );
  DFFX1_LVT u_T_427_reg_8__4_ ( .D(n4328), .CLK(n4231), .Q(n_T_427[1411]) );
  DFFX1_LVT u_T_427_reg_8__3_ ( .D(n4325), .CLK(n4231), .Q(n_T_427[1410]) );
  DFFX1_LVT u_T_427_reg_8__2_ ( .D(n4322), .CLK(n4231), .Q(n_T_427[1409]) );
  DFFX1_LVT u_T_427_reg_8__1_ ( .D(n4320), .CLK(n4231), .Q(n_T_427[1408]) );
  DFFX1_LVT u_T_427_reg_8__0_ ( .D(n4317), .CLK(n4231), .Q(n_T_427[1407]) );
  DFFX1_LVT u_T_427_reg_9__63_ ( .D(n4494), .CLK(n4230), .Q(n_T_427[1406]) );
  DFFX1_LVT u_T_427_reg_9__62_ ( .D(n4491), .CLK(n4230), .Q(n_T_427[1405]) );
  DFFX1_LVT u_T_427_reg_9__61_ ( .D(n4488), .CLK(n4230), .Q(n_T_427[1404]) );
  DFFX1_LVT u_T_427_reg_9__60_ ( .D(n4485), .CLK(n4230), .Q(n_T_427[1403]) );
  DFFX1_LVT u_T_427_reg_9__59_ ( .D(n4482), .CLK(n4229), .Q(n_T_427[1402]) );
  DFFX1_LVT u_T_427_reg_9__58_ ( .D(n4480), .CLK(n4229), .Q(n_T_427[1401]) );
  DFFX1_LVT u_T_427_reg_9__57_ ( .D(n4476), .CLK(n4229), .Q(n_T_427[1400]) );
  DFFX1_LVT u_T_427_reg_9__56_ ( .D(n4474), .CLK(n4229), .Q(n_T_427[1399]) );
  DFFX1_LVT u_T_427_reg_9__55_ ( .D(n4470), .CLK(n4229), .Q(n_T_427[1398]) );
  DFFX1_LVT u_T_427_reg_9__54_ ( .D(n4468), .CLK(n4229), .Q(n_T_427[1397]) );
  DFFX1_LVT u_T_427_reg_9__53_ ( .D(n4464), .CLK(n4229), .Q(n_T_427[1396]) );
  DFFX1_LVT u_T_427_reg_9__52_ ( .D(n4462), .CLK(n4229), .Q(n_T_427[1395]) );
  DFFX1_LVT u_T_427_reg_9__51_ ( .D(n4459), .CLK(n4229), .Q(n_T_427[1394]) );
  DFFX1_LVT u_T_427_reg_9__50_ ( .D(n4455), .CLK(n4229), .Q(n_T_427[1393]) );
  DFFX1_LVT u_T_427_reg_9__49_ ( .D(n4453), .CLK(n4229), .Q(n_T_427[1392]) );
  DFFX1_LVT u_T_427_reg_9__48_ ( .D(n4449), .CLK(n4229), .Q(n_T_427[1391]) );
  DFFX1_LVT u_T_427_reg_9__47_ ( .D(n4446), .CLK(n4228), .Q(n_T_427[1390]) );
  DFFX1_LVT u_T_427_reg_9__46_ ( .D(n4443), .CLK(n4228), .Q(n_T_427[1389]) );
  DFFX1_LVT u_T_427_reg_9__45_ ( .D(n4441), .CLK(n4228), .Q(n_T_427[1388]) );
  DFFX1_LVT u_T_427_reg_9__44_ ( .D(n4437), .CLK(n4228), .Q(n_T_427[1387]) );
  DFFX1_LVT u_T_427_reg_9__43_ ( .D(n4435), .CLK(n4228), .Q(n_T_427[1386]) );
  DFFX1_LVT u_T_427_reg_9__42_ ( .D(n4432), .CLK(n4228), .Q(n_T_427[1385]) );
  DFFX1_LVT u_T_427_reg_9__41_ ( .D(n4429), .CLK(n4228), .Q(n_T_427[1384]) );
  DFFX1_LVT u_T_427_reg_9__40_ ( .D(n4425), .CLK(n4228), .Q(n_T_427[1383]) );
  DFFX1_LVT u_T_427_reg_9__39_ ( .D(n4422), .CLK(n4228), .Q(n_T_427[1382]) );
  DFFX1_LVT u_T_427_reg_9__38_ ( .D(n4420), .CLK(n4228), .Q(n_T_427[1381]) );
  DFFX1_LVT u_T_427_reg_9__37_ ( .D(n4417), .CLK(n4228), .Q(n_T_427[1380]) );
  DFFX1_LVT u_T_427_reg_9__36_ ( .D(n4415), .CLK(n4228), .Q(n_T_427[1379]) );
  DFFX1_LVT u_T_427_reg_9__35_ ( .D(n4412), .CLK(n4227), .Q(n_T_427[1378]) );
  DFFX1_LVT u_T_427_reg_9__34_ ( .D(n4409), .CLK(n4227), .Q(n_T_427[1377]) );
  DFFX1_LVT u_T_427_reg_9__33_ ( .D(n4407), .CLK(n4227), .Q(n_T_427[1376]) );
  DFFX1_LVT u_T_427_reg_9__32_ ( .D(n4404), .CLK(n4227), .Q(n_T_427[1375]) );
  DFFX1_LVT u_T_427_reg_9__31_ ( .D(n4402), .CLK(n4227), .Q(n_T_427[1374]) );
  DFFX1_LVT u_T_427_reg_9__30_ ( .D(n4400), .CLK(n4227), .Q(n_T_427[1373]) );
  DFFX1_LVT u_T_427_reg_9__29_ ( .D(n4397), .CLK(n4227), .Q(n_T_427[1372]) );
  DFFX1_LVT u_T_427_reg_9__28_ ( .D(n4394), .CLK(n4227), .Q(n_T_427[1371]) );
  DFFX1_LVT u_T_427_reg_9__27_ ( .D(n4391), .CLK(n4227), .Q(n_T_427[1370]) );
  DFFX1_LVT u_T_427_reg_9__26_ ( .D(n4389), .CLK(n4227), .Q(n_T_427[1369]) );
  DFFX1_LVT u_T_427_reg_9__25_ ( .D(n4387), .CLK(n4227), .Q(n_T_427[1368]) );
  DFFX1_LVT u_T_427_reg_9__24_ ( .D(n4385), .CLK(n4227), .Q(n_T_427[1367]) );
  DFFX1_LVT u_T_427_reg_9__23_ ( .D(n4381), .CLK(n4226), .Q(n_T_427[1366]) );
  DFFX1_LVT u_T_427_reg_9__22_ ( .D(n4379), .CLK(n4226), .Q(n_T_427[1365]) );
  DFFX1_LVT u_T_427_reg_9__21_ ( .D(n4377), .CLK(n4226), .Q(n_T_427[1364]) );
  DFFX1_LVT u_T_427_reg_9__20_ ( .D(n4375), .CLK(n4226), .Q(n_T_427[1363]) );
  DFFX1_LVT u_T_427_reg_9__19_ ( .D(n4372), .CLK(n4226), .Q(n_T_427[1362]) );
  DFFX1_LVT u_T_427_reg_9__18_ ( .D(n4369), .CLK(n4226), .Q(n_T_427[1361]) );
  DFFX1_LVT u_T_427_reg_9__17_ ( .D(n4365), .CLK(n4226), .Q(n_T_427[1360]) );
  DFFX1_LVT u_T_427_reg_9__16_ ( .D(n4362), .CLK(n4226), .Q(n_T_427[1359]) );
  DFFX1_LVT u_T_427_reg_9__15_ ( .D(n4360), .CLK(n4226), .Q(n_T_427[1358]) );
  DFFX1_LVT u_T_427_reg_9__14_ ( .D(n4357), .CLK(n4226), .Q(n_T_427[1357]) );
  DFFX1_LVT u_T_427_reg_9__13_ ( .D(n4355), .CLK(n4226), .Q(n_T_427[1356]) );
  DFFX1_LVT u_T_427_reg_9__12_ ( .D(n4352), .CLK(n4226), .Q(n_T_427[1355]) );
  DFFX1_LVT u_T_427_reg_9__11_ ( .D(n4350), .CLK(n4225), .Q(n_T_427[1354]) );
  DFFX1_LVT u_T_427_reg_9__10_ ( .D(n4346), .CLK(n4225), .Q(n_T_427[1353]) );
  DFFX1_LVT u_T_427_reg_9__9_ ( .D(n4343), .CLK(n4225), .Q(n_T_427[1352]) );
  DFFX1_LVT u_T_427_reg_9__8_ ( .D(n4340), .CLK(n4225), .Q(n_T_427[1351]) );
  DFFX1_LVT u_T_427_reg_9__7_ ( .D(n4337), .CLK(n4225), .Q(n_T_427[1350]) );
  DFFX1_LVT u_T_427_reg_9__6_ ( .D(n4334), .CLK(n4225), .Q(n_T_427[1349]) );
  DFFX1_LVT u_T_427_reg_9__5_ ( .D(n4331), .CLK(n4225), .Q(n_T_427[1348]) );
  DFFX1_LVT u_T_427_reg_9__4_ ( .D(n4328), .CLK(n4225), .Q(n_T_427[1347]) );
  DFFX1_LVT u_T_427_reg_9__3_ ( .D(n4325), .CLK(n4225), .Q(n_T_427[1346]) );
  DFFX1_LVT u_T_427_reg_9__2_ ( .D(n4322), .CLK(n4225), .Q(n_T_427[1345]) );
  DFFX1_LVT u_T_427_reg_9__1_ ( .D(n4320), .CLK(n4225), .Q(n_T_427[1344]) );
  DFFX1_LVT u_T_427_reg_9__0_ ( .D(n4317), .CLK(n4225), .Q(n_T_427[1343]) );
  DFFX1_LVT u_T_427_reg_10__63_ ( .D(n4494), .CLK(n4224), .Q(n_T_427[1342]) );
  DFFX1_LVT u_T_427_reg_10__62_ ( .D(n4491), .CLK(n4224), .Q(n_T_427[1341]) );
  DFFX1_LVT u_T_427_reg_10__61_ ( .D(n4488), .CLK(n4224), .Q(n_T_427[1340]) );
  DFFX1_LVT u_T_427_reg_10__60_ ( .D(n4485), .CLK(n4224), .Q(n_T_427[1339]) );
  DFFX1_LVT u_T_427_reg_10__59_ ( .D(n4482), .CLK(n4223), .Q(n_T_427[1338]) );
  DFFX1_LVT u_T_427_reg_10__58_ ( .D(n4480), .CLK(n4223), .Q(n_T_427[1337]) );
  DFFX1_LVT u_T_427_reg_10__57_ ( .D(n4476), .CLK(n4223), .Q(n_T_427[1336]) );
  DFFX1_LVT u_T_427_reg_10__56_ ( .D(n4474), .CLK(n4223), .Q(n_T_427[1335]) );
  DFFX1_LVT u_T_427_reg_10__55_ ( .D(n4470), .CLK(n4223), .Q(n_T_427[1334]) );
  DFFX1_LVT u_T_427_reg_10__54_ ( .D(n4468), .CLK(n4223), .Q(n_T_427[1333]) );
  DFFX1_LVT u_T_427_reg_10__53_ ( .D(n4464), .CLK(n4223), .Q(n_T_427[1332]) );
  DFFX1_LVT u_T_427_reg_10__52_ ( .D(n4462), .CLK(n4223), .Q(n_T_427[1331]) );
  DFFX1_LVT u_T_427_reg_10__51_ ( .D(n4459), .CLK(n4223), .Q(n_T_427[1330]) );
  DFFX1_LVT u_T_427_reg_10__50_ ( .D(n4455), .CLK(n4223), .Q(n_T_427[1329]) );
  DFFX1_LVT u_T_427_reg_10__49_ ( .D(n4453), .CLK(n4223), .Q(n_T_427[1328]) );
  DFFX1_LVT u_T_427_reg_10__48_ ( .D(n4449), .CLK(n4223), .Q(n_T_427[1327]) );
  DFFX1_LVT u_T_427_reg_10__47_ ( .D(n4446), .CLK(n4222), .Q(n_T_427[1326]) );
  DFFX1_LVT u_T_427_reg_10__46_ ( .D(n4443), .CLK(n4222), .Q(n_T_427[1325]) );
  DFFX1_LVT u_T_427_reg_10__45_ ( .D(n4441), .CLK(n4222), .Q(n_T_427[1324]) );
  DFFX1_LVT u_T_427_reg_10__44_ ( .D(n4437), .CLK(n4222), .Q(n_T_427[1323]) );
  DFFX1_LVT u_T_427_reg_10__43_ ( .D(n4435), .CLK(n4222), .Q(n_T_427[1322]) );
  DFFX1_LVT u_T_427_reg_10__42_ ( .D(n4432), .CLK(n4222), .Q(n_T_427[1321]) );
  DFFX1_LVT u_T_427_reg_10__41_ ( .D(n4429), .CLK(n4222), .Q(n_T_427[1320]) );
  DFFX1_LVT u_T_427_reg_10__40_ ( .D(n4425), .CLK(n4222), .Q(n_T_427[1319]) );
  DFFX1_LVT u_T_427_reg_10__39_ ( .D(n4422), .CLK(n4222), .Q(n_T_427[1318]) );
  DFFX1_LVT u_T_427_reg_10__38_ ( .D(n4420), .CLK(n4222), .Q(n_T_427[1317]) );
  DFFX1_LVT u_T_427_reg_10__37_ ( .D(n4417), .CLK(n4222), .Q(n_T_427[1316]) );
  DFFX1_LVT u_T_427_reg_10__36_ ( .D(n4415), .CLK(n4222), .Q(n_T_427[1315]) );
  DFFX1_LVT u_T_427_reg_10__35_ ( .D(n4412), .CLK(n4221), .Q(n_T_427[1314]) );
  DFFX1_LVT u_T_427_reg_10__34_ ( .D(n4409), .CLK(n4221), .Q(n_T_427[1313]) );
  DFFX1_LVT u_T_427_reg_10__33_ ( .D(n4407), .CLK(n4221), .Q(n_T_427[1312]) );
  DFFX1_LVT u_T_427_reg_10__32_ ( .D(n4404), .CLK(n4221), .Q(n_T_427[1311]) );
  DFFX1_LVT u_T_427_reg_10__31_ ( .D(n4402), .CLK(n4221), .Q(n_T_427[1310]) );
  DFFX1_LVT u_T_427_reg_10__30_ ( .D(n4400), .CLK(n4221), .Q(n_T_427[1309]) );
  DFFX1_LVT u_T_427_reg_10__29_ ( .D(n4397), .CLK(n4221), .Q(n_T_427[1308]) );
  DFFX1_LVT u_T_427_reg_10__28_ ( .D(n4394), .CLK(n4221), .Q(n_T_427[1307]) );
  DFFX1_LVT u_T_427_reg_10__27_ ( .D(n4391), .CLK(n4221), .Q(n_T_427[1306]) );
  DFFX1_LVT u_T_427_reg_10__26_ ( .D(n4389), .CLK(n4221), .Q(n_T_427[1305]) );
  DFFX1_LVT u_T_427_reg_10__25_ ( .D(n4387), .CLK(n4221), .Q(n_T_427[1304]) );
  DFFX1_LVT u_T_427_reg_10__24_ ( .D(n4385), .CLK(n4221), .Q(n_T_427[1303]) );
  DFFX1_LVT u_T_427_reg_10__23_ ( .D(n4381), .CLK(n4220), .Q(n_T_427[1302]) );
  DFFX1_LVT u_T_427_reg_10__22_ ( .D(n4379), .CLK(n4220), .Q(n_T_427[1301]) );
  DFFX1_LVT u_T_427_reg_10__21_ ( .D(n4377), .CLK(n4220), .Q(n_T_427[1300]) );
  DFFX1_LVT u_T_427_reg_10__20_ ( .D(n4375), .CLK(n4220), .Q(n_T_427[1299]) );
  DFFX1_LVT u_T_427_reg_10__19_ ( .D(n4372), .CLK(n4220), .Q(n_T_427[1298]) );
  DFFX1_LVT u_T_427_reg_10__18_ ( .D(n4369), .CLK(n4220), .Q(n_T_427[1297]) );
  DFFX1_LVT u_T_427_reg_10__17_ ( .D(n4365), .CLK(n4220), .Q(n_T_427[1296]) );
  DFFX1_LVT u_T_427_reg_10__16_ ( .D(n4362), .CLK(n4220), .Q(n_T_427[1295]) );
  DFFX1_LVT u_T_427_reg_10__15_ ( .D(n4360), .CLK(n4220), .Q(n_T_427[1294]) );
  DFFX1_LVT u_T_427_reg_10__14_ ( .D(n4357), .CLK(n4220), .Q(n_T_427[1293]) );
  DFFX1_LVT u_T_427_reg_10__13_ ( .D(n4355), .CLK(n4220), .Q(n_T_427[1292]) );
  DFFX1_LVT u_T_427_reg_10__12_ ( .D(n4352), .CLK(n4220), .Q(n_T_427[1291]) );
  DFFX1_LVT u_T_427_reg_10__11_ ( .D(n4350), .CLK(n4219), .Q(n_T_427[1290]) );
  DFFX1_LVT u_T_427_reg_10__10_ ( .D(n4346), .CLK(n4219), .Q(n_T_427[1289]) );
  DFFX1_LVT u_T_427_reg_10__9_ ( .D(n4343), .CLK(n4219), .Q(n_T_427[1288]) );
  DFFX1_LVT u_T_427_reg_10__8_ ( .D(n4340), .CLK(n4219), .Q(n_T_427[1287]) );
  DFFX1_LVT u_T_427_reg_10__7_ ( .D(n4337), .CLK(n4219), .Q(n_T_427[1286]) );
  DFFX1_LVT u_T_427_reg_10__6_ ( .D(n4334), .CLK(n4219), .Q(n_T_427[1285]) );
  DFFX1_LVT u_T_427_reg_10__5_ ( .D(n4331), .CLK(n4219), .Q(n_T_427[1284]) );
  DFFX1_LVT u_T_427_reg_10__4_ ( .D(n4328), .CLK(n4219), .Q(n_T_427[1283]) );
  DFFX1_LVT u_T_427_reg_10__3_ ( .D(n4325), .CLK(n4219), .Q(n_T_427[1282]) );
  DFFX1_LVT u_T_427_reg_10__2_ ( .D(n4322), .CLK(n4219), .Q(n_T_427[1281]) );
  DFFX1_LVT u_T_427_reg_10__1_ ( .D(n4320), .CLK(n4219), .Q(n_T_427[1280]) );
  DFFX1_LVT u_T_427_reg_10__0_ ( .D(n4317), .CLK(n4219), .Q(n_T_427[1279]) );
  DFFX1_LVT u_T_427_reg_11__63_ ( .D(n4494), .CLK(n4218), .Q(n_T_427[1278]) );
  DFFX1_LVT u_T_427_reg_11__62_ ( .D(n4491), .CLK(n4218), .Q(n_T_427[1277]) );
  DFFX1_LVT u_T_427_reg_11__61_ ( .D(n4488), .CLK(n4218), .Q(n_T_427[1276]) );
  DFFX1_LVT u_T_427_reg_11__60_ ( .D(n4485), .CLK(n4218), .Q(n_T_427[1275]) );
  DFFX1_LVT u_T_427_reg_11__59_ ( .D(n4482), .CLK(n4217), .Q(n_T_427[1274]) );
  DFFX1_LVT u_T_427_reg_11__58_ ( .D(n4480), .CLK(n4217), .Q(n_T_427[1273]) );
  DFFX1_LVT u_T_427_reg_11__57_ ( .D(n4476), .CLK(n4217), .Q(n_T_427[1272]) );
  DFFX1_LVT u_T_427_reg_11__56_ ( .D(n4474), .CLK(n4217), .Q(n_T_427[1271]) );
  DFFX1_LVT u_T_427_reg_11__55_ ( .D(n4470), .CLK(n4217), .Q(n_T_427[1270]) );
  DFFX1_LVT u_T_427_reg_11__54_ ( .D(n4468), .CLK(n4217), .Q(n_T_427[1269]) );
  DFFX1_LVT u_T_427_reg_11__53_ ( .D(n4464), .CLK(n4217), .Q(n_T_427[1268]) );
  DFFX1_LVT u_T_427_reg_11__52_ ( .D(n4462), .CLK(n4217), .Q(n_T_427[1267]) );
  DFFX1_LVT u_T_427_reg_11__51_ ( .D(n4459), .CLK(n4217), .Q(n_T_427[1266]) );
  DFFX1_LVT u_T_427_reg_11__50_ ( .D(n4455), .CLK(n4217), .Q(n_T_427[1265]) );
  DFFX1_LVT u_T_427_reg_11__49_ ( .D(n4453), .CLK(n4217), .Q(n_T_427[1264]) );
  DFFX1_LVT u_T_427_reg_11__48_ ( .D(n4449), .CLK(n4217), .Q(n_T_427[1263]) );
  DFFX1_LVT u_T_427_reg_11__47_ ( .D(n4446), .CLK(n4216), .Q(n_T_427[1262]) );
  DFFX1_LVT u_T_427_reg_11__46_ ( .D(n4443), .CLK(n4216), .Q(n_T_427[1261]) );
  DFFX1_LVT u_T_427_reg_11__45_ ( .D(n4441), .CLK(n4216), .Q(n_T_427[1260]) );
  DFFX1_LVT u_T_427_reg_11__44_ ( .D(n4437), .CLK(n4216), .Q(n_T_427[1259]) );
  DFFX1_LVT u_T_427_reg_11__43_ ( .D(n4435), .CLK(n4216), .Q(n_T_427[1258]) );
  DFFX1_LVT u_T_427_reg_11__42_ ( .D(n4432), .CLK(n4216), .Q(n_T_427[1257]) );
  DFFX1_LVT u_T_427_reg_11__41_ ( .D(n4429), .CLK(n4216), .Q(n_T_427[1256]) );
  DFFX1_LVT u_T_427_reg_11__40_ ( .D(n4425), .CLK(n4216), .Q(n_T_427[1255]) );
  DFFX1_LVT u_T_427_reg_11__39_ ( .D(n4422), .CLK(n4216), .Q(n_T_427[1254]) );
  DFFX1_LVT u_T_427_reg_11__38_ ( .D(n4420), .CLK(n4216), .Q(n_T_427[1253]) );
  DFFX1_LVT u_T_427_reg_11__37_ ( .D(n4417), .CLK(n4216), .Q(n_T_427[1252]) );
  DFFX1_LVT u_T_427_reg_11__36_ ( .D(n4415), .CLK(n4216), .Q(n_T_427[1251]) );
  DFFX1_LVT u_T_427_reg_11__35_ ( .D(n4412), .CLK(n4215), .Q(n_T_427[1250]) );
  DFFX1_LVT u_T_427_reg_11__34_ ( .D(n4409), .CLK(n4215), .Q(n_T_427[1249]) );
  DFFX1_LVT u_T_427_reg_11__33_ ( .D(n4407), .CLK(n4215), .Q(n_T_427[1248]) );
  DFFX1_LVT u_T_427_reg_11__32_ ( .D(n4404), .CLK(n4215), .Q(n_T_427[1247]) );
  DFFX1_LVT u_T_427_reg_11__31_ ( .D(n4402), .CLK(n4215), .Q(n_T_427[1246]) );
  DFFX1_LVT u_T_427_reg_11__30_ ( .D(n4400), .CLK(n4215), .Q(n_T_427[1245]) );
  DFFX1_LVT u_T_427_reg_11__29_ ( .D(n4397), .CLK(n4215), .Q(n_T_427[1244]) );
  DFFX1_LVT u_T_427_reg_11__28_ ( .D(n4394), .CLK(n4215), .Q(n_T_427[1243]) );
  DFFX1_LVT u_T_427_reg_11__27_ ( .D(n4391), .CLK(n4215), .Q(n_T_427[1242]) );
  DFFX1_LVT u_T_427_reg_11__26_ ( .D(n4389), .CLK(n4215), .Q(n_T_427[1241]) );
  DFFX1_LVT u_T_427_reg_11__25_ ( .D(n4387), .CLK(n4215), .Q(n_T_427[1240]) );
  DFFX1_LVT u_T_427_reg_11__24_ ( .D(n4385), .CLK(n4215), .Q(n_T_427[1239]) );
  DFFX1_LVT u_T_427_reg_11__23_ ( .D(n4381), .CLK(n4214), .Q(n_T_427[1238]) );
  DFFX1_LVT u_T_427_reg_11__22_ ( .D(n4379), .CLK(n4214), .Q(n_T_427[1237]) );
  DFFX1_LVT u_T_427_reg_11__21_ ( .D(n4377), .CLK(n4214), .Q(n_T_427[1236]) );
  DFFX1_LVT u_T_427_reg_11__20_ ( .D(n4375), .CLK(n4214), .Q(n_T_427[1235]) );
  DFFX1_LVT u_T_427_reg_11__19_ ( .D(n4372), .CLK(n4214), .Q(n_T_427[1234]) );
  DFFX1_LVT u_T_427_reg_11__18_ ( .D(n4369), .CLK(n4214), .Q(n_T_427[1233]) );
  DFFX1_LVT u_T_427_reg_11__17_ ( .D(n4365), .CLK(n4214), .Q(n_T_427[1232]) );
  DFFX1_LVT u_T_427_reg_11__16_ ( .D(n4362), .CLK(n4214), .Q(n_T_427[1231]) );
  DFFX1_LVT u_T_427_reg_11__15_ ( .D(n4360), .CLK(n4214), .Q(n_T_427[1230]) );
  DFFX1_LVT u_T_427_reg_11__14_ ( .D(n4357), .CLK(n4214), .Q(n_T_427[1229]) );
  DFFX1_LVT u_T_427_reg_11__13_ ( .D(n4355), .CLK(n4214), .Q(n_T_427[1228]) );
  DFFX1_LVT u_T_427_reg_11__12_ ( .D(n4352), .CLK(n4214), .Q(n_T_427[1227]) );
  DFFX1_LVT u_T_427_reg_11__11_ ( .D(n4350), .CLK(n4213), .Q(n_T_427[1226]) );
  DFFX1_LVT u_T_427_reg_11__10_ ( .D(n4346), .CLK(n4213), .Q(n_T_427[1225]) );
  DFFX1_LVT u_T_427_reg_11__9_ ( .D(n4343), .CLK(n4213), .Q(n_T_427[1224]) );
  DFFX1_LVT u_T_427_reg_11__8_ ( .D(n4340), .CLK(n4213), .Q(n_T_427[1223]) );
  DFFX1_LVT u_T_427_reg_11__7_ ( .D(n4337), .CLK(n4213), .Q(n_T_427[1222]) );
  DFFX1_LVT u_T_427_reg_11__6_ ( .D(n4334), .CLK(n4213), .Q(n_T_427[1221]) );
  DFFX1_LVT u_T_427_reg_11__5_ ( .D(n4331), .CLK(n4213), .Q(n_T_427[1220]) );
  DFFX1_LVT u_T_427_reg_11__4_ ( .D(n4328), .CLK(n4213), .Q(n_T_427[1219]) );
  DFFX1_LVT u_T_427_reg_11__3_ ( .D(n4325), .CLK(n4213), .Q(n_T_427[1218]) );
  DFFX1_LVT u_T_427_reg_11__2_ ( .D(n4322), .CLK(n4213), .Q(n_T_427[1217]) );
  DFFX1_LVT u_T_427_reg_11__1_ ( .D(n4320), .CLK(n4213), .Q(n_T_427[1216]) );
  DFFX1_LVT u_T_427_reg_11__0_ ( .D(n4317), .CLK(n4213), .Q(n_T_427[1215]) );
  DFFX1_LVT u_T_427_reg_12__63_ ( .D(n4495), .CLK(n4212), .Q(n_T_427[1214]), 
        .QN(n3308) );
  DFFX1_LVT u_T_427_reg_12__62_ ( .D(n4492), .CLK(n4212), .Q(n_T_427[1213]), 
        .QN(n3306) );
  DFFX1_LVT u_T_427_reg_12__61_ ( .D(n4489), .CLK(n4212), .Q(n_T_427[1212]), 
        .QN(n3305) );
  DFFX1_LVT u_T_427_reg_12__60_ ( .D(n4486), .CLK(n4212), .Q(n_T_427[1211]), 
        .QN(n3304) );
  DFFX1_LVT u_T_427_reg_12__58_ ( .D(n4480), .CLK(n4211), .Q(n_T_427[1209]), 
        .QN(n3365) );
  DFFX1_LVT u_T_427_reg_12__56_ ( .D(n4474), .CLK(n4211), .Q(n_T_427[1207]), 
        .QN(n3362) );
  DFFX1_LVT u_T_427_reg_12__54_ ( .D(n4468), .CLK(n4211), .Q(n_T_427[1205]), 
        .QN(n3360) );
  DFFX1_LVT u_T_427_reg_12__52_ ( .D(n4462), .CLK(n4211), .Q(n_T_427[1203]), 
        .QN(n3355) );
  DFFX1_LVT u_T_427_reg_12__51_ ( .D(n4459), .CLK(n4211), .Q(n_T_427[1202]), 
        .QN(n3354) );
  DFFX1_LVT u_T_427_reg_12__49_ ( .D(n4453), .CLK(n4211), .Q(n_T_427[1200]), 
        .QN(n3349) );
  DFFX1_LVT u_T_427_reg_12__45_ ( .D(n4441), .CLK(n4210), .Q(n_T_427[1196]), 
        .QN(n3343) );
  DFFX1_LVT u_T_427_reg_12__43_ ( .D(n4435), .CLK(n4210), .Q(n_T_427[1194]), 
        .QN(n3340) );
  DFFX1_LVT u_T_427_reg_12__42_ ( .D(n4432), .CLK(n4210), .Q(n_T_427[1193]) );
  DFFX1_LVT u_T_427_reg_12__41_ ( .D(n4429), .CLK(n4210), .Q(n_T_427[1192]), 
        .QN(n3339) );
  DFFX1_LVT u_T_427_reg_12__39_ ( .D(n4423), .CLK(n4210), .Q(n_T_427[1190]) );
  DFFX1_LVT u_T_427_reg_12__38_ ( .D(n4420), .CLK(n4210), .Q(n_T_427[1189]) );
  DFFX1_LVT u_T_427_reg_12__36_ ( .D(n4415), .CLK(n4210), .Q(n_T_427[1187]) );
  DFFX1_LVT u_T_427_reg_12__30_ ( .D(n4400), .CLK(n4209), .Q(n_T_427[1181]), 
        .QN(n3331) );
  DFFX1_LVT u_T_427_reg_12__29_ ( .D(n4397), .CLK(n4209), .Q(n_T_427[1180]), 
        .QN(n3294) );
  DFFX1_LVT u_T_427_reg_12__27_ ( .D(n4392), .CLK(n4209), .Q(n_T_427[1178]), 
        .QN(n3328) );
  DFFX1_LVT u_T_427_reg_12__24_ ( .D(n4385), .CLK(n4209), .Q(n_T_427[1175]), 
        .QN(n3326) );
  DFFX1_LVT u_T_427_reg_12__20_ ( .D(n4375), .CLK(n4208), .Q(n_T_427[1171]), 
        .QN(n3320) );
  DFFX1_LVT u_T_427_reg_12__19_ ( .D(n4372), .CLK(n4208), .Q(n_T_427[1170]), 
        .QN(n3317) );
  DFFX1_LVT u_T_427_reg_12__18_ ( .D(n4369), .CLK(n4208), .Q(n_T_427[1169]), 
        .QN(n3314) );
  DFFX1_LVT u_T_427_reg_12__1_ ( .D(n4320), .CLK(n4207), .Q(n_T_427[1152]) );
  DFFX1_LVT u_T_427_reg_12__0_ ( .D(n4317), .CLK(n4207), .Q(n_T_427[1151]) );
  DFFX1_LVT u_T_427_reg_13__63_ ( .D(n4495), .CLK(n4206), .Q(n_T_427[1150]) );
  DFFX1_LVT u_T_427_reg_13__62_ ( .D(n4492), .CLK(n4206), .Q(n_T_427[1149]) );
  DFFX1_LVT u_T_427_reg_13__61_ ( .D(n4489), .CLK(n4206), .Q(n_T_427[1148]) );
  DFFX1_LVT u_T_427_reg_13__60_ ( .D(n4486), .CLK(n4206), .Q(n_T_427[1147]) );
  DFFX1_LVT u_T_427_reg_13__59_ ( .D(n4483), .CLK(n4205), .Q(n_T_427[1146]) );
  DFFX1_LVT u_T_427_reg_13__58_ ( .D(n4480), .CLK(n4205), .Q(n_T_427[1145]) );
  DFFX1_LVT u_T_427_reg_13__57_ ( .D(n4477), .CLK(n4205), .Q(n_T_427[1144]) );
  DFFX1_LVT u_T_427_reg_13__56_ ( .D(n4474), .CLK(n4205), .Q(n_T_427[1143]) );
  DFFX1_LVT u_T_427_reg_13__55_ ( .D(n4471), .CLK(n4205), .Q(n_T_427[1142]) );
  DFFX1_LVT u_T_427_reg_13__54_ ( .D(n4468), .CLK(n4205), .Q(n_T_427[1141]) );
  DFFX1_LVT u_T_427_reg_13__53_ ( .D(n4465), .CLK(n4205), .Q(n_T_427[1140]) );
  DFFX1_LVT u_T_427_reg_13__52_ ( .D(n4462), .CLK(n4205), .Q(n_T_427[1139]) );
  DFFX1_LVT u_T_427_reg_13__51_ ( .D(n4459), .CLK(n4205), .Q(n_T_427[1138]) );
  DFFX1_LVT u_T_427_reg_13__50_ ( .D(n4456), .CLK(n4205), .Q(n_T_427[1137]) );
  DFFX1_LVT u_T_427_reg_13__49_ ( .D(n4453), .CLK(n4205), .Q(n_T_427[1136]) );
  DFFX1_LVT u_T_427_reg_13__48_ ( .D(n4450), .CLK(n4205), .Q(n_T_427[1135]) );
  DFFX1_LVT u_T_427_reg_13__47_ ( .D(n4447), .CLK(n4204), .Q(n_T_427[1134]) );
  DFFX1_LVT u_T_427_reg_13__46_ ( .D(n4444), .CLK(n4204), .Q(n_T_427[1133]) );
  DFFX1_LVT u_T_427_reg_13__45_ ( .D(n4441), .CLK(n4204), .Q(n_T_427[1132]) );
  DFFX1_LVT u_T_427_reg_13__44_ ( .D(n4438), .CLK(n4204), .Q(n_T_427[1131]) );
  DFFX1_LVT u_T_427_reg_13__43_ ( .D(n4435), .CLK(n4204), .Q(n_T_427[1130]) );
  DFFX1_LVT u_T_427_reg_13__42_ ( .D(n4432), .CLK(n4204), .Q(n_T_427[1129]) );
  DFFX1_LVT u_T_427_reg_13__41_ ( .D(n4429), .CLK(n4204), .Q(n_T_427[1128]) );
  DFFX1_LVT u_T_427_reg_13__40_ ( .D(n4426), .CLK(n4204), .Q(n_T_427[1127]) );
  DFFX1_LVT u_T_427_reg_13__39_ ( .D(n4423), .CLK(n4204), .Q(n_T_427[1126]) );
  DFFX1_LVT u_T_427_reg_13__38_ ( .D(n4420), .CLK(n4204), .Q(n_T_427[1125]) );
  DFFX1_LVT u_T_427_reg_13__37_ ( .D(n4418), .CLK(n4204), .Q(n_T_427[1124]) );
  DFFX1_LVT u_T_427_reg_13__36_ ( .D(n4415), .CLK(n4204), .Q(n_T_427[1123]) );
  DFFX1_LVT u_T_427_reg_13__35_ ( .D(n4412), .CLK(n4203), .Q(n_T_427[1122]) );
  DFFX1_LVT u_T_427_reg_13__34_ ( .D(n4410), .CLK(n4203), .Q(n_T_427[1121]) );
  DFFX1_LVT u_T_427_reg_13__33_ ( .D(n4407), .CLK(n4203), .Q(n_T_427[1120]) );
  DFFX1_LVT u_T_427_reg_13__32_ ( .D(n4405), .CLK(n4203), .Q(n_T_427[1119]) );
  DFFX1_LVT u_T_427_reg_13__31_ ( .D(n4402), .CLK(n4203), .Q(n_T_427[1118]) );
  DFFX1_LVT u_T_427_reg_13__30_ ( .D(n4400), .CLK(n4203), .Q(n_T_427[1117]) );
  DFFX1_LVT u_T_427_reg_13__29_ ( .D(n4397), .CLK(n4203), .Q(n_T_427[1116]) );
  DFFX1_LVT u_T_427_reg_13__28_ ( .D(n4394), .CLK(n4203), .Q(n_T_427[1115]) );
  DFFX1_LVT u_T_427_reg_13__27_ ( .D(n4392), .CLK(n4203), .Q(n_T_427[1114]) );
  DFFX1_LVT u_T_427_reg_13__26_ ( .D(n4389), .CLK(n4203), .Q(n_T_427[1113]) );
  DFFX1_LVT u_T_427_reg_13__25_ ( .D(n4387), .CLK(n4203), .Q(n_T_427[1112]) );
  DFFX1_LVT u_T_427_reg_13__24_ ( .D(n4385), .CLK(n4203), .Q(n_T_427[1111]) );
  DFFX1_LVT u_T_427_reg_13__23_ ( .D(n4382), .CLK(n4202), .Q(n_T_427[1110]) );
  DFFX1_LVT u_T_427_reg_13__22_ ( .D(n4379), .CLK(n4202), .Q(n_T_427[1109]) );
  DFFX1_LVT u_T_427_reg_13__21_ ( .D(n4377), .CLK(n4202), .Q(n_T_427[1108]) );
  DFFX1_LVT u_T_427_reg_13__20_ ( .D(n4375), .CLK(n4202), .Q(n_T_427[1107]) );
  DFFX1_LVT u_T_427_reg_13__19_ ( .D(n4372), .CLK(n4202), .Q(n_T_427[1106]) );
  DFFX1_LVT u_T_427_reg_13__18_ ( .D(n4369), .CLK(n4202), .Q(n_T_427[1105]) );
  DFFX1_LVT u_T_427_reg_13__17_ ( .D(n4366), .CLK(n4202), .Q(n_T_427[1104]) );
  DFFX1_LVT u_T_427_reg_13__16_ ( .D(n4363), .CLK(n4202), .Q(n_T_427[1103]) );
  DFFX1_LVT u_T_427_reg_13__15_ ( .D(n4360), .CLK(n4202), .Q(n_T_427[1102]) );
  DFFX1_LVT u_T_427_reg_13__14_ ( .D(n4358), .CLK(n4202), .Q(n_T_427[1101]) );
  DFFX1_LVT u_T_427_reg_13__13_ ( .D(n4355), .CLK(n4202), .Q(n_T_427[1100]) );
  DFFX1_LVT u_T_427_reg_13__12_ ( .D(n4353), .CLK(n4202), .Q(n_T_427[1099]) );
  DFFX1_LVT u_T_427_reg_13__11_ ( .D(n4350), .CLK(n4201), .Q(n_T_427[1098]) );
  DFFX1_LVT u_T_427_reg_13__10_ ( .D(n4347), .CLK(n4201), .Q(n_T_427[1097]) );
  DFFX1_LVT u_T_427_reg_13__9_ ( .D(n4344), .CLK(n4201), .Q(n_T_427[1096]) );
  DFFX1_LVT u_T_427_reg_13__8_ ( .D(n4341), .CLK(n4201), .Q(n_T_427[1095]) );
  DFFX1_LVT u_T_427_reg_13__7_ ( .D(n4338), .CLK(n4201), .Q(n_T_427[1094]) );
  DFFX1_LVT u_T_427_reg_13__6_ ( .D(n4335), .CLK(n4201), .Q(n_T_427[1093]) );
  DFFX1_LVT u_T_427_reg_13__5_ ( .D(n4332), .CLK(n4201), .Q(n_T_427[1092]) );
  DFFX1_LVT u_T_427_reg_13__4_ ( .D(n4329), .CLK(n4201), .Q(n_T_427[1091]) );
  DFFX1_LVT u_T_427_reg_13__3_ ( .D(n4326), .CLK(n4201), .Q(n_T_427[1090]) );
  DFFX1_LVT u_T_427_reg_13__2_ ( .D(n4323), .CLK(n4201), .Q(n_T_427[1089]) );
  DFFX1_LVT u_T_427_reg_13__1_ ( .D(n4320), .CLK(n4201), .Q(n_T_427[1088]) );
  DFFX1_LVT u_T_427_reg_13__0_ ( .D(n4317), .CLK(n4201), .Q(n_T_427[1087]) );
  DFFX1_LVT u_T_427_reg_14__63_ ( .D(n4495), .CLK(n4200), .Q(n_T_427[1086]), 
        .QN(n3309) );
  DFFX1_LVT u_T_427_reg_14__62_ ( .D(n4492), .CLK(n4200), .Q(n_T_427[1085]), 
        .QN(n3307) );
  DFFX1_LVT u_T_427_reg_14__61_ ( .D(n4489), .CLK(n4200), .Q(n_T_427[1084]), 
        .QN(n3281) );
  DFFX1_LVT u_T_427_reg_14__60_ ( .D(n4486), .CLK(n4200), .Q(n_T_427[1083]), 
        .QN(n3303) );
  DFFX1_LVT u_T_427_reg_14__58_ ( .D(n4480), .CLK(n4199), .Q(n_T_427[1081]), 
        .QN(n3366) );
  DFFX1_LVT u_T_427_reg_14__56_ ( .D(n4474), .CLK(n4199), .Q(n_T_427[1079]) );
  DFFX1_LVT u_T_427_reg_14__55_ ( .D(n4471), .CLK(n4199), .Q(n_T_427[1078]) );
  DFFX1_LVT u_T_427_reg_14__54_ ( .D(n4468), .CLK(n4199), .Q(n_T_427[1077]), 
        .QN(n3359) );
  DFFX1_LVT u_T_427_reg_14__52_ ( .D(n4462), .CLK(n4199), .Q(n_T_427[1075]), 
        .QN(n3356) );
  DFFX1_LVT u_T_427_reg_14__51_ ( .D(n4459), .CLK(n4199), .Q(n_T_427[1074]), 
        .QN(n3353) );
  DFFX1_LVT u_T_427_reg_14__49_ ( .D(n4453), .CLK(n4199), .Q(n_T_427[1072]), 
        .QN(n3350) );
  DFFX1_LVT u_T_427_reg_14__48_ ( .D(n4450), .CLK(n4199), .Q(n_T_427[1071]) );
  DFFX1_LVT u_T_427_reg_14__45_ ( .D(n4441), .CLK(n4198), .Q(n_T_427[1068]), 
        .QN(n3344) );
  DFFX1_LVT u_T_427_reg_14__44_ ( .D(n4438), .CLK(n4198), .Q(n_T_427[1067]) );
  DFFX1_LVT u_T_427_reg_14__43_ ( .D(n4435), .CLK(n4198), .Q(n_T_427[1066]), 
        .QN(n3341) );
  DFFX1_LVT u_T_427_reg_14__42_ ( .D(n4432), .CLK(n4198), .Q(n_T_427[1065]) );
  DFFX1_LVT u_T_427_reg_14__41_ ( .D(n4429), .CLK(n4198), .Q(n_T_427[1064]) );
  DFFX1_LVT u_T_427_reg_14__39_ ( .D(n4423), .CLK(n4198), .Q(n_T_427[1062]) );
  DFFX1_LVT u_T_427_reg_14__38_ ( .D(n4420), .CLK(n4198), .Q(n_T_427[1061]) );
  DFFX1_LVT u_T_427_reg_14__37_ ( .D(n4418), .CLK(n4198), .Q(n_T_427[1060]) );
  DFFX1_LVT u_T_427_reg_14__36_ ( .D(n4415), .CLK(n4198), .Q(n_T_427[1059]) );
  DFFX1_LVT u_T_427_reg_14__35_ ( .D(n4412), .CLK(n4197), .Q(n_T_427[1058]) );
  DFFX1_LVT u_T_427_reg_14__34_ ( .D(n4410), .CLK(n4197), .Q(n_T_427[1057]) );
  DFFX1_LVT u_T_427_reg_14__33_ ( .D(n4407), .CLK(n4197), .Q(n_T_427[1056]) );
  DFFX1_LVT u_T_427_reg_14__30_ ( .D(n4400), .CLK(n4197), .Q(n_T_427[1053]), 
        .QN(n3332) );
  DFFX1_LVT u_T_427_reg_14__29_ ( .D(n4397), .CLK(n4197), .Q(n_T_427[1052]), 
        .QN(n3295) );
  DFFX1_LVT u_T_427_reg_14__27_ ( .D(n4392), .CLK(n4197), .Q(n_T_427[1050]), 
        .QN(n3329) );
  DFFX1_LVT u_T_427_reg_14__24_ ( .D(n4385), .CLK(n4197), .Q(n_T_427[1047]), 
        .QN(n3327) );
  DFFX1_LVT u_T_427_reg_14__20_ ( .D(n4375), .CLK(n4196), .Q(n_T_427[1043]), 
        .QN(n3321) );
  DFFX1_LVT u_T_427_reg_14__19_ ( .D(n4372), .CLK(n4196), .Q(n_T_427[1042]), 
        .QN(n3318) );
  DFFX1_LVT u_T_427_reg_14__18_ ( .D(n4369), .CLK(n4196), .Q(n_T_427[1041]), 
        .QN(n3315) );
  DFFX1_LVT u_T_427_reg_14__15_ ( .D(n4360), .CLK(n4196), .Q(n_T_427[1038]) );
  DFFX1_LVT u_T_427_reg_14__14_ ( .D(n4358), .CLK(n4196), .Q(n_T_427[1037]) );
  DFFX1_LVT u_T_427_reg_14__13_ ( .D(n4355), .CLK(n4196), .Q(n_T_427[1036]) );
  DFFX1_LVT u_T_427_reg_14__12_ ( .D(n4353), .CLK(n4196), .Q(n_T_427[1035]) );
  DFFX1_LVT u_T_427_reg_14__11_ ( .D(n4350), .CLK(n4195), .Q(n_T_427[1034]) );
  DFFX1_LVT u_T_427_reg_14__10_ ( .D(n4347), .CLK(n4195), .Q(n_T_427[1033]) );
  DFFX1_LVT u_T_427_reg_14__9_ ( .D(n4344), .CLK(n4195), .Q(n_T_427[1032]) );
  DFFX1_LVT u_T_427_reg_14__8_ ( .D(n4341), .CLK(n4195), .Q(n_T_427[1031]) );
  DFFX1_LVT u_T_427_reg_14__7_ ( .D(n4338), .CLK(n4195), .Q(n_T_427[1030]) );
  DFFX1_LVT u_T_427_reg_14__6_ ( .D(n4335), .CLK(n4195), .Q(n_T_427[1029]) );
  DFFX1_LVT u_T_427_reg_14__5_ ( .D(n4332), .CLK(n4195), .Q(n_T_427[1028]) );
  DFFX1_LVT u_T_427_reg_14__4_ ( .D(n4329), .CLK(n4195), .Q(n_T_427[1027]) );
  DFFX1_LVT u_T_427_reg_14__3_ ( .D(n4326), .CLK(n4195), .Q(n_T_427[1026]) );
  DFFX1_LVT u_T_427_reg_14__2_ ( .D(n4323), .CLK(n4195), .Q(n_T_427[1025]) );
  DFFX1_LVT u_T_427_reg_14__1_ ( .D(n4320), .CLK(n4195), .Q(n_T_427[1024]) );
  DFFX1_LVT u_T_427_reg_14__0_ ( .D(n4317), .CLK(n4195), .Q(n_T_427[1023]) );
  DFFX1_LVT u_T_427_reg_15__63_ ( .D(n4495), .CLK(n4194), .Q(n_T_427[1022]) );
  DFFX1_LVT u_T_427_reg_15__62_ ( .D(n4492), .CLK(n4194), .Q(n_T_427[1021]) );
  DFFX1_LVT u_T_427_reg_15__61_ ( .D(n4489), .CLK(n4194), .Q(n_T_427[1020]) );
  DFFX1_LVT u_T_427_reg_15__60_ ( .D(n4486), .CLK(n4194), .Q(n_T_427[1019]) );
  DFFX1_LVT u_T_427_reg_15__59_ ( .D(n4483), .CLK(n4193), .Q(n_T_427[1018]) );
  DFFX1_LVT u_T_427_reg_15__58_ ( .D(n4480), .CLK(n4193), .Q(n_T_427[1017]) );
  DFFX1_LVT u_T_427_reg_15__57_ ( .D(n4477), .CLK(n4193), .Q(n_T_427[1016]) );
  DFFX1_LVT u_T_427_reg_15__56_ ( .D(n4474), .CLK(n4193), .Q(n_T_427[1015]) );
  DFFX1_LVT u_T_427_reg_15__55_ ( .D(n4471), .CLK(n4193), .Q(n_T_427[1014]) );
  DFFX1_LVT u_T_427_reg_15__54_ ( .D(n4468), .CLK(n4193), .Q(n_T_427[1013]) );
  DFFX1_LVT u_T_427_reg_15__53_ ( .D(n4465), .CLK(n4193), .Q(n_T_427[1012]) );
  DFFX1_LVT u_T_427_reg_15__52_ ( .D(n4462), .CLK(n4193), .Q(n_T_427[1011]) );
  DFFX1_LVT u_T_427_reg_15__51_ ( .D(n4459), .CLK(n4193), .Q(n_T_427[1010]) );
  DFFX1_LVT u_T_427_reg_15__50_ ( .D(n4456), .CLK(n4193), .Q(n_T_427[1009]) );
  DFFX1_LVT u_T_427_reg_15__49_ ( .D(n4453), .CLK(n4193), .Q(n_T_427[1008]) );
  DFFX1_LVT u_T_427_reg_15__48_ ( .D(n4450), .CLK(n4193), .Q(n_T_427[1007]) );
  DFFX1_LVT u_T_427_reg_15__47_ ( .D(n4447), .CLK(n4192), .Q(n_T_427[1006]) );
  DFFX1_LVT u_T_427_reg_15__46_ ( .D(n4444), .CLK(n4192), .Q(n_T_427[1005]) );
  DFFX1_LVT u_T_427_reg_15__45_ ( .D(n4441), .CLK(n4192), .Q(n_T_427[1004]) );
  DFFX1_LVT u_T_427_reg_15__44_ ( .D(n4438), .CLK(n4192), .Q(n_T_427[1003]) );
  DFFX1_LVT u_T_427_reg_15__43_ ( .D(n4435), .CLK(n4192), .Q(n_T_427[1002]) );
  DFFX1_LVT u_T_427_reg_15__42_ ( .D(n4432), .CLK(n4192), .Q(n_T_427[1001]) );
  DFFX1_LVT u_T_427_reg_15__41_ ( .D(n4429), .CLK(n4192), .Q(n_T_427[1000]) );
  DFFX1_LVT u_T_427_reg_15__40_ ( .D(n4426), .CLK(n4192), .Q(n_T_427[999]) );
  DFFX1_LVT u_T_427_reg_15__39_ ( .D(n4423), .CLK(n4192), .Q(n_T_427[998]) );
  DFFX1_LVT u_T_427_reg_15__38_ ( .D(n4420), .CLK(n4192), .Q(n_T_427[997]) );
  DFFX1_LVT u_T_427_reg_15__37_ ( .D(n4418), .CLK(n4192), .Q(n_T_427[996]) );
  DFFX1_LVT u_T_427_reg_15__36_ ( .D(n4415), .CLK(n4192), .Q(n_T_427[995]) );
  DFFX1_LVT u_T_427_reg_15__35_ ( .D(n4412), .CLK(n4191), .Q(n_T_427[994]) );
  DFFX1_LVT u_T_427_reg_15__34_ ( .D(n4410), .CLK(n4191), .Q(n_T_427[993]) );
  DFFX1_LVT u_T_427_reg_15__33_ ( .D(n4407), .CLK(n4191), .Q(n_T_427[992]) );
  DFFX1_LVT u_T_427_reg_15__32_ ( .D(n4405), .CLK(n4191), .Q(n_T_427[991]) );
  DFFX1_LVT u_T_427_reg_15__31_ ( .D(n4402), .CLK(n4191), .Q(n_T_427[990]) );
  DFFX1_LVT u_T_427_reg_15__30_ ( .D(n4400), .CLK(n4191), .Q(n_T_427[989]) );
  DFFX1_LVT u_T_427_reg_15__29_ ( .D(n4397), .CLK(n4191), .Q(n_T_427[988]) );
  DFFX1_LVT u_T_427_reg_15__28_ ( .D(n4394), .CLK(n4191), .Q(n_T_427[987]) );
  DFFX1_LVT u_T_427_reg_15__27_ ( .D(n4392), .CLK(n4191), .Q(n_T_427[986]) );
  DFFX1_LVT u_T_427_reg_15__26_ ( .D(n4389), .CLK(n4191), .Q(n_T_427[985]) );
  DFFX1_LVT u_T_427_reg_15__25_ ( .D(n4387), .CLK(n4191), .Q(n_T_427[984]) );
  DFFX1_LVT u_T_427_reg_15__24_ ( .D(n4385), .CLK(n4191), .Q(n_T_427[983]) );
  DFFX1_LVT u_T_427_reg_15__23_ ( .D(n4382), .CLK(n4190), .Q(n_T_427[982]) );
  DFFX1_LVT u_T_427_reg_15__22_ ( .D(n4379), .CLK(n4190), .Q(n_T_427[981]) );
  DFFX1_LVT u_T_427_reg_15__21_ ( .D(n4377), .CLK(n4190), .Q(n_T_427[980]) );
  DFFX1_LVT u_T_427_reg_15__20_ ( .D(n4375), .CLK(n4190), .Q(n_T_427[979]) );
  DFFX1_LVT u_T_427_reg_15__19_ ( .D(n4372), .CLK(n4190), .Q(n_T_427[978]) );
  DFFX1_LVT u_T_427_reg_15__18_ ( .D(n4369), .CLK(n4190), .Q(n_T_427[977]) );
  DFFX1_LVT u_T_427_reg_15__17_ ( .D(n4366), .CLK(n4190), .Q(n_T_427[976]) );
  DFFX1_LVT u_T_427_reg_15__16_ ( .D(n4363), .CLK(n4190), .Q(n_T_427[975]) );
  DFFX1_LVT u_T_427_reg_15__15_ ( .D(n4360), .CLK(n4190), .Q(n_T_427[974]) );
  DFFX1_LVT u_T_427_reg_15__14_ ( .D(n4358), .CLK(n4190), .Q(n_T_427[973]) );
  DFFX1_LVT u_T_427_reg_15__13_ ( .D(n4355), .CLK(n4190), .Q(n_T_427[972]) );
  DFFX1_LVT u_T_427_reg_15__12_ ( .D(n4353), .CLK(n4190), .Q(n_T_427[971]) );
  DFFX1_LVT u_T_427_reg_15__11_ ( .D(n4350), .CLK(n4189), .Q(n_T_427[970]) );
  DFFX1_LVT u_T_427_reg_15__10_ ( .D(n4347), .CLK(n4189), .Q(n_T_427[969]) );
  DFFX1_LVT u_T_427_reg_15__9_ ( .D(n4344), .CLK(n4189), .Q(n_T_427[968]) );
  DFFX1_LVT u_T_427_reg_15__8_ ( .D(n4341), .CLK(n4189), .Q(n_T_427[967]) );
  DFFX1_LVT u_T_427_reg_15__7_ ( .D(n4338), .CLK(n4189), .Q(n_T_427[966]) );
  DFFX1_LVT u_T_427_reg_15__6_ ( .D(n4335), .CLK(n4189), .Q(n_T_427[965]) );
  DFFX1_LVT u_T_427_reg_15__5_ ( .D(n4332), .CLK(n4189), .Q(n_T_427[964]) );
  DFFX1_LVT u_T_427_reg_15__4_ ( .D(n4329), .CLK(n4189), .Q(n_T_427[963]) );
  DFFX1_LVT u_T_427_reg_15__3_ ( .D(n4326), .CLK(n4189), .Q(n_T_427[962]) );
  DFFX1_LVT u_T_427_reg_15__2_ ( .D(n4323), .CLK(n4189), .Q(n_T_427[961]) );
  DFFX1_LVT u_T_427_reg_15__1_ ( .D(n4320), .CLK(n4189), .Q(n_T_427[960]) );
  DFFX1_LVT u_T_427_reg_15__0_ ( .D(n4317), .CLK(n4189), .Q(n_T_427[959]) );
  DFFX1_LVT u_T_427_reg_16__63_ ( .D(n4495), .CLK(n4188), .Q(n_T_427[958]) );
  DFFX1_LVT u_T_427_reg_16__62_ ( .D(n4492), .CLK(n4188), .Q(n_T_427[957]) );
  DFFX1_LVT u_T_427_reg_16__61_ ( .D(n4489), .CLK(n4188), .Q(n_T_427[956]) );
  DFFX1_LVT u_T_427_reg_16__60_ ( .D(n4486), .CLK(n4188), .Q(n_T_427[955]) );
  DFFX1_LVT u_T_427_reg_16__59_ ( .D(n4483), .CLK(n4187), .Q(n_T_427[954]) );
  DFFX1_LVT u_T_427_reg_16__58_ ( .D(n4480), .CLK(n4187), .Q(n_T_427[953]) );
  DFFX1_LVT u_T_427_reg_16__57_ ( .D(n4477), .CLK(n4187), .Q(n_T_427[952]) );
  DFFX1_LVT u_T_427_reg_16__56_ ( .D(n4474), .CLK(n4187), .Q(n_T_427[951]) );
  DFFX1_LVT u_T_427_reg_16__55_ ( .D(n4471), .CLK(n4187), .Q(n_T_427[950]) );
  DFFX1_LVT u_T_427_reg_16__54_ ( .D(n4468), .CLK(n4187), .Q(n_T_427[949]) );
  DFFX1_LVT u_T_427_reg_16__53_ ( .D(n4465), .CLK(n4187), .Q(n_T_427[948]) );
  DFFX1_LVT u_T_427_reg_16__52_ ( .D(n4462), .CLK(n4187), .Q(n_T_427[947]) );
  DFFX1_LVT u_T_427_reg_16__51_ ( .D(n4459), .CLK(n4187), .Q(n_T_427[946]) );
  DFFX1_LVT u_T_427_reg_16__50_ ( .D(n4456), .CLK(n4187), .Q(n_T_427[945]) );
  DFFX1_LVT u_T_427_reg_16__49_ ( .D(n4453), .CLK(n4187), .Q(n_T_427[944]) );
  DFFX1_LVT u_T_427_reg_16__48_ ( .D(n4450), .CLK(n4187), .Q(n_T_427[943]) );
  DFFX1_LVT u_T_427_reg_16__47_ ( .D(n4447), .CLK(n4186), .Q(n_T_427[942]) );
  DFFX1_LVT u_T_427_reg_16__46_ ( .D(n4444), .CLK(n4186), .Q(n_T_427[941]) );
  DFFX1_LVT u_T_427_reg_16__45_ ( .D(n4441), .CLK(n4186), .Q(n_T_427[940]) );
  DFFX1_LVT u_T_427_reg_16__44_ ( .D(n4438), .CLK(n4186), .Q(n_T_427[939]) );
  DFFX1_LVT u_T_427_reg_16__43_ ( .D(n4435), .CLK(n4186), .Q(n_T_427[938]) );
  DFFX1_LVT u_T_427_reg_16__42_ ( .D(n4432), .CLK(n4186), .Q(n_T_427[937]) );
  DFFX1_LVT u_T_427_reg_16__41_ ( .D(n4429), .CLK(n4186), .Q(n_T_427[936]) );
  DFFX1_LVT u_T_427_reg_16__40_ ( .D(n4426), .CLK(n4186), .Q(n_T_427[935]) );
  DFFX1_LVT u_T_427_reg_16__39_ ( .D(n4423), .CLK(n4186), .Q(n_T_427[934]) );
  DFFX1_LVT u_T_427_reg_16__38_ ( .D(n4420), .CLK(n4186), .Q(n_T_427[933]) );
  DFFX1_LVT u_T_427_reg_16__37_ ( .D(n4418), .CLK(n4186), .Q(n_T_427[932]) );
  DFFX1_LVT u_T_427_reg_16__36_ ( .D(n4415), .CLK(n4186), .Q(n_T_427[931]) );
  DFFX1_LVT u_T_427_reg_16__35_ ( .D(n4412), .CLK(n4185), .Q(n_T_427[930]) );
  DFFX1_LVT u_T_427_reg_16__34_ ( .D(n4410), .CLK(n4185), .Q(n_T_427[929]) );
  DFFX1_LVT u_T_427_reg_16__33_ ( .D(n4407), .CLK(n4185), .Q(n_T_427[928]) );
  DFFX1_LVT u_T_427_reg_16__32_ ( .D(n4405), .CLK(n4185), .Q(n_T_427[927]) );
  DFFX1_LVT u_T_427_reg_16__31_ ( .D(n4402), .CLK(n4185), .Q(n_T_427[926]) );
  DFFX1_LVT u_T_427_reg_16__30_ ( .D(n4400), .CLK(n4185), .Q(n_T_427[925]) );
  DFFX1_LVT u_T_427_reg_16__29_ ( .D(n4397), .CLK(n4185), .Q(n_T_427[924]) );
  DFFX1_LVT u_T_427_reg_16__28_ ( .D(n4394), .CLK(n4185), .Q(n_T_427[923]) );
  DFFX1_LVT u_T_427_reg_16__27_ ( .D(n4392), .CLK(n4185), .Q(n_T_427[922]) );
  DFFX1_LVT u_T_427_reg_16__26_ ( .D(n4389), .CLK(n4185), .Q(n_T_427[921]) );
  DFFX1_LVT u_T_427_reg_16__25_ ( .D(n4387), .CLK(n4185), .Q(n_T_427[920]) );
  DFFX1_LVT u_T_427_reg_16__24_ ( .D(n4385), .CLK(n4185), .Q(n_T_427[919]) );
  DFFX1_LVT u_T_427_reg_16__23_ ( .D(n4382), .CLK(n4184), .Q(n_T_427[918]) );
  DFFX1_LVT u_T_427_reg_16__22_ ( .D(n4379), .CLK(n4184), .Q(n_T_427[917]) );
  DFFX1_LVT u_T_427_reg_16__21_ ( .D(n4377), .CLK(n4184), .Q(n_T_427[916]) );
  DFFX1_LVT u_T_427_reg_16__20_ ( .D(n4375), .CLK(n4184), .Q(n_T_427[915]) );
  DFFX1_LVT u_T_427_reg_16__19_ ( .D(n4372), .CLK(n4184), .Q(n_T_427[914]) );
  DFFX1_LVT u_T_427_reg_16__18_ ( .D(n4369), .CLK(n4184), .Q(n_T_427[913]) );
  DFFX1_LVT u_T_427_reg_16__17_ ( .D(n4366), .CLK(n4184), .Q(n_T_427[912]) );
  DFFX1_LVT u_T_427_reg_16__16_ ( .D(n4363), .CLK(n4184), .Q(n_T_427[911]) );
  DFFX1_LVT u_T_427_reg_16__15_ ( .D(n4360), .CLK(n4184), .Q(n_T_427[910]) );
  DFFX1_LVT u_T_427_reg_16__14_ ( .D(n4358), .CLK(n4184), .Q(n_T_427[909]) );
  DFFX1_LVT u_T_427_reg_16__13_ ( .D(n4355), .CLK(n4184), .Q(n_T_427[908]) );
  DFFX1_LVT u_T_427_reg_16__12_ ( .D(n4353), .CLK(n4184), .Q(n_T_427[907]) );
  DFFX1_LVT u_T_427_reg_16__11_ ( .D(n4350), .CLK(n4183), .Q(n_T_427[906]) );
  DFFX1_LVT u_T_427_reg_16__10_ ( .D(n4347), .CLK(n4183), .Q(n_T_427[905]) );
  DFFX1_LVT u_T_427_reg_16__9_ ( .D(n4344), .CLK(n4183), .Q(n_T_427[904]) );
  DFFX1_LVT u_T_427_reg_16__8_ ( .D(n4341), .CLK(n4183), .Q(n_T_427[903]) );
  DFFX1_LVT u_T_427_reg_16__7_ ( .D(n4338), .CLK(n4183), .Q(n_T_427[902]) );
  DFFX1_LVT u_T_427_reg_16__6_ ( .D(n4335), .CLK(n4183), .Q(n_T_427[901]) );
  DFFX1_LVT u_T_427_reg_16__5_ ( .D(n4332), .CLK(n4183), .Q(n_T_427[900]) );
  DFFX1_LVT u_T_427_reg_16__4_ ( .D(n4329), .CLK(n4183), .Q(n_T_427[899]) );
  DFFX1_LVT u_T_427_reg_16__3_ ( .D(n4326), .CLK(n4183), .Q(n_T_427[898]) );
  DFFX1_LVT u_T_427_reg_16__2_ ( .D(n4323), .CLK(n4183), .Q(n_T_427[897]) );
  DFFX1_LVT u_T_427_reg_16__1_ ( .D(n4320), .CLK(n4183), .Q(n_T_427[896]) );
  DFFX1_LVT u_T_427_reg_16__0_ ( .D(n4317), .CLK(n4183), .Q(n_T_427[895]) );
  DFFX1_LVT u_T_427_reg_17__63_ ( .D(n4495), .CLK(n4182), .Q(n_T_427[894]) );
  DFFX1_LVT u_T_427_reg_17__62_ ( .D(n4492), .CLK(n4182), .Q(n_T_427[893]) );
  DFFX1_LVT u_T_427_reg_17__61_ ( .D(n4489), .CLK(n4182), .Q(n_T_427[892]) );
  DFFX1_LVT u_T_427_reg_17__60_ ( .D(n4486), .CLK(n4182), .Q(n_T_427[891]) );
  DFFX1_LVT u_T_427_reg_17__59_ ( .D(n4483), .CLK(n4181), .Q(n_T_427[890]) );
  DFFX1_LVT u_T_427_reg_17__58_ ( .D(n4480), .CLK(n4181), .Q(n_T_427[889]) );
  DFFX1_LVT u_T_427_reg_17__57_ ( .D(n4477), .CLK(n4181), .Q(n_T_427[888]) );
  DFFX1_LVT u_T_427_reg_17__56_ ( .D(n4474), .CLK(n4181), .Q(n_T_427[887]) );
  DFFX1_LVT u_T_427_reg_17__55_ ( .D(n4471), .CLK(n4181), .Q(n_T_427[886]) );
  DFFX1_LVT u_T_427_reg_17__54_ ( .D(n4468), .CLK(n4181), .Q(n_T_427[885]) );
  DFFX1_LVT u_T_427_reg_17__53_ ( .D(n4465), .CLK(n4181), .Q(n_T_427[884]) );
  DFFX1_LVT u_T_427_reg_17__52_ ( .D(n4462), .CLK(n4181), .Q(n_T_427[883]) );
  DFFX1_LVT u_T_427_reg_17__51_ ( .D(n4459), .CLK(n4181), .Q(n_T_427[882]) );
  DFFX1_LVT u_T_427_reg_17__50_ ( .D(n4456), .CLK(n4181), .Q(n_T_427[881]) );
  DFFX1_LVT u_T_427_reg_17__49_ ( .D(n4453), .CLK(n4181), .Q(n_T_427[880]) );
  DFFX1_LVT u_T_427_reg_17__48_ ( .D(n4450), .CLK(n4181), .Q(n_T_427[879]) );
  DFFX1_LVT u_T_427_reg_17__47_ ( .D(n4447), .CLK(n4180), .Q(n_T_427[878]) );
  DFFX1_LVT u_T_427_reg_17__46_ ( .D(n4444), .CLK(n4180), .Q(n_T_427[877]) );
  DFFX1_LVT u_T_427_reg_17__45_ ( .D(n4441), .CLK(n4180), .Q(n_T_427[876]) );
  DFFX1_LVT u_T_427_reg_17__44_ ( .D(n4438), .CLK(n4180), .Q(n_T_427[875]) );
  DFFX1_LVT u_T_427_reg_17__43_ ( .D(n4435), .CLK(n4180), .Q(n_T_427[874]) );
  DFFX1_LVT u_T_427_reg_17__42_ ( .D(n4432), .CLK(n4180), .Q(n_T_427[873]) );
  DFFX1_LVT u_T_427_reg_17__41_ ( .D(n4429), .CLK(n4180), .Q(n_T_427[872]) );
  DFFX1_LVT u_T_427_reg_17__40_ ( .D(n4426), .CLK(n4180), .Q(n_T_427[871]) );
  DFFX1_LVT u_T_427_reg_17__39_ ( .D(n4423), .CLK(n4180), .Q(n_T_427[870]) );
  DFFX1_LVT u_T_427_reg_17__38_ ( .D(n4420), .CLK(n4180), .Q(n_T_427[869]) );
  DFFX1_LVT u_T_427_reg_17__37_ ( .D(n4418), .CLK(n4180), .Q(n_T_427[868]) );
  DFFX1_LVT u_T_427_reg_17__36_ ( .D(n4415), .CLK(n4180), .Q(n_T_427[867]) );
  DFFX1_LVT u_T_427_reg_17__35_ ( .D(n4412), .CLK(n4179), .Q(n_T_427[866]) );
  DFFX1_LVT u_T_427_reg_17__34_ ( .D(n4410), .CLK(n4179), .Q(n_T_427[865]) );
  DFFX1_LVT u_T_427_reg_17__33_ ( .D(n4407), .CLK(n4179), .Q(n_T_427[864]) );
  DFFX1_LVT u_T_427_reg_17__32_ ( .D(n4405), .CLK(n4179), .Q(n_T_427[863]) );
  DFFX1_LVT u_T_427_reg_17__31_ ( .D(n4402), .CLK(n4179), .Q(n_T_427[862]) );
  DFFX1_LVT u_T_427_reg_17__30_ ( .D(n4400), .CLK(n4179), .Q(n_T_427[861]) );
  DFFX1_LVT u_T_427_reg_17__29_ ( .D(n4397), .CLK(n4179), .Q(n_T_427[860]) );
  DFFX1_LVT u_T_427_reg_17__28_ ( .D(n4394), .CLK(n4179), .Q(n_T_427[859]) );
  DFFX1_LVT u_T_427_reg_17__27_ ( .D(n4392), .CLK(n4179), .Q(n_T_427[858]) );
  DFFX1_LVT u_T_427_reg_17__26_ ( .D(n4389), .CLK(n4179), .Q(n_T_427[857]) );
  DFFX1_LVT u_T_427_reg_17__25_ ( .D(n4387), .CLK(n4179), .Q(n_T_427[856]) );
  DFFX1_LVT u_T_427_reg_17__24_ ( .D(n4385), .CLK(n4179), .Q(n_T_427[855]) );
  DFFX1_LVT u_T_427_reg_17__23_ ( .D(n4382), .CLK(n4178), .Q(n_T_427[854]) );
  DFFX1_LVT u_T_427_reg_17__22_ ( .D(n4379), .CLK(n4178), .Q(n_T_427[853]) );
  DFFX1_LVT u_T_427_reg_17__21_ ( .D(n4377), .CLK(n4178), .Q(n_T_427[852]) );
  DFFX1_LVT u_T_427_reg_17__20_ ( .D(n4375), .CLK(n4178), .Q(n_T_427[851]) );
  DFFX1_LVT u_T_427_reg_17__19_ ( .D(n4372), .CLK(n4178), .Q(n_T_427[850]) );
  DFFX1_LVT u_T_427_reg_17__18_ ( .D(n4369), .CLK(n4178), .Q(n_T_427[849]) );
  DFFX1_LVT u_T_427_reg_17__17_ ( .D(n4366), .CLK(n4178), .Q(n_T_427[848]) );
  DFFX1_LVT u_T_427_reg_17__16_ ( .D(n4363), .CLK(n4178), .Q(n_T_427[847]) );
  DFFX1_LVT u_T_427_reg_17__15_ ( .D(n4360), .CLK(n4178), .Q(n_T_427[846]) );
  DFFX1_LVT u_T_427_reg_17__14_ ( .D(n4358), .CLK(n4178), .Q(n_T_427[845]) );
  DFFX1_LVT u_T_427_reg_17__13_ ( .D(n4355), .CLK(n4178), .Q(n_T_427[844]) );
  DFFX1_LVT u_T_427_reg_17__12_ ( .D(n4353), .CLK(n4178), .Q(n_T_427[843]) );
  DFFX1_LVT u_T_427_reg_17__11_ ( .D(n4350), .CLK(n4177), .Q(n_T_427[842]) );
  DFFX1_LVT u_T_427_reg_17__10_ ( .D(n4347), .CLK(n4177), .Q(n_T_427[841]) );
  DFFX1_LVT u_T_427_reg_17__9_ ( .D(n4344), .CLK(n4177), .Q(n_T_427[840]) );
  DFFX1_LVT u_T_427_reg_17__8_ ( .D(n4341), .CLK(n4177), .Q(n_T_427[839]) );
  DFFX1_LVT u_T_427_reg_17__7_ ( .D(n4338), .CLK(n4177), .Q(n_T_427[838]) );
  DFFX1_LVT u_T_427_reg_17__6_ ( .D(n4335), .CLK(n4177), .Q(n_T_427[837]) );
  DFFX1_LVT u_T_427_reg_17__5_ ( .D(n4332), .CLK(n4177), .Q(n_T_427[836]) );
  DFFX1_LVT u_T_427_reg_17__4_ ( .D(n4329), .CLK(n4177), .Q(n_T_427[835]) );
  DFFX1_LVT u_T_427_reg_17__3_ ( .D(n4326), .CLK(n4177), .Q(n_T_427[834]) );
  DFFX1_LVT u_T_427_reg_17__2_ ( .D(n4323), .CLK(n4177), .Q(n_T_427[833]) );
  DFFX1_LVT u_T_427_reg_17__1_ ( .D(n4320), .CLK(n4177), .Q(n_T_427[832]) );
  DFFX1_LVT u_T_427_reg_17__0_ ( .D(n4317), .CLK(n4177), .Q(n_T_427[831]) );
  DFFX1_LVT u_T_427_reg_18__63_ ( .D(n4495), .CLK(n4176), .Q(n_T_427[830]) );
  DFFX1_LVT u_T_427_reg_18__62_ ( .D(n4492), .CLK(n4176), .Q(n_T_427[829]) );
  DFFX1_LVT u_T_427_reg_18__61_ ( .D(n4489), .CLK(n4176), .Q(n_T_427[828]) );
  DFFX1_LVT u_T_427_reg_18__60_ ( .D(n4486), .CLK(n4176), .Q(n_T_427[827]) );
  DFFX1_LVT u_T_427_reg_18__59_ ( .D(n4483), .CLK(n4175), .Q(n_T_427[826]) );
  DFFX1_LVT u_T_427_reg_18__58_ ( .D(n4480), .CLK(n4175), .Q(n_T_427[825]) );
  DFFX1_LVT u_T_427_reg_18__57_ ( .D(n4477), .CLK(n4175), .Q(n_T_427[824]) );
  DFFX1_LVT u_T_427_reg_18__56_ ( .D(n4474), .CLK(n4175), .Q(n_T_427[823]) );
  DFFX1_LVT u_T_427_reg_18__55_ ( .D(n4471), .CLK(n4175), .Q(n_T_427[822]) );
  DFFX1_LVT u_T_427_reg_18__54_ ( .D(n4468), .CLK(n4175), .Q(n_T_427[821]) );
  DFFX1_LVT u_T_427_reg_18__53_ ( .D(n4465), .CLK(n4175), .Q(n_T_427[820]) );
  DFFX1_LVT u_T_427_reg_18__52_ ( .D(n4462), .CLK(n4175), .Q(n_T_427[819]) );
  DFFX1_LVT u_T_427_reg_18__51_ ( .D(n4459), .CLK(n4175), .Q(n_T_427[818]) );
  DFFX1_LVT u_T_427_reg_18__50_ ( .D(n4456), .CLK(n4175), .Q(n_T_427[817]) );
  DFFX1_LVT u_T_427_reg_18__49_ ( .D(n4453), .CLK(n4175), .Q(n_T_427[816]) );
  DFFX1_LVT u_T_427_reg_18__48_ ( .D(n4450), .CLK(n4175), .Q(n_T_427[815]) );
  DFFX1_LVT u_T_427_reg_18__47_ ( .D(n4447), .CLK(n4174), .Q(n_T_427[814]) );
  DFFX1_LVT u_T_427_reg_18__46_ ( .D(n4444), .CLK(n4174), .Q(n_T_427[813]) );
  DFFX1_LVT u_T_427_reg_18__45_ ( .D(n4441), .CLK(n4174), .Q(n_T_427[812]) );
  DFFX1_LVT u_T_427_reg_18__44_ ( .D(n4438), .CLK(n4174), .Q(n_T_427[811]) );
  DFFX1_LVT u_T_427_reg_18__43_ ( .D(n4435), .CLK(n4174), .Q(n_T_427[810]) );
  DFFX1_LVT u_T_427_reg_18__42_ ( .D(n4432), .CLK(n4174), .Q(n_T_427[809]) );
  DFFX1_LVT u_T_427_reg_18__41_ ( .D(n4429), .CLK(n4174), .Q(n_T_427[808]) );
  DFFX1_LVT u_T_427_reg_18__40_ ( .D(n4426), .CLK(n4174), .Q(n_T_427[807]) );
  DFFX1_LVT u_T_427_reg_18__39_ ( .D(n4423), .CLK(n4174), .Q(n_T_427[806]) );
  DFFX1_LVT u_T_427_reg_18__38_ ( .D(n4420), .CLK(n4174), .Q(n_T_427[805]) );
  DFFX1_LVT u_T_427_reg_18__37_ ( .D(n4418), .CLK(n4174), .Q(n_T_427[804]) );
  DFFX1_LVT u_T_427_reg_18__36_ ( .D(n4415), .CLK(n4174), .Q(n_T_427[803]) );
  DFFX1_LVT u_T_427_reg_18__35_ ( .D(n4412), .CLK(n4173), .Q(n_T_427[802]) );
  DFFX1_LVT u_T_427_reg_18__34_ ( .D(n4410), .CLK(n4173), .Q(n_T_427[801]) );
  DFFX1_LVT u_T_427_reg_18__33_ ( .D(n4407), .CLK(n4173), .Q(n_T_427[800]) );
  DFFX1_LVT u_T_427_reg_18__32_ ( .D(n4405), .CLK(n4173), .Q(n_T_427[799]) );
  DFFX1_LVT u_T_427_reg_18__31_ ( .D(n4402), .CLK(n4173), .Q(n_T_427[798]) );
  DFFX1_LVT u_T_427_reg_18__30_ ( .D(n4400), .CLK(n4173), .Q(n_T_427[797]) );
  DFFX1_LVT u_T_427_reg_18__29_ ( .D(n4397), .CLK(n4173), .Q(n_T_427[796]) );
  DFFX1_LVT u_T_427_reg_18__28_ ( .D(n4394), .CLK(n4173), .Q(n_T_427[795]) );
  DFFX1_LVT u_T_427_reg_18__27_ ( .D(n4392), .CLK(n4173), .Q(n_T_427[794]) );
  DFFX1_LVT u_T_427_reg_18__26_ ( .D(n4389), .CLK(n4173), .Q(n_T_427[793]) );
  DFFX1_LVT u_T_427_reg_18__25_ ( .D(n4387), .CLK(n4173), .Q(n_T_427[792]) );
  DFFX1_LVT u_T_427_reg_18__24_ ( .D(n4385), .CLK(n4173), .Q(n_T_427[791]) );
  DFFX1_LVT u_T_427_reg_18__23_ ( .D(n4382), .CLK(n4172), .Q(n_T_427[790]) );
  DFFX1_LVT u_T_427_reg_18__22_ ( .D(n4379), .CLK(n4172), .Q(n_T_427[789]) );
  DFFX1_LVT u_T_427_reg_18__21_ ( .D(n4377), .CLK(n4172), .Q(n_T_427[788]) );
  DFFX1_LVT u_T_427_reg_18__20_ ( .D(n4375), .CLK(n4172), .Q(n_T_427[787]) );
  DFFX1_LVT u_T_427_reg_18__19_ ( .D(n4372), .CLK(n4172), .Q(n_T_427[786]) );
  DFFX1_LVT u_T_427_reg_18__18_ ( .D(n4369), .CLK(n4172), .Q(n_T_427[785]) );
  DFFX1_LVT u_T_427_reg_18__17_ ( .D(n4366), .CLK(n4172), .Q(n_T_427[784]) );
  DFFX1_LVT u_T_427_reg_18__16_ ( .D(n4363), .CLK(n4172), .Q(n_T_427[783]) );
  DFFX1_LVT u_T_427_reg_18__15_ ( .D(n4360), .CLK(n4172), .Q(n_T_427[782]) );
  DFFX1_LVT u_T_427_reg_18__14_ ( .D(n4358), .CLK(n4172), .Q(n_T_427[781]) );
  DFFX1_LVT u_T_427_reg_18__13_ ( .D(n4355), .CLK(n4172), .Q(n_T_427[780]) );
  DFFX1_LVT u_T_427_reg_18__12_ ( .D(n4353), .CLK(n4172), .Q(n_T_427[779]) );
  DFFX1_LVT u_T_427_reg_18__11_ ( .D(n4350), .CLK(n4171), .Q(n_T_427[778]) );
  DFFX1_LVT u_T_427_reg_18__10_ ( .D(n4347), .CLK(n4171), .Q(n_T_427[777]) );
  DFFX1_LVT u_T_427_reg_18__9_ ( .D(n4344), .CLK(n4171), .Q(n_T_427[776]) );
  DFFX1_LVT u_T_427_reg_18__8_ ( .D(n4341), .CLK(n4171), .Q(n_T_427[775]) );
  DFFX1_LVT u_T_427_reg_18__7_ ( .D(n4338), .CLK(n4171), .Q(n_T_427[774]) );
  DFFX1_LVT u_T_427_reg_18__6_ ( .D(n4335), .CLK(n4171), .Q(n_T_427[773]) );
  DFFX1_LVT u_T_427_reg_18__5_ ( .D(n4332), .CLK(n4171), .Q(n_T_427[772]) );
  DFFX1_LVT u_T_427_reg_18__4_ ( .D(n4329), .CLK(n4171), .Q(n_T_427[771]) );
  DFFX1_LVT u_T_427_reg_18__3_ ( .D(n4326), .CLK(n4171), .Q(n_T_427[770]) );
  DFFX1_LVT u_T_427_reg_18__2_ ( .D(n4323), .CLK(n4171), .Q(n_T_427[769]) );
  DFFX1_LVT u_T_427_reg_18__1_ ( .D(n4320), .CLK(n4171), .Q(n_T_427[768]) );
  DFFX1_LVT u_T_427_reg_18__0_ ( .D(n4317), .CLK(n4171), .Q(n_T_427[767]) );
  DFFX1_LVT u_T_427_reg_19__63_ ( .D(n4495), .CLK(n4170), .Q(n_T_427[766]) );
  DFFX1_LVT u_T_427_reg_19__62_ ( .D(n4492), .CLK(n4170), .Q(n_T_427[765]) );
  DFFX1_LVT u_T_427_reg_19__61_ ( .D(n4489), .CLK(n4170), .Q(n_T_427[764]), 
        .QN(n3280) );
  DFFX1_LVT u_T_427_reg_19__60_ ( .D(n4486), .CLK(n4170), .Q(n_T_427[763]) );
  DFFX1_LVT u_T_427_reg_19__59_ ( .D(n4483), .CLK(n4169), .Q(n_T_427[762]) );
  DFFX1_LVT u_T_427_reg_19__58_ ( .D(n4479), .CLK(n4169), .Q(n_T_427[761]) );
  DFFX1_LVT u_T_427_reg_19__56_ ( .D(n4473), .CLK(n4169), .Q(n_T_427[759]) );
  DFFX1_LVT u_T_427_reg_19__54_ ( .D(n4467), .CLK(n4169), .Q(n_T_427[757]) );
  DFFX1_LVT u_T_427_reg_19__53_ ( .D(n4465), .CLK(n4169), .Q(n_T_427[756]) );
  DFFX1_LVT u_T_427_reg_19__52_ ( .D(n4461), .CLK(n4169), .Q(n_T_427[755]), 
        .QN(n3408) );
  DFFX1_LVT u_T_427_reg_19__51_ ( .D(n4458), .CLK(n4169), .Q(n_T_427[754]) );
  DFFX1_LVT u_T_427_reg_19__49_ ( .D(n4452), .CLK(n4169), .Q(n_T_427[752]) );
  DFFX1_LVT u_T_427_reg_19__48_ ( .D(n4450), .CLK(n4169), .Q(n_T_427[751]) );
  DFFX1_LVT u_T_427_reg_19__47_ ( .D(n4447), .CLK(n4168), .Q(n_T_427[750]) );
  DFFX1_LVT u_T_427_reg_19__45_ ( .D(n4440), .CLK(n4168), .Q(n_T_427[748]) );
  DFFX1_LVT u_T_427_reg_19__44_ ( .D(n4438), .CLK(n4168), .Q(n_T_427[747]) );
  DFFX1_LVT u_T_427_reg_19__43_ ( .D(n4434), .CLK(n4168), .Q(n_T_427[746]), 
        .QN(n3405) );
  DFFX1_LVT u_T_427_reg_19__42_ ( .D(n4431), .CLK(n4168), .Q(n_T_427[745]) );
  DFFX1_LVT u_T_427_reg_19__41_ ( .D(n4428), .CLK(n4168), .Q(n_T_427[744]) );
  DFFX1_LVT u_T_427_reg_19__39_ ( .D(n4423), .CLK(n4168), .Q(n_T_427[742]) );
  DFFX1_LVT u_T_427_reg_19__38_ ( .D(n4420), .CLK(n4168), .Q(n_T_427[741]) );
  DFFX1_LVT u_T_427_reg_19__37_ ( .D(n4418), .CLK(n4168), .Q(n_T_427[740]) );
  DFFX1_LVT u_T_427_reg_19__36_ ( .D(n4414), .CLK(n4168), .Q(n_T_427[739]) );
  DFFX1_LVT u_T_427_reg_19__33_ ( .D(n4407), .CLK(n4167), .Q(n_T_427[737]) );
  DFFX1_LVT u_T_427_reg_19__31_ ( .D(n4402), .CLK(n4167), .Q(n_T_427[735]) );
  DFFX1_LVT u_T_427_reg_19__30_ ( .D(n4399), .CLK(n4167), .Q(n_T_427[734]) );
  DFFX1_LVT u_T_427_reg_19__29_ ( .D(n4396), .CLK(n4167), .Q(n_T_427[733]) );
  DFFX1_LVT u_T_427_reg_19__28_ ( .D(n4394), .CLK(n4167), .Q(n_T_427[732]) );
  DFFX1_LVT u_T_427_reg_19__27_ ( .D(n4392), .CLK(n4167), .Q(n_T_427[731]) );
  DFFX1_LVT u_T_427_reg_19__26_ ( .D(n4389), .CLK(n4167), .Q(n_T_427[730]) );
  DFFX1_LVT u_T_427_reg_19__25_ ( .D(n4387), .CLK(n4167), .Q(n_T_427[729]) );
  DFFX1_LVT u_T_427_reg_19__24_ ( .D(n4384), .CLK(n4167), .Q(n_T_427[728]) );
  DFFX1_LVT u_T_427_reg_19__23_ ( .D(n4382), .CLK(n4166), .Q(n_T_427[727]) );
  DFFX1_LVT u_T_427_reg_19__22_ ( .D(n4379), .CLK(n4166), .Q(n_T_427[726]) );
  DFFX1_LVT u_T_427_reg_19__21_ ( .D(n4377), .CLK(n4166), .Q(n_T_427[725]) );
  DFFX1_LVT u_T_427_reg_19__20_ ( .D(n4374), .CLK(n4166), .Q(n_T_427[724]) );
  DFFX1_LVT u_T_427_reg_19__19_ ( .D(n4371), .CLK(n4166), .Q(n_T_427[723]) );
  DFFX1_LVT u_T_427_reg_19__18_ ( .D(n4368), .CLK(n4166), .Q(n_T_427[722]) );
  DFFX1_LVT u_T_427_reg_19__17_ ( .D(n4366), .CLK(n4166), .Q(n_T_427[721]) );
  DFFX1_LVT u_T_427_reg_19__16_ ( .D(n4363), .CLK(n4166), .Q(n_T_427[720]) );
  DFFX1_LVT u_T_427_reg_19__15_ ( .D(n4360), .CLK(n4166), .Q(n_T_427[719]) );
  DFFX1_LVT u_T_427_reg_19__14_ ( .D(n4358), .CLK(n4166), .Q(n_T_427[718]) );
  DFFX1_LVT u_T_427_reg_19__13_ ( .D(n4355), .CLK(n4166), .Q(n_T_427[717]) );
  DFFX1_LVT u_T_427_reg_19__12_ ( .D(n4353), .CLK(n4166), .Q(n_T_427[716]) );
  DFFX1_LVT u_T_427_reg_19__11_ ( .D(n4349), .CLK(n4165), .Q(n_T_427[715]) );
  DFFX1_LVT u_T_427_reg_19__10_ ( .D(n4347), .CLK(n4165), .Q(n_T_427[714]) );
  DFFX1_LVT u_T_427_reg_19__9_ ( .D(n4344), .CLK(n4165), .Q(n_T_427[713]) );
  DFFX1_LVT u_T_427_reg_19__8_ ( .D(n4341), .CLK(n4165), .Q(n_T_427[712]) );
  DFFX1_LVT u_T_427_reg_19__7_ ( .D(n4338), .CLK(n4165), .Q(n_T_427[711]) );
  DFFX1_LVT u_T_427_reg_19__6_ ( .D(n4335), .CLK(n4165), .Q(n_T_427[710]) );
  DFFX1_LVT u_T_427_reg_19__5_ ( .D(n4332), .CLK(n4165), .Q(n_T_427[709]) );
  DFFX1_LVT u_T_427_reg_19__4_ ( .D(n4329), .CLK(n4165), .Q(n_T_427[708]) );
  DFFX1_LVT u_T_427_reg_19__3_ ( .D(n4326), .CLK(n4165), .Q(n_T_427[707]) );
  DFFX1_LVT u_T_427_reg_19__2_ ( .D(n4323), .CLK(n4165), .Q(n_T_427[706]) );
  DFFX1_LVT u_T_427_reg_19__1_ ( .D(n4319), .CLK(n4165), .Q(n_T_427[705]) );
  DFFX1_LVT u_T_427_reg_19__0_ ( .D(n4316), .CLK(n4165), .Q(n_T_427[704]) );
  DFFX1_LVT u_T_427_reg_20__63_ ( .D(n4495), .CLK(n4164), .Q(n_T_427[703]) );
  DFFX1_LVT u_T_427_reg_20__62_ ( .D(n4492), .CLK(n4164), .Q(n_T_427[702]), 
        .QN(n3478) );
  DFFX1_LVT u_T_427_reg_20__61_ ( .D(n4489), .CLK(n4164), .Q(n_T_427[701]) );
  DFFX1_LVT u_T_427_reg_20__60_ ( .D(n4486), .CLK(n4164), .Q(n_T_427[700]) );
  DFFX1_LVT u_T_427_reg_20__59_ ( .D(n4483), .CLK(n4163), .Q(n_T_427[699]) );
  DFFX1_LVT u_T_427_reg_20__58_ ( .D(n4479), .CLK(n4163), .Q(n_T_427[698]) );
  DFFX1_LVT u_T_427_reg_20__57_ ( .D(n4477), .CLK(n4163), .Q(n_T_427[697]) );
  DFFX1_LVT u_T_427_reg_20__56_ ( .D(n4473), .CLK(n4163), .Q(n_T_427[696]) );
  DFFX1_LVT u_T_427_reg_20__55_ ( .D(n4471), .CLK(n4163), .Q(n_T_427[695]) );
  DFFX1_LVT u_T_427_reg_20__54_ ( .D(n4467), .CLK(n4163), .Q(n_T_427[694]) );
  DFFX1_LVT u_T_427_reg_20__53_ ( .D(n4465), .CLK(n4163), .Q(n_T_427[693]) );
  DFFX1_LVT u_T_427_reg_20__52_ ( .D(n4461), .CLK(n4163), .Q(n_T_427[692]) );
  DFFX1_LVT u_T_427_reg_20__51_ ( .D(n4458), .CLK(n4163), .Q(n_T_427[691]) );
  DFFX1_LVT u_T_427_reg_20__50_ ( .D(n4456), .CLK(n4163), .Q(n_T_427[690]) );
  DFFX1_LVT u_T_427_reg_20__49_ ( .D(n4452), .CLK(n4163), .Q(n_T_427[689]) );
  DFFX1_LVT u_T_427_reg_20__48_ ( .D(n4450), .CLK(n4163), .Q(n_T_427[688]) );
  DFFX1_LVT u_T_427_reg_20__46_ ( .D(n4444), .CLK(n4162), .Q(n_T_427[686]) );
  DFFX1_LVT u_T_427_reg_20__45_ ( .D(n4440), .CLK(n4162), .Q(n_T_427[685]) );
  DFFX1_LVT u_T_427_reg_20__44_ ( .D(n4438), .CLK(n4162), .Q(n_T_427[684]) );
  DFFX1_LVT u_T_427_reg_20__43_ ( .D(n4434), .CLK(n4162), .Q(n_T_427[683]) );
  DFFX1_LVT u_T_427_reg_20__42_ ( .D(n4431), .CLK(n4162), .Q(n_T_427[682]) );
  DFFX1_LVT u_T_427_reg_20__41_ ( .D(n4428), .CLK(n4162), .Q(n_T_427[681]), 
        .QN(n3404) );
  DFFX1_LVT u_T_427_reg_20__40_ ( .D(n4426), .CLK(n4162), .Q(n_T_427[680]) );
  DFFX1_LVT u_T_427_reg_20__38_ ( .D(n4420), .CLK(n4162), .Q(n_T_427[678]) );
  DFFX1_LVT u_T_427_reg_20__37_ ( .D(n4418), .CLK(n4162), .Q(n_T_427[677]) );
  DFFX1_LVT u_T_427_reg_20__36_ ( .D(n4414), .CLK(n4162), .Q(n_T_427[676]) );
  DFFX1_LVT u_T_427_reg_20__34_ ( .D(n4410), .CLK(n4161), .Q(n_T_427[674]) );
  DFFX1_LVT u_T_427_reg_20__33_ ( .D(n4407), .CLK(n4161), .Q(n_T_427[673]) );
  DFFX1_LVT u_T_427_reg_20__32_ ( .D(n4405), .CLK(n4161), .Q(n_T_427[672]) );
  DFFX1_LVT u_T_427_reg_20__31_ ( .D(n4402), .CLK(n4161), .Q(n_T_427[671]) );
  DFFX1_LVT u_T_427_reg_20__30_ ( .D(n4399), .CLK(n4161), .Q(n_T_427[670]) );
  DFFX1_LVT u_T_427_reg_20__29_ ( .D(n4396), .CLK(n4161), .Q(n_T_427[669]) );
  DFFX1_LVT u_T_427_reg_20__28_ ( .D(n4394), .CLK(n4161), .Q(n_T_427[668]) );
  DFFX1_LVT u_T_427_reg_20__27_ ( .D(n4392), .CLK(n4161), .Q(n_T_427[667]) );
  DFFX1_LVT u_T_427_reg_20__26_ ( .D(n4389), .CLK(n4161), .Q(n_T_427[666]) );
  DFFX1_LVT u_T_427_reg_20__25_ ( .D(n4387), .CLK(n4161), .Q(n_T_427[665]) );
  DFFX1_LVT u_T_427_reg_20__24_ ( .D(n4384), .CLK(n4161), .Q(n_T_427[664]) );
  DFFX1_LVT u_T_427_reg_20__23_ ( .D(n4382), .CLK(n4160), .Q(n_T_427[663]) );
  DFFX1_LVT u_T_427_reg_20__22_ ( .D(n4379), .CLK(n4160), .Q(n_T_427[662]) );
  DFFX1_LVT u_T_427_reg_20__21_ ( .D(n4377), .CLK(n4160), .Q(n_T_427[661]) );
  DFFX1_LVT u_T_427_reg_20__20_ ( .D(n4374), .CLK(n4160), .Q(n_T_427[660]) );
  DFFX1_LVT u_T_427_reg_20__19_ ( .D(n4371), .CLK(n4160), .Q(n_T_427[659]) );
  DFFX1_LVT u_T_427_reg_20__18_ ( .D(n4368), .CLK(n4160), .Q(n_T_427[658]) );
  DFFX1_LVT u_T_427_reg_20__17_ ( .D(n4366), .CLK(n4160), .Q(n_T_427[657]) );
  DFFX1_LVT u_T_427_reg_20__16_ ( .D(n4363), .CLK(n4160), .Q(n_T_427[656]) );
  DFFX1_LVT u_T_427_reg_20__15_ ( .D(n4360), .CLK(n4160), .Q(n_T_427[655]) );
  DFFX1_LVT u_T_427_reg_20__14_ ( .D(n4358), .CLK(n4160), .Q(n_T_427[654]) );
  DFFX1_LVT u_T_427_reg_20__13_ ( .D(n4355), .CLK(n4160), .Q(n_T_427[653]) );
  DFFX1_LVT u_T_427_reg_20__12_ ( .D(n4353), .CLK(n4160), .Q(n_T_427[652]) );
  DFFX1_LVT u_T_427_reg_20__11_ ( .D(n4349), .CLK(n4159), .Q(n_T_427[651]) );
  DFFX1_LVT u_T_427_reg_20__10_ ( .D(n4347), .CLK(n4159), .Q(n_T_427[650]) );
  DFFX1_LVT u_T_427_reg_20__9_ ( .D(n4344), .CLK(n4159), .Q(n_T_427[649]) );
  DFFX1_LVT u_T_427_reg_20__8_ ( .D(n4341), .CLK(n4159), .Q(n_T_427[648]) );
  DFFX1_LVT u_T_427_reg_20__7_ ( .D(n4338), .CLK(n4159), .Q(n_T_427[647]) );
  DFFX1_LVT u_T_427_reg_20__6_ ( .D(n4335), .CLK(n4159), .Q(n_T_427[646]) );
  DFFX1_LVT u_T_427_reg_20__5_ ( .D(n4332), .CLK(n4159), .Q(n_T_427[645]) );
  DFFX1_LVT u_T_427_reg_20__3_ ( .D(n4326), .CLK(n4159), .Q(n_T_427[643]) );
  DFFX1_LVT u_T_427_reg_20__1_ ( .D(n4319), .CLK(n4159), .Q(n_T_427[641]) );
  DFFX1_LVT u_T_427_reg_20__0_ ( .D(n4316), .CLK(n4159), .Q(n_T_427[640]) );
  DFFX1_LVT u_T_427_reg_21__63_ ( .D(n4495), .CLK(n4158), .Q(n_T_427[639]) );
  DFFX1_LVT u_T_427_reg_21__62_ ( .D(n4492), .CLK(n4158), .Q(n_T_427[638]) );
  DFFX1_LVT u_T_427_reg_21__61_ ( .D(n4489), .CLK(n4158), .Q(n_T_427[637]) );
  DFFX1_LVT u_T_427_reg_21__60_ ( .D(n4486), .CLK(n4158), .Q(n_T_427[636]) );
  DFFX1_LVT u_T_427_reg_21__59_ ( .D(n4483), .CLK(n4157), .Q(n_T_427[635]) );
  DFFX1_LVT u_T_427_reg_21__58_ ( .D(n4479), .CLK(n4157), .Q(n_T_427[634]) );
  DFFX1_LVT u_T_427_reg_21__57_ ( .D(n4477), .CLK(n4157), .Q(n_T_427[633]) );
  DFFX1_LVT u_T_427_reg_21__56_ ( .D(n4473), .CLK(n4157), .Q(n_T_427[632]) );
  DFFX1_LVT u_T_427_reg_21__55_ ( .D(n4471), .CLK(n4157), .Q(n_T_427[631]) );
  DFFX1_LVT u_T_427_reg_21__54_ ( .D(n4467), .CLK(n4157), .Q(n_T_427[630]) );
  DFFX1_LVT u_T_427_reg_21__53_ ( .D(n4465), .CLK(n4157), .Q(n_T_427[629]) );
  DFFX1_LVT u_T_427_reg_21__52_ ( .D(n4461), .CLK(n4157), .Q(n_T_427[628]) );
  DFFX1_LVT u_T_427_reg_21__51_ ( .D(n4458), .CLK(n4157), .Q(n_T_427[627]) );
  DFFX1_LVT u_T_427_reg_21__50_ ( .D(n4456), .CLK(n4157), .Q(n_T_427[626]) );
  DFFX1_LVT u_T_427_reg_21__49_ ( .D(n4452), .CLK(n4157), .Q(n_T_427[625]) );
  DFFX1_LVT u_T_427_reg_21__48_ ( .D(n4450), .CLK(n4157), .Q(n_T_427[624]) );
  DFFX1_LVT u_T_427_reg_21__47_ ( .D(n4447), .CLK(n4156), .Q(n_T_427[623]) );
  DFFX1_LVT u_T_427_reg_21__46_ ( .D(n4444), .CLK(n4156), .Q(n_T_427[622]) );
  DFFX1_LVT u_T_427_reg_21__45_ ( .D(n4440), .CLK(n4156), .Q(n_T_427[621]) );
  DFFX1_LVT u_T_427_reg_21__44_ ( .D(n4438), .CLK(n4156), .Q(n_T_427[620]) );
  DFFX1_LVT u_T_427_reg_21__43_ ( .D(n4434), .CLK(n4156), .Q(n_T_427[619]) );
  DFFX1_LVT u_T_427_reg_21__42_ ( .D(n4431), .CLK(n4156), .Q(n_T_427[618]) );
  DFFX1_LVT u_T_427_reg_21__41_ ( .D(n4428), .CLK(n4156), .Q(n_T_427[617]) );
  DFFX1_LVT u_T_427_reg_21__40_ ( .D(n4426), .CLK(n4156), .Q(n_T_427[616]) );
  DFFX1_LVT u_T_427_reg_21__39_ ( .D(n4423), .CLK(n4156), .Q(n_T_427[615]) );
  DFFX1_LVT u_T_427_reg_21__38_ ( .D(n4420), .CLK(n4156), .Q(n_T_427[614]) );
  DFFX1_LVT u_T_427_reg_21__37_ ( .D(n4418), .CLK(n4156), .Q(n_T_427[613]) );
  DFFX1_LVT u_T_427_reg_21__36_ ( .D(n4414), .CLK(n4156), .Q(n_T_427[612]) );
  DFFX1_LVT u_T_427_reg_21__35_ ( .D(n4412), .CLK(n4155), .Q(n_T_427[611]) );
  DFFX1_LVT u_T_427_reg_21__34_ ( .D(n4410), .CLK(n4155), .Q(n_T_427[610]) );
  DFFX1_LVT u_T_427_reg_21__33_ ( .D(n4407), .CLK(n4155), .Q(n_T_427[609]) );
  DFFX1_LVT u_T_427_reg_21__32_ ( .D(n4405), .CLK(n4155), .Q(n_T_427[608]) );
  DFFX1_LVT u_T_427_reg_21__31_ ( .D(n4402), .CLK(n4155), .Q(n_T_427[607]) );
  DFFX1_LVT u_T_427_reg_21__30_ ( .D(n4399), .CLK(n4155), .Q(n_T_427[606]) );
  DFFX1_LVT u_T_427_reg_21__29_ ( .D(n4396), .CLK(n4155), .Q(n_T_427[605]) );
  DFFX1_LVT u_T_427_reg_21__28_ ( .D(n4394), .CLK(n4155), .Q(n_T_427[604]) );
  DFFX1_LVT u_T_427_reg_21__27_ ( .D(n4392), .CLK(n4155), .Q(n_T_427[603]) );
  DFFX1_LVT u_T_427_reg_21__26_ ( .D(n4389), .CLK(n4155), .Q(n_T_427[602]) );
  DFFX1_LVT u_T_427_reg_21__25_ ( .D(n4387), .CLK(n4155), .Q(n_T_427[601]) );
  DFFX1_LVT u_T_427_reg_21__24_ ( .D(n4384), .CLK(n4155), .Q(n_T_427[600]) );
  DFFX1_LVT u_T_427_reg_21__23_ ( .D(n4382), .CLK(n4154), .Q(n_T_427[599]) );
  DFFX1_LVT u_T_427_reg_21__22_ ( .D(n4379), .CLK(n4154), .Q(n_T_427[598]) );
  DFFX1_LVT u_T_427_reg_21__21_ ( .D(n4377), .CLK(n4154), .Q(n_T_427[597]) );
  DFFX1_LVT u_T_427_reg_21__20_ ( .D(n4374), .CLK(n4154), .Q(n_T_427[596]) );
  DFFX1_LVT u_T_427_reg_21__19_ ( .D(n4371), .CLK(n4154), .Q(n_T_427[595]) );
  DFFX1_LVT u_T_427_reg_21__18_ ( .D(n4368), .CLK(n4154), .Q(n_T_427[594]) );
  DFFX1_LVT u_T_427_reg_21__17_ ( .D(n4366), .CLK(n4154), .Q(n_T_427[593]) );
  DFFX1_LVT u_T_427_reg_21__16_ ( .D(n4363), .CLK(n4154), .Q(n_T_427[592]) );
  DFFX1_LVT u_T_427_reg_21__15_ ( .D(n4360), .CLK(n4154), .Q(n_T_427[591]) );
  DFFX1_LVT u_T_427_reg_21__14_ ( .D(n4358), .CLK(n4154), .Q(n_T_427[590]) );
  DFFX1_LVT u_T_427_reg_21__13_ ( .D(n4355), .CLK(n4154), .Q(n_T_427[589]) );
  DFFX1_LVT u_T_427_reg_21__12_ ( .D(n4353), .CLK(n4154), .Q(n_T_427[588]) );
  DFFX1_LVT u_T_427_reg_21__11_ ( .D(n4349), .CLK(n4153), .Q(n_T_427[587]) );
  DFFX1_LVT u_T_427_reg_21__10_ ( .D(n4347), .CLK(n4153), .Q(n_T_427[586]) );
  DFFX1_LVT u_T_427_reg_21__9_ ( .D(n4344), .CLK(n4153), .Q(n_T_427[585]) );
  DFFX1_LVT u_T_427_reg_21__8_ ( .D(n4341), .CLK(n4153), .Q(n_T_427[584]) );
  DFFX1_LVT u_T_427_reg_21__7_ ( .D(n4338), .CLK(n4153), .Q(n_T_427[583]) );
  DFFX1_LVT u_T_427_reg_21__6_ ( .D(n4335), .CLK(n4153), .Q(n_T_427[582]) );
  DFFX1_LVT u_T_427_reg_21__5_ ( .D(n4332), .CLK(n4153), .Q(n_T_427[581]) );
  DFFX1_LVT u_T_427_reg_21__4_ ( .D(n4329), .CLK(n4153), .Q(n_T_427[580]) );
  DFFX1_LVT u_T_427_reg_21__3_ ( .D(n4326), .CLK(n4153), .Q(n_T_427[579]) );
  DFFX1_LVT u_T_427_reg_21__2_ ( .D(n4323), .CLK(n4153), .Q(n_T_427[578]) );
  DFFX1_LVT u_T_427_reg_21__1_ ( .D(n4319), .CLK(n4153), .Q(n_T_427[577]) );
  DFFX1_LVT u_T_427_reg_21__0_ ( .D(n4316), .CLK(n4153), .Q(n_T_427[576]) );
  DFFX1_LVT u_T_427_reg_22__63_ ( .D(n4495), .CLK(n4152), .Q(n_T_427[575]) );
  DFFX1_LVT u_T_427_reg_22__62_ ( .D(n4492), .CLK(n4152), .Q(n_T_427[574]) );
  DFFX1_LVT u_T_427_reg_22__61_ ( .D(n4489), .CLK(n4152), .Q(n_T_427[573]) );
  DFFX1_LVT u_T_427_reg_22__60_ ( .D(n4486), .CLK(n4152), .Q(n_T_427[572]) );
  DFFX1_LVT u_T_427_reg_22__59_ ( .D(n4483), .CLK(n4151), .Q(n_T_427[571]) );
  DFFX1_LVT u_T_427_reg_22__58_ ( .D(n4479), .CLK(n4151), .Q(n_T_427[570]) );
  DFFX1_LVT u_T_427_reg_22__57_ ( .D(n4477), .CLK(n4151), .Q(n_T_427[569]) );
  DFFX1_LVT u_T_427_reg_22__56_ ( .D(n4473), .CLK(n4151), .Q(n_T_427[568]) );
  DFFX1_LVT u_T_427_reg_22__55_ ( .D(n4471), .CLK(n4151), .Q(n_T_427[567]) );
  DFFX1_LVT u_T_427_reg_22__54_ ( .D(n4467), .CLK(n4151), .Q(n_T_427[566]) );
  DFFX1_LVT u_T_427_reg_22__53_ ( .D(n4465), .CLK(n4151), .Q(n_T_427[565]) );
  DFFX1_LVT u_T_427_reg_22__52_ ( .D(n4461), .CLK(n4151), .Q(n_T_427[564]) );
  DFFX1_LVT u_T_427_reg_22__51_ ( .D(n4458), .CLK(n4151), .Q(n_T_427[563]) );
  DFFX1_LVT u_T_427_reg_22__50_ ( .D(n4456), .CLK(n4151), .Q(n_T_427[562]) );
  DFFX1_LVT u_T_427_reg_22__49_ ( .D(n4452), .CLK(n4151), .Q(n_T_427[561]) );
  DFFX1_LVT u_T_427_reg_22__48_ ( .D(n4450), .CLK(n4151), .Q(n_T_427[560]) );
  DFFX1_LVT u_T_427_reg_22__47_ ( .D(n4447), .CLK(n4150), .Q(n_T_427[559]) );
  DFFX1_LVT u_T_427_reg_22__46_ ( .D(n4444), .CLK(n4150), .Q(n_T_427[558]) );
  DFFX1_LVT u_T_427_reg_22__45_ ( .D(n4440), .CLK(n4150), .Q(n_T_427[557]) );
  DFFX1_LVT u_T_427_reg_22__44_ ( .D(n4438), .CLK(n4150), .Q(n_T_427[556]) );
  DFFX1_LVT u_T_427_reg_22__43_ ( .D(n4434), .CLK(n4150), .Q(n_T_427[555]) );
  DFFX1_LVT u_T_427_reg_22__42_ ( .D(n4431), .CLK(n4150), .Q(n_T_427[554]) );
  DFFX1_LVT u_T_427_reg_22__41_ ( .D(n4428), .CLK(n4150), .Q(n_T_427[553]) );
  DFFX1_LVT u_T_427_reg_22__40_ ( .D(n4426), .CLK(n4150), .Q(n_T_427[552]) );
  DFFX1_LVT u_T_427_reg_22__39_ ( .D(n4423), .CLK(n4150), .Q(n_T_427[551]) );
  DFFX1_LVT u_T_427_reg_22__38_ ( .D(n4420), .CLK(n4150), .Q(n_T_427[550]) );
  DFFX1_LVT u_T_427_reg_22__37_ ( .D(n4418), .CLK(n4150), .Q(n_T_427[549]) );
  DFFX1_LVT u_T_427_reg_22__36_ ( .D(n4414), .CLK(n4150), .Q(n_T_427[548]) );
  DFFX1_LVT u_T_427_reg_22__35_ ( .D(n4412), .CLK(n4149), .Q(n_T_427[547]) );
  DFFX1_LVT u_T_427_reg_22__34_ ( .D(n4410), .CLK(n4149), .Q(n_T_427[546]) );
  DFFX1_LVT u_T_427_reg_22__33_ ( .D(n4407), .CLK(n4149), .Q(n_T_427[545]) );
  DFFX1_LVT u_T_427_reg_22__32_ ( .D(n4405), .CLK(n4149), .Q(n_T_427[544]) );
  DFFX1_LVT u_T_427_reg_22__31_ ( .D(n4402), .CLK(n4149), .Q(n_T_427[543]) );
  DFFX1_LVT u_T_427_reg_22__30_ ( .D(n4399), .CLK(n4149), .Q(n_T_427[542]) );
  DFFX1_LVT u_T_427_reg_22__29_ ( .D(n4396), .CLK(n4149), .Q(n_T_427[541]) );
  DFFX1_LVT u_T_427_reg_22__28_ ( .D(n4394), .CLK(n4149), .Q(n_T_427[540]) );
  DFFX1_LVT u_T_427_reg_22__27_ ( .D(n4392), .CLK(n4149), .Q(n_T_427[539]) );
  DFFX1_LVT u_T_427_reg_22__26_ ( .D(n4389), .CLK(n4149), .Q(n_T_427[538]) );
  DFFX1_LVT u_T_427_reg_22__25_ ( .D(n4387), .CLK(n4149), .Q(n_T_427[537]) );
  DFFX1_LVT u_T_427_reg_22__24_ ( .D(n4384), .CLK(n4149), .Q(n_T_427[536]) );
  DFFX1_LVT u_T_427_reg_22__23_ ( .D(n4382), .CLK(n4148), .Q(n_T_427[535]) );
  DFFX1_LVT u_T_427_reg_22__22_ ( .D(n4379), .CLK(n4148), .Q(n_T_427[534]) );
  DFFX1_LVT u_T_427_reg_22__21_ ( .D(n4377), .CLK(n4148), .Q(n_T_427[533]) );
  DFFX1_LVT u_T_427_reg_22__20_ ( .D(n4374), .CLK(n4148), .Q(n_T_427[532]) );
  DFFX1_LVT u_T_427_reg_22__19_ ( .D(n4371), .CLK(n4148), .Q(n_T_427[531]) );
  DFFX1_LVT u_T_427_reg_22__18_ ( .D(n4368), .CLK(n4148), .Q(n_T_427[530]) );
  DFFX1_LVT u_T_427_reg_22__17_ ( .D(n4366), .CLK(n4148), .Q(n_T_427[529]) );
  DFFX1_LVT u_T_427_reg_22__16_ ( .D(n4363), .CLK(n4148), .Q(n_T_427[528]) );
  DFFX1_LVT u_T_427_reg_22__15_ ( .D(n4360), .CLK(n4148), .Q(n_T_427[527]) );
  DFFX1_LVT u_T_427_reg_22__14_ ( .D(n4358), .CLK(n4148), .Q(n_T_427[526]) );
  DFFX1_LVT u_T_427_reg_22__13_ ( .D(n4355), .CLK(n4148), .Q(n_T_427[525]) );
  DFFX1_LVT u_T_427_reg_22__12_ ( .D(n4353), .CLK(n4148), .Q(n_T_427[524]) );
  DFFX1_LVT u_T_427_reg_22__11_ ( .D(n4349), .CLK(n4147), .Q(n_T_427[523]) );
  DFFX1_LVT u_T_427_reg_22__10_ ( .D(n4347), .CLK(n4147), .Q(n_T_427[522]) );
  DFFX1_LVT u_T_427_reg_22__9_ ( .D(n4344), .CLK(n4147), .Q(n_T_427[521]) );
  DFFX1_LVT u_T_427_reg_22__8_ ( .D(n4341), .CLK(n4147), .Q(n_T_427[520]) );
  DFFX1_LVT u_T_427_reg_22__7_ ( .D(n4338), .CLK(n4147), .Q(n_T_427[519]) );
  DFFX1_LVT u_T_427_reg_22__6_ ( .D(n4335), .CLK(n4147), .Q(n_T_427[518]) );
  DFFX1_LVT u_T_427_reg_22__5_ ( .D(n4332), .CLK(n4147), .Q(n_T_427[517]) );
  DFFX1_LVT u_T_427_reg_22__4_ ( .D(n4329), .CLK(n4147), .Q(n_T_427[516]) );
  DFFX1_LVT u_T_427_reg_22__3_ ( .D(n4326), .CLK(n4147), .Q(n_T_427[515]) );
  DFFX1_LVT u_T_427_reg_22__2_ ( .D(n4323), .CLK(n4147), .Q(n_T_427[514]) );
  DFFX1_LVT u_T_427_reg_22__1_ ( .D(n4319), .CLK(n4147), .Q(n_T_427[513]) );
  DFFX1_LVT u_T_427_reg_22__0_ ( .D(n4316), .CLK(n4147), .Q(n_T_427[512]) );
  DFFX1_LVT u_T_427_reg_23__63_ ( .D(n4495), .CLK(n4146), .Q(n_T_427[511]) );
  DFFX1_LVT u_T_427_reg_23__62_ ( .D(n4492), .CLK(n4146), .Q(n_T_427[510]) );
  DFFX1_LVT u_T_427_reg_23__61_ ( .D(n4489), .CLK(n4146), .Q(n_T_427[509]) );
  DFFX1_LVT u_T_427_reg_23__60_ ( .D(n4486), .CLK(n4146), .Q(n_T_427[508]) );
  DFFX1_LVT u_T_427_reg_23__59_ ( .D(n4483), .CLK(n4145), .Q(n_T_427[507]) );
  DFFX1_LVT u_T_427_reg_23__58_ ( .D(n4479), .CLK(n4145), .Q(n_T_427[506]) );
  DFFX1_LVT u_T_427_reg_23__57_ ( .D(n4477), .CLK(n4145), .Q(n_T_427[505]) );
  DFFX1_LVT u_T_427_reg_23__56_ ( .D(n4473), .CLK(n4145), .Q(n_T_427[504]) );
  DFFX1_LVT u_T_427_reg_23__55_ ( .D(n4471), .CLK(n4145), .Q(n_T_427[503]) );
  DFFX1_LVT u_T_427_reg_23__54_ ( .D(n4467), .CLK(n4145), .Q(n_T_427[502]) );
  DFFX1_LVT u_T_427_reg_23__53_ ( .D(n4465), .CLK(n4145), .Q(n_T_427[501]) );
  DFFX1_LVT u_T_427_reg_23__52_ ( .D(n4461), .CLK(n4145), .Q(n_T_427[500]) );
  DFFX1_LVT u_T_427_reg_23__51_ ( .D(n4458), .CLK(n4145), .Q(n_T_427[499]) );
  DFFX1_LVT u_T_427_reg_23__50_ ( .D(n4456), .CLK(n4145), .Q(n_T_427[498]) );
  DFFX1_LVT u_T_427_reg_23__49_ ( .D(n4452), .CLK(n4145), .Q(n_T_427[497]) );
  DFFX1_LVT u_T_427_reg_23__48_ ( .D(n4450), .CLK(n4145), .Q(n_T_427[496]) );
  DFFX1_LVT u_T_427_reg_23__47_ ( .D(n4447), .CLK(n4144), .Q(n_T_427[495]) );
  DFFX1_LVT u_T_427_reg_23__46_ ( .D(n4444), .CLK(n4144), .Q(n_T_427[494]) );
  DFFX1_LVT u_T_427_reg_23__45_ ( .D(n4440), .CLK(n4144), .Q(n_T_427[493]) );
  DFFX1_LVT u_T_427_reg_23__44_ ( .D(n4438), .CLK(n4144), .Q(n_T_427[492]) );
  DFFX1_LVT u_T_427_reg_23__43_ ( .D(n4434), .CLK(n4144), .Q(n_T_427[491]) );
  DFFX1_LVT u_T_427_reg_23__42_ ( .D(n4431), .CLK(n4144), .Q(n_T_427[490]) );
  DFFX1_LVT u_T_427_reg_23__41_ ( .D(n4428), .CLK(n4144), .Q(n_T_427[489]) );
  DFFX1_LVT u_T_427_reg_23__40_ ( .D(n4426), .CLK(n4144), .Q(n_T_427[488]) );
  DFFX1_LVT u_T_427_reg_23__39_ ( .D(n4423), .CLK(n4144), .Q(n_T_427[487]) );
  DFFX1_LVT u_T_427_reg_23__38_ ( .D(n4420), .CLK(n4144), .Q(n_T_427[486]) );
  DFFX1_LVT u_T_427_reg_23__37_ ( .D(n4418), .CLK(n4144), .Q(n_T_427[485]) );
  DFFX1_LVT u_T_427_reg_23__36_ ( .D(n4414), .CLK(n4144), .Q(n_T_427[484]) );
  DFFX1_LVT u_T_427_reg_23__35_ ( .D(n4412), .CLK(n4143), .Q(n_T_427[483]) );
  DFFX1_LVT u_T_427_reg_23__34_ ( .D(n4410), .CLK(n4143), .Q(n_T_427[482]) );
  DFFX1_LVT u_T_427_reg_23__33_ ( .D(n4407), .CLK(n4143), .Q(n_T_427[481]) );
  DFFX1_LVT u_T_427_reg_23__32_ ( .D(n4405), .CLK(n4143), .Q(n_T_427[480]) );
  DFFX1_LVT u_T_427_reg_23__31_ ( .D(n4402), .CLK(n4143), .Q(n_T_427[479]) );
  DFFX1_LVT u_T_427_reg_23__30_ ( .D(n4399), .CLK(n4143), .Q(n_T_427[478]) );
  DFFX1_LVT u_T_427_reg_23__29_ ( .D(n4396), .CLK(n4143), .Q(n_T_427[477]) );
  DFFX1_LVT u_T_427_reg_23__28_ ( .D(n4394), .CLK(n4143), .Q(n_T_427[476]) );
  DFFX1_LVT u_T_427_reg_23__27_ ( .D(n4392), .CLK(n4143), .Q(n_T_427[475]) );
  DFFX1_LVT u_T_427_reg_23__26_ ( .D(n4389), .CLK(n4143), .Q(n_T_427[474]) );
  DFFX1_LVT u_T_427_reg_23__25_ ( .D(n4387), .CLK(n4143), .Q(n_T_427[473]) );
  DFFX1_LVT u_T_427_reg_23__24_ ( .D(n4384), .CLK(n4143), .Q(n_T_427[472]) );
  DFFX1_LVT u_T_427_reg_23__23_ ( .D(n4382), .CLK(n4142), .Q(n_T_427[471]) );
  DFFX1_LVT u_T_427_reg_23__22_ ( .D(n4379), .CLK(n4142), .Q(n_T_427[470]) );
  DFFX1_LVT u_T_427_reg_23__21_ ( .D(n4377), .CLK(n4142), .Q(n_T_427[469]) );
  DFFX1_LVT u_T_427_reg_23__20_ ( .D(n4374), .CLK(n4142), .Q(n_T_427[468]) );
  DFFX1_LVT u_T_427_reg_23__19_ ( .D(n4371), .CLK(n4142), .Q(n_T_427[467]) );
  DFFX1_LVT u_T_427_reg_23__18_ ( .D(n4368), .CLK(n4142), .Q(n_T_427[466]) );
  DFFX1_LVT u_T_427_reg_23__17_ ( .D(n4366), .CLK(n4142), .Q(n_T_427[465]) );
  DFFX1_LVT u_T_427_reg_23__16_ ( .D(n4363), .CLK(n4142), .Q(n_T_427[464]) );
  DFFX1_LVT u_T_427_reg_23__15_ ( .D(n4360), .CLK(n4142), .Q(n_T_427[463]) );
  DFFX1_LVT u_T_427_reg_23__14_ ( .D(n4358), .CLK(n4142), .Q(n_T_427[462]) );
  DFFX1_LVT u_T_427_reg_23__13_ ( .D(n4355), .CLK(n4142), .Q(n_T_427[461]) );
  DFFX1_LVT u_T_427_reg_23__12_ ( .D(n4353), .CLK(n4142), .Q(n_T_427[460]) );
  DFFX1_LVT u_T_427_reg_23__11_ ( .D(n4349), .CLK(n4141), .Q(n_T_427[459]) );
  DFFX1_LVT u_T_427_reg_23__10_ ( .D(n4347), .CLK(n4141), .Q(n_T_427[458]) );
  DFFX1_LVT u_T_427_reg_23__9_ ( .D(n4344), .CLK(n4141), .Q(n_T_427[457]) );
  DFFX1_LVT u_T_427_reg_23__8_ ( .D(n4341), .CLK(n4141), .Q(n_T_427[456]) );
  DFFX1_LVT u_T_427_reg_23__7_ ( .D(n4338), .CLK(n4141), .Q(n_T_427[455]) );
  DFFX1_LVT u_T_427_reg_23__6_ ( .D(n4335), .CLK(n4141), .Q(n_T_427[454]) );
  DFFX1_LVT u_T_427_reg_23__5_ ( .D(n4332), .CLK(n4141), .Q(n_T_427[453]) );
  DFFX1_LVT u_T_427_reg_23__4_ ( .D(n4329), .CLK(n4141), .Q(n_T_427[452]) );
  DFFX1_LVT u_T_427_reg_23__3_ ( .D(n4326), .CLK(n4141), .Q(n_T_427[451]) );
  DFFX1_LVT u_T_427_reg_23__2_ ( .D(n4323), .CLK(n4141), .Q(n_T_427[450]) );
  DFFX1_LVT u_T_427_reg_23__1_ ( .D(n4319), .CLK(n4141), .Q(n_T_427[449]) );
  DFFX1_LVT u_T_427_reg_23__0_ ( .D(n4316), .CLK(n4141), .Q(n_T_427[448]) );
  DFFX1_LVT u_T_427_reg_24__63_ ( .D(n4496), .CLK(n4140), .Q(n_T_427[447]) );
  DFFX1_LVT u_T_427_reg_24__62_ ( .D(n4493), .CLK(n4140), .Q(n_T_427[446]) );
  DFFX1_LVT u_T_427_reg_24__61_ ( .D(n4490), .CLK(n4140), .Q(n_T_427[445]) );
  DFFX1_LVT u_T_427_reg_24__60_ ( .D(n4487), .CLK(n4140), .Q(n_T_427[444]), 
        .QN(n3525) );
  DFFX1_LVT u_T_427_reg_24__59_ ( .D(n4484), .CLK(n4139), .Q(n_T_427[443]) );
  DFFX1_LVT u_T_427_reg_24__58_ ( .D(n4480), .CLK(n4139), .Q(n_T_427[442]) );
  DFFX1_LVT u_T_427_reg_24__57_ ( .D(n4478), .CLK(n4139), .Q(n_T_427[441]) );
  DFFX1_LVT u_T_427_reg_24__56_ ( .D(n4474), .CLK(n4139), .Q(n_T_427[440]) );
  DFFX1_LVT u_T_427_reg_24__55_ ( .D(n4472), .CLK(n4139), .Q(n_T_427[439]) );
  DFFX1_LVT u_T_427_reg_24__54_ ( .D(n4468), .CLK(n4139), .Q(n_T_427[438]) );
  DFFX1_LVT u_T_427_reg_24__53_ ( .D(n4466), .CLK(n4139), .Q(n_T_427[437]) );
  DFFX1_LVT u_T_427_reg_24__52_ ( .D(n4462), .CLK(n4139), .Q(n_T_427[436]) );
  DFFX1_LVT u_T_427_reg_24__51_ ( .D(n4459), .CLK(n4139), .Q(n_T_427[435]) );
  DFFX1_LVT u_T_427_reg_24__50_ ( .D(n4457), .CLK(n4139), .Q(n_T_427[434]) );
  DFFX1_LVT u_T_427_reg_24__49_ ( .D(n4453), .CLK(n4139), .Q(n_T_427[433]) );
  DFFX1_LVT u_T_427_reg_24__48_ ( .D(n4451), .CLK(n4139), .Q(n_T_427[432]) );
  DFFX1_LVT u_T_427_reg_24__47_ ( .D(n4448), .CLK(n4138), .Q(n_T_427[431]) );
  DFFX1_LVT u_T_427_reg_24__46_ ( .D(n4445), .CLK(n4138), .Q(n_T_427[430]) );
  DFFX1_LVT u_T_427_reg_24__45_ ( .D(n4441), .CLK(n4138), .Q(n_T_427[429]) );
  DFFX1_LVT u_T_427_reg_24__44_ ( .D(n4439), .CLK(n4138), .Q(n_T_427[428]) );
  DFFX1_LVT u_T_427_reg_24__43_ ( .D(n4435), .CLK(n4138), .Q(n_T_427[427]) );
  DFFX1_LVT u_T_427_reg_24__42_ ( .D(n4432), .CLK(n4138), .Q(n_T_427[426]) );
  DFFX1_LVT u_T_427_reg_24__41_ ( .D(n4429), .CLK(n4138), .Q(n_T_427[425]) );
  DFFX1_LVT u_T_427_reg_24__40_ ( .D(n4427), .CLK(n4138), .Q(n_T_427[424]) );
  DFFX1_LVT u_T_427_reg_24__39_ ( .D(n4424), .CLK(n4138), .Q(n_T_427[423]) );
  DFFX1_LVT u_T_427_reg_24__38_ ( .D(n4421), .CLK(n4138), .Q(n_T_427[422]) );
  DFFX1_LVT u_T_427_reg_24__37_ ( .D(n4419), .CLK(n4138), .Q(n_T_427[421]) );
  DFFX1_LVT u_T_427_reg_24__36_ ( .D(n4415), .CLK(n4138), .Q(n_T_427[420]) );
  DFFX1_LVT u_T_427_reg_24__35_ ( .D(n4413), .CLK(n4137), .Q(n_T_427[419]) );
  DFFX1_LVT u_T_427_reg_24__34_ ( .D(n4411), .CLK(n4137), .Q(n_T_427[418]), 
        .QN(n3527) );
  DFFX1_LVT u_T_427_reg_24__33_ ( .D(n4408), .CLK(n4137), .Q(n_T_427[417]) );
  DFFX1_LVT u_T_427_reg_24__32_ ( .D(n4406), .CLK(n4137), .Q(n_T_427[416]) );
  DFFX1_LVT u_T_427_reg_24__31_ ( .D(n4403), .CLK(n4137), .Q(n_T_427[415]) );
  DFFX1_LVT u_T_427_reg_24__30_ ( .D(n4400), .CLK(n4137), .Q(n_T_427[414]) );
  DFFX1_LVT u_T_427_reg_24__29_ ( .D(n4397), .CLK(n4137), .Q(n_T_427[413]) );
  DFFX1_LVT u_T_427_reg_24__28_ ( .D(n4395), .CLK(n4137), .Q(n_T_427[412]) );
  DFFX1_LVT u_T_427_reg_24__27_ ( .D(n4393), .CLK(n4137), .Q(n_T_427[411]) );
  DFFX1_LVT u_T_427_reg_24__26_ ( .D(n4390), .CLK(n4137), .Q(n_T_427[410]) );
  DFFX1_LVT u_T_427_reg_24__25_ ( .D(n4388), .CLK(n4137), .Q(n_T_427[409]) );
  DFFX1_LVT u_T_427_reg_24__24_ ( .D(n4385), .CLK(n4137), .Q(n_T_427[408]) );
  DFFX1_LVT u_T_427_reg_24__23_ ( .D(n4383), .CLK(n4136), .Q(n_T_427[407]) );
  DFFX1_LVT u_T_427_reg_24__22_ ( .D(n4380), .CLK(n4136), .Q(n_T_427[406]) );
  DFFX1_LVT u_T_427_reg_24__21_ ( .D(n4378), .CLK(n4136), .Q(n_T_427[405]) );
  DFFX1_LVT u_T_427_reg_24__20_ ( .D(n4375), .CLK(n4136), .Q(n_T_427[404]) );
  DFFX1_LVT u_T_427_reg_24__19_ ( .D(n4372), .CLK(n4136), .Q(n_T_427[403]) );
  DFFX1_LVT u_T_427_reg_24__18_ ( .D(n4369), .CLK(n4136), .Q(n_T_427[402]) );
  DFFX1_LVT u_T_427_reg_24__17_ ( .D(n4367), .CLK(n4136), .Q(n_T_427[401]) );
  DFFX1_LVT u_T_427_reg_24__16_ ( .D(n4364), .CLK(n4136), .Q(n_T_427[400]) );
  DFFX1_LVT u_T_427_reg_24__15_ ( .D(n4361), .CLK(n4136), .Q(n_T_427[399]) );
  DFFX1_LVT u_T_427_reg_24__14_ ( .D(n4359), .CLK(n4136), .Q(n_T_427[398]) );
  DFFX1_LVT u_T_427_reg_24__13_ ( .D(n4356), .CLK(n4136), .Q(n_T_427[397]) );
  DFFX1_LVT u_T_427_reg_24__12_ ( .D(n4354), .CLK(n4136), .Q(n_T_427[396]) );
  DFFX1_LVT u_T_427_reg_24__11_ ( .D(n4349), .CLK(n4135), .Q(n_T_427[395]) );
  DFFX1_LVT u_T_427_reg_24__10_ ( .D(n4348), .CLK(n4135), .Q(n_T_427[394]) );
  DFFX1_LVT u_T_427_reg_24__9_ ( .D(n4345), .CLK(n4135), .Q(n_T_427[393]) );
  DFFX1_LVT u_T_427_reg_24__8_ ( .D(n4342), .CLK(n4135), .Q(n_T_427[392]) );
  DFFX1_LVT u_T_427_reg_24__7_ ( .D(n4339), .CLK(n4135), .Q(n_T_427[391]) );
  DFFX1_LVT u_T_427_reg_24__6_ ( .D(n4336), .CLK(n4135), .Q(n_T_427[390]) );
  DFFX1_LVT u_T_427_reg_24__5_ ( .D(n4333), .CLK(n4135), .Q(n_T_427[389]) );
  DFFX1_LVT u_T_427_reg_24__4_ ( .D(n4330), .CLK(n4135), .Q(n_T_427[388]) );
  DFFX1_LVT u_T_427_reg_24__3_ ( .D(n4327), .CLK(n4135), .Q(n_T_427[387]) );
  DFFX1_LVT u_T_427_reg_24__2_ ( .D(n4324), .CLK(n4135), .Q(n_T_427[386]) );
  DFFX1_LVT u_T_427_reg_24__1_ ( .D(n4320), .CLK(n4135), .Q(n_T_427[385]) );
  DFFX1_LVT u_T_427_reg_24__0_ ( .D(n4317), .CLK(n4135), .Q(n_T_427[384]) );
  DFFX1_LVT u_T_427_reg_25__63_ ( .D(n4496), .CLK(n4134), .Q(n_T_427[383]) );
  DFFX1_LVT u_T_427_reg_25__62_ ( .D(n4493), .CLK(n4134), .Q(n_T_427[382]) );
  DFFX1_LVT u_T_427_reg_25__61_ ( .D(n4490), .CLK(n4134), .Q(n_T_427[381]) );
  DFFX1_LVT u_T_427_reg_25__60_ ( .D(n4487), .CLK(n4134), .Q(n_T_427[380]), 
        .QN(n3172) );
  DFFX1_LVT u_T_427_reg_25__59_ ( .D(n4484), .CLK(n4133), .Q(n_T_427[379]) );
  DFFX1_LVT u_T_427_reg_25__58_ ( .D(n4479), .CLK(n4133), .Q(n_T_427[378]) );
  DFFX1_LVT u_T_427_reg_25__57_ ( .D(n4478), .CLK(n4133), .Q(n_T_427[377]) );
  DFFX1_LVT u_T_427_reg_25__56_ ( .D(n4473), .CLK(n4133), .Q(n_T_427[376]) );
  DFFX1_LVT u_T_427_reg_25__55_ ( .D(n4472), .CLK(n4133), .Q(n_T_427[375]) );
  DFFX1_LVT u_T_427_reg_25__54_ ( .D(n4467), .CLK(n4133), .Q(n_T_427[374]) );
  DFFX1_LVT u_T_427_reg_25__53_ ( .D(n4466), .CLK(n4133), .Q(n_T_427[373]) );
  DFFX1_LVT u_T_427_reg_25__52_ ( .D(n4461), .CLK(n4133), .Q(n_T_427[372]) );
  DFFX1_LVT u_T_427_reg_25__51_ ( .D(n4458), .CLK(n4133), .Q(n_T_427[371]) );
  DFFX1_LVT u_T_427_reg_25__50_ ( .D(n4457), .CLK(n4133), .Q(n_T_427[370]) );
  DFFX1_LVT u_T_427_reg_25__49_ ( .D(n4452), .CLK(n4133), .Q(n_T_427[369]) );
  DFFX1_LVT u_T_427_reg_25__48_ ( .D(n4451), .CLK(n4133), .Q(n_T_427[368]) );
  DFFX1_LVT u_T_427_reg_25__47_ ( .D(n4448), .CLK(n4132), .Q(n_T_427[367]) );
  DFFX1_LVT u_T_427_reg_25__46_ ( .D(n4445), .CLK(n4132), .Q(n_T_427[366]) );
  DFFX1_LVT u_T_427_reg_25__45_ ( .D(n4440), .CLK(n4132), .Q(n_T_427[365]) );
  DFFX1_LVT u_T_427_reg_25__44_ ( .D(n4439), .CLK(n4132), .Q(n_T_427[364]) );
  DFFX1_LVT u_T_427_reg_25__43_ ( .D(n4434), .CLK(n4132), .Q(n_T_427[363]) );
  DFFX1_LVT u_T_427_reg_25__42_ ( .D(n4431), .CLK(n4132), .Q(n_T_427[362]) );
  DFFX1_LVT u_T_427_reg_25__41_ ( .D(n4428), .CLK(n4132), .Q(n_T_427[361]) );
  DFFX1_LVT u_T_427_reg_25__40_ ( .D(n4427), .CLK(n4132), .Q(n_T_427[360]) );
  DFFX1_LVT u_T_427_reg_25__39_ ( .D(n4424), .CLK(n4132), .Q(n_T_427[359]) );
  DFFX1_LVT u_T_427_reg_25__38_ ( .D(n4421), .CLK(n4132), .Q(n_T_427[358]) );
  DFFX1_LVT u_T_427_reg_25__37_ ( .D(n4419), .CLK(n4132), .Q(n_T_427[357]) );
  DFFX1_LVT u_T_427_reg_25__36_ ( .D(n4414), .CLK(n4132), .Q(n_T_427[356]) );
  DFFX1_LVT u_T_427_reg_25__35_ ( .D(n4413), .CLK(n4131), .Q(n_T_427[355]) );
  DFFX1_LVT u_T_427_reg_25__34_ ( .D(n4411), .CLK(n4131), .Q(n_T_427[354]) );
  DFFX1_LVT u_T_427_reg_25__33_ ( .D(n4408), .CLK(n4131), .Q(n_T_427[353]) );
  DFFX1_LVT u_T_427_reg_25__32_ ( .D(n4406), .CLK(n4131), .Q(n_T_427[352]) );
  DFFX1_LVT u_T_427_reg_25__31_ ( .D(n4403), .CLK(n4131), .Q(n_T_427[351]) );
  DFFX1_LVT u_T_427_reg_25__30_ ( .D(n4399), .CLK(n4131), .Q(n_T_427[350]) );
  DFFX1_LVT u_T_427_reg_25__29_ ( .D(n4396), .CLK(n4131), .Q(n_T_427[349]) );
  DFFX1_LVT u_T_427_reg_25__28_ ( .D(n4395), .CLK(n4131), .Q(n_T_427[348]) );
  DFFX1_LVT u_T_427_reg_25__27_ ( .D(n4393), .CLK(n4131), .Q(n_T_427[347]) );
  DFFX1_LVT u_T_427_reg_25__26_ ( .D(n4390), .CLK(n4131), .Q(n_T_427[346]) );
  DFFX1_LVT u_T_427_reg_25__25_ ( .D(n4388), .CLK(n4131), .Q(n_T_427[345]) );
  DFFX1_LVT u_T_427_reg_25__24_ ( .D(n4384), .CLK(n4131), .Q(n_T_427[344]) );
  DFFX1_LVT u_T_427_reg_25__23_ ( .D(n4383), .CLK(n4130), .Q(n_T_427[343]) );
  DFFX1_LVT u_T_427_reg_25__22_ ( .D(n4380), .CLK(n4130), .Q(n_T_427[342]) );
  DFFX1_LVT u_T_427_reg_25__21_ ( .D(n4378), .CLK(n4130), .Q(n_T_427[341]) );
  DFFX1_LVT u_T_427_reg_25__20_ ( .D(n4374), .CLK(n4130), .Q(n_T_427[340]) );
  DFFX1_LVT u_T_427_reg_25__19_ ( .D(n4371), .CLK(n4130), .Q(n_T_427[339]) );
  DFFX1_LVT u_T_427_reg_25__18_ ( .D(n4368), .CLK(n4130), .Q(n_T_427[338]) );
  DFFX1_LVT u_T_427_reg_25__17_ ( .D(n4367), .CLK(n4130), .Q(n_T_427[337]) );
  DFFX1_LVT u_T_427_reg_25__16_ ( .D(n4364), .CLK(n4130), .Q(n_T_427[336]) );
  DFFX1_LVT u_T_427_reg_25__15_ ( .D(n4361), .CLK(n4130), .Q(n_T_427[335]) );
  DFFX1_LVT u_T_427_reg_25__14_ ( .D(n4359), .CLK(n4130), .Q(n_T_427[334]) );
  DFFX1_LVT u_T_427_reg_25__13_ ( .D(n4356), .CLK(n4130), .Q(n_T_427[333]) );
  DFFX1_LVT u_T_427_reg_25__12_ ( .D(n4354), .CLK(n4130), .Q(n_T_427[332]) );
  DFFX1_LVT u_T_427_reg_25__11_ ( .D(n4349), .CLK(n4129), .Q(n_T_427[331]) );
  DFFX1_LVT u_T_427_reg_25__10_ ( .D(n4348), .CLK(n4129), .Q(n_T_427[330]) );
  DFFX1_LVT u_T_427_reg_25__9_ ( .D(n4345), .CLK(n4129), .Q(n_T_427[329]) );
  DFFX1_LVT u_T_427_reg_25__8_ ( .D(n4342), .CLK(n4129), .Q(n_T_427[328]) );
  DFFX1_LVT u_T_427_reg_25__7_ ( .D(n4339), .CLK(n4129), .Q(n_T_427[327]) );
  DFFX1_LVT u_T_427_reg_25__6_ ( .D(n4336), .CLK(n4129), .Q(n_T_427[326]) );
  DFFX1_LVT u_T_427_reg_25__5_ ( .D(n4333), .CLK(n4129), .Q(n_T_427[325]) );
  DFFX1_LVT u_T_427_reg_25__4_ ( .D(n4330), .CLK(n4129), .Q(n_T_427[324]), 
        .QN(n3520) );
  DFFX1_LVT u_T_427_reg_25__3_ ( .D(n4327), .CLK(n4129), .Q(n_T_427[323]) );
  DFFX1_LVT u_T_427_reg_25__2_ ( .D(n4324), .CLK(n4129), .Q(n_T_427[322]), 
        .QN(n3519) );
  DFFX1_LVT u_T_427_reg_25__1_ ( .D(n4319), .CLK(n4129), .Q(n_T_427[321]) );
  DFFX1_LVT u_T_427_reg_25__0_ ( .D(n4316), .CLK(n4129), .Q(n_T_427[320]) );
  DFFX1_LVT u_T_427_reg_26__63_ ( .D(n4496), .CLK(n4128), .Q(n_T_427[319]) );
  DFFX1_LVT u_T_427_reg_26__62_ ( .D(n4493), .CLK(n4128), .Q(n_T_427[318]) );
  DFFX1_LVT u_T_427_reg_26__61_ ( .D(n4490), .CLK(n4128), .Q(n_T_427[317]) );
  DFFX1_LVT u_T_427_reg_26__60_ ( .D(n4487), .CLK(n4128), .Q(n_T_427[316]) );
  DFFX1_LVT u_T_427_reg_26__59_ ( .D(n4484), .CLK(n4127), .Q(n_T_427[315]) );
  DFFX1_LVT u_T_427_reg_26__58_ ( .D(n4479), .CLK(n4127), .Q(n_T_427[314]) );
  DFFX1_LVT u_T_427_reg_26__57_ ( .D(n4478), .CLK(n4127), .Q(n_T_427[313]) );
  DFFX1_LVT u_T_427_reg_26__56_ ( .D(n4473), .CLK(n4127), .Q(n_T_427[312]) );
  DFFX1_LVT u_T_427_reg_26__55_ ( .D(n4472), .CLK(n4127), .Q(n_T_427[311]) );
  DFFX1_LVT u_T_427_reg_26__54_ ( .D(n4467), .CLK(n4127), .Q(n_T_427[310]) );
  DFFX1_LVT u_T_427_reg_26__53_ ( .D(n4466), .CLK(n4127), .Q(n_T_427[309]) );
  DFFX1_LVT u_T_427_reg_26__52_ ( .D(n4461), .CLK(n4127), .Q(n_T_427[308]) );
  DFFX1_LVT u_T_427_reg_26__51_ ( .D(n4458), .CLK(n4127), .Q(n_T_427[307]) );
  DFFX1_LVT u_T_427_reg_26__50_ ( .D(n4457), .CLK(n4127), .Q(n_T_427[306]) );
  DFFX1_LVT u_T_427_reg_26__49_ ( .D(n4452), .CLK(n4127), .Q(n_T_427[305]) );
  DFFX1_LVT u_T_427_reg_26__48_ ( .D(n4451), .CLK(n4127), .Q(n_T_427[304]) );
  DFFX1_LVT u_T_427_reg_26__47_ ( .D(n4448), .CLK(n4126), .Q(n_T_427[303]) );
  DFFX1_LVT u_T_427_reg_26__46_ ( .D(n4445), .CLK(n4126), .Q(n_T_427[302]) );
  DFFX1_LVT u_T_427_reg_26__45_ ( .D(n4440), .CLK(n4126), .Q(n_T_427[301]) );
  DFFX1_LVT u_T_427_reg_26__44_ ( .D(n4439), .CLK(n4126), .Q(n_T_427[300]) );
  DFFX1_LVT u_T_427_reg_26__43_ ( .D(n4434), .CLK(n4126), .Q(n_T_427[299]) );
  DFFX1_LVT u_T_427_reg_26__42_ ( .D(n4431), .CLK(n4126), .Q(n_T_427[298]) );
  DFFX1_LVT u_T_427_reg_26__41_ ( .D(n4428), .CLK(n4126), .Q(n_T_427[297]) );
  DFFX1_LVT u_T_427_reg_26__40_ ( .D(n4427), .CLK(n4126), .Q(n_T_427[296]) );
  DFFX1_LVT u_T_427_reg_26__39_ ( .D(n4424), .CLK(n4126), .Q(n_T_427[295]) );
  DFFX1_LVT u_T_427_reg_26__38_ ( .D(n4421), .CLK(n4126), .Q(n_T_427[294]) );
  DFFX1_LVT u_T_427_reg_26__37_ ( .D(n4419), .CLK(n4126), .Q(n_T_427[293]) );
  DFFX1_LVT u_T_427_reg_26__36_ ( .D(n4414), .CLK(n4126), .Q(n_T_427[292]) );
  DFFX1_LVT u_T_427_reg_26__35_ ( .D(n4413), .CLK(n4125), .Q(n_T_427[291]) );
  DFFX1_LVT u_T_427_reg_26__34_ ( .D(n4411), .CLK(n4125), .Q(n_T_427[290]) );
  DFFX1_LVT u_T_427_reg_26__33_ ( .D(n4408), .CLK(n4125), .Q(n_T_427[289]) );
  DFFX1_LVT u_T_427_reg_26__32_ ( .D(n4406), .CLK(n4125), .Q(n_T_427[288]) );
  DFFX1_LVT u_T_427_reg_26__31_ ( .D(n4403), .CLK(n4125), .Q(n_T_427[287]) );
  DFFX1_LVT u_T_427_reg_26__30_ ( .D(n4399), .CLK(n4125), .Q(n_T_427[286]) );
  DFFX1_LVT u_T_427_reg_26__29_ ( .D(n4396), .CLK(n4125), .Q(n_T_427[285]) );
  DFFX1_LVT u_T_427_reg_26__28_ ( .D(n4395), .CLK(n4125), .Q(n_T_427[284]) );
  DFFX1_LVT u_T_427_reg_26__27_ ( .D(n4393), .CLK(n4125), .Q(n_T_427[283]) );
  DFFX1_LVT u_T_427_reg_26__26_ ( .D(n4390), .CLK(n4125), .Q(n_T_427[282]) );
  DFFX1_LVT u_T_427_reg_26__25_ ( .D(n4388), .CLK(n4125), .Q(n_T_427[281]) );
  DFFX1_LVT u_T_427_reg_26__24_ ( .D(n4384), .CLK(n4125), .Q(n_T_427[280]) );
  DFFX1_LVT u_T_427_reg_26__23_ ( .D(n4383), .CLK(n4124), .Q(n_T_427[279]) );
  DFFX1_LVT u_T_427_reg_26__22_ ( .D(n4380), .CLK(n4124), .Q(n_T_427[278]) );
  DFFX1_LVT u_T_427_reg_26__21_ ( .D(n4378), .CLK(n4124), .Q(n_T_427[277]) );
  DFFX1_LVT u_T_427_reg_26__20_ ( .D(n4374), .CLK(n4124), .Q(n_T_427[276]) );
  DFFX1_LVT u_T_427_reg_26__19_ ( .D(n4371), .CLK(n4124), .Q(n_T_427[275]) );
  DFFX1_LVT u_T_427_reg_26__18_ ( .D(n4368), .CLK(n4124), .Q(n_T_427[274]) );
  DFFX1_LVT u_T_427_reg_26__17_ ( .D(n4367), .CLK(n4124), .Q(n_T_427[273]) );
  DFFX1_LVT u_T_427_reg_26__16_ ( .D(n4364), .CLK(n4124), .Q(n_T_427[272]) );
  DFFX1_LVT u_T_427_reg_26__15_ ( .D(n4361), .CLK(n4124), .Q(n_T_427[271]) );
  DFFX1_LVT u_T_427_reg_26__14_ ( .D(n4359), .CLK(n4124), .Q(n_T_427[270]) );
  DFFX1_LVT u_T_427_reg_26__13_ ( .D(n4356), .CLK(n4124), .Q(n_T_427[269]) );
  DFFX1_LVT u_T_427_reg_26__12_ ( .D(n4354), .CLK(n4124), .Q(n_T_427[268]) );
  DFFX1_LVT u_T_427_reg_26__11_ ( .D(n4349), .CLK(n4123), .Q(n_T_427[267]) );
  DFFX1_LVT u_T_427_reg_26__10_ ( .D(n4348), .CLK(n4123), .Q(n_T_427[266]) );
  DFFX1_LVT u_T_427_reg_26__9_ ( .D(n4345), .CLK(n4123), .Q(n_T_427[265]) );
  DFFX1_LVT u_T_427_reg_26__8_ ( .D(n4342), .CLK(n4123), .Q(n_T_427[264]) );
  DFFX1_LVT u_T_427_reg_26__7_ ( .D(n4339), .CLK(n4123), .Q(n_T_427[263]) );
  DFFX1_LVT u_T_427_reg_26__6_ ( .D(n4336), .CLK(n4123), .Q(n_T_427[262]) );
  DFFX1_LVT u_T_427_reg_26__5_ ( .D(n4333), .CLK(n4123), .Q(n_T_427[261]) );
  DFFX1_LVT u_T_427_reg_26__4_ ( .D(n4330), .CLK(n4123), .Q(n_T_427[260]) );
  DFFX1_LVT u_T_427_reg_26__3_ ( .D(n4327), .CLK(n4123), .Q(n_T_427[259]) );
  DFFX1_LVT u_T_427_reg_26__2_ ( .D(n4324), .CLK(n4123), .Q(n_T_427[258]) );
  DFFX1_LVT u_T_427_reg_26__1_ ( .D(n4319), .CLK(n4123), .Q(n_T_427[257]) );
  DFFX1_LVT u_T_427_reg_26__0_ ( .D(n4316), .CLK(n4123), .Q(n_T_427[256]) );
  DFFX1_LVT u_T_427_reg_27__63_ ( .D(n4496), .CLK(n4122), .Q(n_T_427[255]) );
  DFFX1_LVT u_T_427_reg_27__62_ ( .D(n4493), .CLK(n4122), .Q(n_T_427[254]) );
  DFFX1_LVT u_T_427_reg_27__61_ ( .D(n4490), .CLK(n4122), .Q(n_T_427[253]) );
  DFFX1_LVT u_T_427_reg_27__60_ ( .D(n4487), .CLK(n4122), .Q(n_T_427[252]) );
  DFFX1_LVT u_T_427_reg_27__59_ ( .D(n4484), .CLK(n4121), .Q(n_T_427[251]) );
  DFFX1_LVT u_T_427_reg_27__58_ ( .D(n4479), .CLK(n4121), .Q(n_T_427[250]) );
  DFFX1_LVT u_T_427_reg_27__57_ ( .D(n4478), .CLK(n4121), .Q(n_T_427[249]) );
  DFFX1_LVT u_T_427_reg_27__56_ ( .D(n4473), .CLK(n4121), .Q(n_T_427[248]) );
  DFFX1_LVT u_T_427_reg_27__55_ ( .D(n4472), .CLK(n4121), .Q(n_T_427[247]) );
  DFFX1_LVT u_T_427_reg_27__54_ ( .D(n4467), .CLK(n4121), .Q(n_T_427[246]) );
  DFFX1_LVT u_T_427_reg_27__53_ ( .D(n4466), .CLK(n4121), .Q(n_T_427[245]) );
  DFFX1_LVT u_T_427_reg_27__52_ ( .D(n4461), .CLK(n4121), .Q(n_T_427[244]) );
  DFFX1_LVT u_T_427_reg_27__51_ ( .D(n4458), .CLK(n4121), .Q(n_T_427[243]) );
  DFFX1_LVT u_T_427_reg_27__50_ ( .D(n4457), .CLK(n4121), .Q(n_T_427[242]) );
  DFFX1_LVT u_T_427_reg_27__49_ ( .D(n4452), .CLK(n4121), .Q(n_T_427[241]) );
  DFFX1_LVT u_T_427_reg_27__48_ ( .D(n4451), .CLK(n4121), .Q(n_T_427[240]) );
  DFFX1_LVT u_T_427_reg_27__47_ ( .D(n4448), .CLK(n4120), .Q(n_T_427[239]) );
  DFFX1_LVT u_T_427_reg_27__46_ ( .D(n4445), .CLK(n4120), .Q(n_T_427[238]), 
        .QN(n3522) );
  DFFX1_LVT u_T_427_reg_27__45_ ( .D(n4440), .CLK(n4120), .Q(n_T_427[237]) );
  DFFX1_LVT u_T_427_reg_27__44_ ( .D(n4439), .CLK(n4120), .Q(n_T_427[236]) );
  DFFX1_LVT u_T_427_reg_27__43_ ( .D(n4434), .CLK(n4120), .Q(n_T_427[235]) );
  DFFX1_LVT u_T_427_reg_27__42_ ( .D(n4431), .CLK(n4120), .Q(n_T_427[234]) );
  DFFX1_LVT u_T_427_reg_27__41_ ( .D(n4428), .CLK(n4120), .Q(n_T_427[233]) );
  DFFX1_LVT u_T_427_reg_27__40_ ( .D(n4427), .CLK(n4120), .Q(n_T_427[232]) );
  DFFX1_LVT u_T_427_reg_27__39_ ( .D(n4424), .CLK(n4120), .Q(n_T_427[231]), 
        .QN(n3523) );
  DFFX1_LVT u_T_427_reg_27__38_ ( .D(n4421), .CLK(n4120), .Q(n_T_427[230]) );
  DFFX1_LVT u_T_427_reg_27__37_ ( .D(n4419), .CLK(n4120), .Q(n_T_427[229]) );
  DFFX1_LVT u_T_427_reg_27__36_ ( .D(n4414), .CLK(n4120), .Q(n_T_427[228]) );
  DFFX1_LVT u_T_427_reg_27__35_ ( .D(n4413), .CLK(n4119), .Q(n_T_427[227]) );
  DFFX1_LVT u_T_427_reg_27__34_ ( .D(n4411), .CLK(n4119), .Q(n_T_427[226]) );
  DFFX1_LVT u_T_427_reg_27__33_ ( .D(n4408), .CLK(n4119), .Q(n_T_427[225]) );
  DFFX1_LVT u_T_427_reg_27__32_ ( .D(n4406), .CLK(n4119), .Q(n_T_427[224]) );
  DFFX1_LVT u_T_427_reg_27__31_ ( .D(n4403), .CLK(n4119), .Q(n_T_427[223]) );
  DFFX1_LVT u_T_427_reg_27__30_ ( .D(n4399), .CLK(n4119), .Q(n_T_427[222]) );
  DFFX1_LVT u_T_427_reg_27__29_ ( .D(n4396), .CLK(n4119), .Q(n_T_427[221]) );
  DFFX1_LVT u_T_427_reg_27__28_ ( .D(n4395), .CLK(n4119), .Q(n_T_427[220]) );
  DFFX1_LVT u_T_427_reg_27__27_ ( .D(n4393), .CLK(n4119), .Q(n_T_427[219]) );
  DFFX1_LVT u_T_427_reg_27__26_ ( .D(n4390), .CLK(n4119), .Q(n_T_427[218]) );
  DFFX1_LVT u_T_427_reg_27__25_ ( .D(n4388), .CLK(n4119), .Q(n_T_427[217]) );
  DFFX1_LVT u_T_427_reg_27__24_ ( .D(n4384), .CLK(n4119), .Q(n_T_427[216]) );
  DFFX1_LVT u_T_427_reg_27__23_ ( .D(n4383), .CLK(n4118), .Q(n_T_427[215]) );
  DFFX1_LVT u_T_427_reg_27__22_ ( .D(n4380), .CLK(n4118), .Q(n_T_427[214]) );
  DFFX1_LVT u_T_427_reg_27__21_ ( .D(n4378), .CLK(n4118), .Q(n_T_427[213]) );
  DFFX1_LVT u_T_427_reg_27__20_ ( .D(n4374), .CLK(n4118), .Q(n_T_427[212]) );
  DFFX1_LVT u_T_427_reg_27__19_ ( .D(n4371), .CLK(n4118), .Q(n_T_427[211]) );
  DFFX1_LVT u_T_427_reg_27__18_ ( .D(n4368), .CLK(n4118), .Q(n_T_427[210]) );
  DFFX1_LVT u_T_427_reg_27__17_ ( .D(n4367), .CLK(n4118), .Q(n_T_427[209]) );
  DFFX1_LVT u_T_427_reg_27__16_ ( .D(n4364), .CLK(n4118), .Q(n_T_427[208]), 
        .QN(n3521) );
  DFFX1_LVT u_T_427_reg_27__15_ ( .D(n4361), .CLK(n4118), .Q(n_T_427[207]) );
  DFFX1_LVT u_T_427_reg_27__14_ ( .D(n4359), .CLK(n4118), .Q(n_T_427[206]) );
  DFFX1_LVT u_T_427_reg_27__13_ ( .D(n4356), .CLK(n4118), .Q(n_T_427[205]) );
  DFFX1_LVT u_T_427_reg_27__12_ ( .D(n4354), .CLK(n4118), .Q(n_T_427[204]) );
  DFFX1_LVT u_T_427_reg_27__11_ ( .D(n4349), .CLK(n4117), .Q(n_T_427[203]) );
  DFFX1_LVT u_T_427_reg_27__10_ ( .D(n4348), .CLK(n4117), .Q(n_T_427[202]) );
  DFFX1_LVT u_T_427_reg_27__9_ ( .D(n4345), .CLK(n4117), .Q(n_T_427[201]) );
  DFFX1_LVT u_T_427_reg_27__8_ ( .D(n4342), .CLK(n4117), .Q(n_T_427[200]) );
  DFFX1_LVT u_T_427_reg_27__7_ ( .D(n4339), .CLK(n4117), .Q(n_T_427[199]) );
  DFFX1_LVT u_T_427_reg_27__6_ ( .D(n4336), .CLK(n4117), .Q(n_T_427[198]) );
  DFFX1_LVT u_T_427_reg_27__5_ ( .D(n4333), .CLK(n4117), .Q(n_T_427[197]) );
  DFFX1_LVT u_T_427_reg_27__4_ ( .D(n4330), .CLK(n4117), .Q(n_T_427[196]) );
  DFFX1_LVT u_T_427_reg_27__3_ ( .D(n4327), .CLK(n4117), .Q(n_T_427[195]) );
  DFFX1_LVT u_T_427_reg_27__2_ ( .D(n4324), .CLK(n4117), .Q(n_T_427[194]) );
  DFFX1_LVT u_T_427_reg_27__1_ ( .D(n4319), .CLK(n4117), .Q(n_T_427[193]) );
  DFFX1_LVT u_T_427_reg_27__0_ ( .D(n4316), .CLK(n4117), .Q(n_T_427[192]) );
  DFFX1_LVT u_T_427_reg_28__63_ ( .D(n4496), .CLK(n4116), .Q(n_T_427[191]) );
  DFFX1_LVT u_T_427_reg_28__62_ ( .D(n4493), .CLK(n4116), .Q(n_T_427[190]) );
  DFFX1_LVT u_T_427_reg_28__61_ ( .D(n4490), .CLK(n4116), .Q(n_T_427[189]) );
  DFFX1_LVT u_T_427_reg_28__60_ ( .D(n4487), .CLK(n4116), .Q(n_T_427[188]) );
  DFFX1_LVT u_T_427_reg_28__59_ ( .D(n4484), .CLK(n4115), .Q(n_T_427[187]) );
  DFFX1_LVT u_T_427_reg_28__58_ ( .D(n4479), .CLK(n4115), .Q(n_T_427[186]) );
  DFFX1_LVT u_T_427_reg_28__57_ ( .D(n4478), .CLK(n4115), .Q(n_T_427[185]) );
  DFFX1_LVT u_T_427_reg_28__56_ ( .D(n4473), .CLK(n4115), .Q(n_T_427[184]) );
  DFFX1_LVT u_T_427_reg_28__55_ ( .D(n4472), .CLK(n4115), .Q(n_T_427[183]) );
  DFFX1_LVT u_T_427_reg_28__54_ ( .D(n4467), .CLK(n4115), .Q(n_T_427[182]) );
  DFFX1_LVT u_T_427_reg_28__53_ ( .D(n4466), .CLK(n4115), .Q(n_T_427[181]) );
  DFFX1_LVT u_T_427_reg_28__52_ ( .D(n4461), .CLK(n4115), .Q(n_T_427[180]) );
  DFFX1_LVT u_T_427_reg_28__51_ ( .D(n4458), .CLK(n4115), .Q(n_T_427[179]) );
  DFFX1_LVT u_T_427_reg_28__50_ ( .D(n4457), .CLK(n4115), .Q(n_T_427[178]) );
  DFFX1_LVT u_T_427_reg_28__49_ ( .D(n4452), .CLK(n4115), .Q(n_T_427[177]) );
  DFFX1_LVT u_T_427_reg_28__48_ ( .D(n4451), .CLK(n4115), .Q(n_T_427[176]) );
  DFFX1_LVT u_T_427_reg_28__47_ ( .D(n4448), .CLK(n4114), .Q(n_T_427[175]) );
  DFFX1_LVT u_T_427_reg_28__46_ ( .D(n4445), .CLK(n4114), .Q(n_T_427[174]) );
  DFFX1_LVT u_T_427_reg_28__45_ ( .D(n4440), .CLK(n4114), .Q(n_T_427[173]) );
  DFFX1_LVT u_T_427_reg_28__44_ ( .D(n4439), .CLK(n4114), .Q(n_T_427[172]) );
  DFFX1_LVT u_T_427_reg_28__43_ ( .D(n4434), .CLK(n4114), .Q(n_T_427[171]) );
  DFFX1_LVT u_T_427_reg_28__42_ ( .D(n4431), .CLK(n4114), .Q(n_T_427[170]) );
  DFFX1_LVT u_T_427_reg_28__41_ ( .D(n4428), .CLK(n4114), .Q(n_T_427[169]) );
  DFFX1_LVT u_T_427_reg_28__40_ ( .D(n4427), .CLK(n4114), .Q(n_T_427[168]) );
  DFFX1_LVT u_T_427_reg_28__39_ ( .D(n4424), .CLK(n4114), .Q(n_T_427[167]) );
  DFFX1_LVT u_T_427_reg_28__38_ ( .D(n4421), .CLK(n4114), .Q(n_T_427[166]) );
  DFFX1_LVT u_T_427_reg_28__37_ ( .D(n4419), .CLK(n4114), .Q(n_T_427[165]) );
  DFFX1_LVT u_T_427_reg_28__36_ ( .D(n4414), .CLK(n4114), .Q(n_T_427[164]) );
  DFFX1_LVT u_T_427_reg_28__35_ ( .D(n4413), .CLK(n4113), .Q(n_T_427[163]) );
  DFFX1_LVT u_T_427_reg_28__34_ ( .D(n4411), .CLK(n4113), .Q(n_T_427[162]) );
  DFFX1_LVT u_T_427_reg_28__33_ ( .D(n4408), .CLK(n4113), .Q(n_T_427[161]) );
  DFFX1_LVT u_T_427_reg_28__32_ ( .D(n4406), .CLK(n4113), .Q(n_T_427[160]) );
  DFFX1_LVT u_T_427_reg_28__31_ ( .D(n4403), .CLK(n4113), .Q(n_T_427[159]) );
  DFFX1_LVT u_T_427_reg_28__30_ ( .D(n4399), .CLK(n4113), .Q(n_T_427[158]) );
  DFFX1_LVT u_T_427_reg_28__29_ ( .D(n4396), .CLK(n4113), .Q(n_T_427[157]) );
  DFFX1_LVT u_T_427_reg_28__28_ ( .D(n4395), .CLK(n4113), .Q(n_T_427[156]) );
  DFFX1_LVT u_T_427_reg_28__27_ ( .D(n4393), .CLK(n4113), .Q(n_T_427[155]) );
  DFFX1_LVT u_T_427_reg_28__26_ ( .D(n4390), .CLK(n4113), .Q(n_T_427[154]) );
  DFFX1_LVT u_T_427_reg_28__25_ ( .D(n4388), .CLK(n4113), .Q(n_T_427[153]) );
  DFFX1_LVT u_T_427_reg_28__24_ ( .D(n4384), .CLK(n4113), .Q(n_T_427[152]) );
  DFFX1_LVT u_T_427_reg_28__23_ ( .D(n4383), .CLK(n4112), .Q(n_T_427[151]), 
        .QN(n3526) );
  DFFX1_LVT u_T_427_reg_28__22_ ( .D(n4380), .CLK(n4112), .Q(n_T_427[150]) );
  DFFX1_LVT u_T_427_reg_28__21_ ( .D(n4378), .CLK(n4112), .Q(n_T_427[149]) );
  DFFX1_LVT u_T_427_reg_28__20_ ( .D(n4374), .CLK(n4112), .Q(n_T_427[148]) );
  DFFX1_LVT u_T_427_reg_28__19_ ( .D(n4371), .CLK(n4112), .Q(n_T_427[147]) );
  DFFX1_LVT u_T_427_reg_28__18_ ( .D(n4368), .CLK(n4112), .Q(n_T_427[146]) );
  DFFX1_LVT u_T_427_reg_28__17_ ( .D(n4367), .CLK(n4112), .Q(n_T_427[145]) );
  DFFX1_LVT u_T_427_reg_28__16_ ( .D(n4364), .CLK(n4112), .Q(n_T_427[144]) );
  DFFX1_LVT u_T_427_reg_28__15_ ( .D(n4361), .CLK(n4112), .Q(n_T_427[143]) );
  DFFX1_LVT u_T_427_reg_28__14_ ( .D(n4359), .CLK(n4112), .Q(n_T_427[142]) );
  DFFX1_LVT u_T_427_reg_28__13_ ( .D(n4356), .CLK(n4112), .Q(n_T_427[141]) );
  DFFX1_LVT u_T_427_reg_28__12_ ( .D(n4354), .CLK(n4112), .Q(n_T_427[140]) );
  DFFX1_LVT u_T_427_reg_28__11_ ( .D(n4349), .CLK(n4111), .Q(n_T_427[139]) );
  DFFX1_LVT u_T_427_reg_28__10_ ( .D(n4348), .CLK(n4111), .Q(n_T_427[138]) );
  DFFX1_LVT u_T_427_reg_28__9_ ( .D(n4345), .CLK(n4111), .Q(n_T_427[137]) );
  DFFX1_LVT u_T_427_reg_28__8_ ( .D(n4342), .CLK(n4111), .Q(n_T_427[136]) );
  DFFX1_LVT u_T_427_reg_28__7_ ( .D(n4339), .CLK(n4111), .Q(n_T_427[135]) );
  DFFX1_LVT u_T_427_reg_28__6_ ( .D(n4336), .CLK(n4111), .Q(n_T_427[134]) );
  DFFX1_LVT u_T_427_reg_28__5_ ( .D(n4333), .CLK(n4111), .Q(n_T_427[133]) );
  DFFX1_LVT u_T_427_reg_28__4_ ( .D(n4330), .CLK(n4111), .Q(n_T_427[132]) );
  DFFX1_LVT u_T_427_reg_28__3_ ( .D(n4327), .CLK(n4111), .Q(n_T_427[131]) );
  DFFX1_LVT u_T_427_reg_28__2_ ( .D(n4324), .CLK(n4111), .Q(n_T_427[130]) );
  DFFX1_LVT u_T_427_reg_28__1_ ( .D(n4319), .CLK(n4111), .Q(n_T_427[129]) );
  DFFX1_LVT u_T_427_reg_28__0_ ( .D(n4316), .CLK(n4111), .Q(n_T_427[128]) );
  DFFX1_LVT u_T_427_reg_29__63_ ( .D(n4496), .CLK(n4110), .Q(n_T_427[127]) );
  DFFX1_LVT u_T_427_reg_29__62_ ( .D(n4493), .CLK(n4110), .Q(n_T_427[126]) );
  DFFX1_LVT u_T_427_reg_29__61_ ( .D(n4490), .CLK(n4110), .Q(n_T_427[125]) );
  DFFX1_LVT u_T_427_reg_29__60_ ( .D(n4487), .CLK(n4110), .Q(n_T_427[124]) );
  DFFX1_LVT u_T_427_reg_29__59_ ( .D(n4484), .CLK(n4109), .Q(n_T_427[123]) );
  DFFX1_LVT u_T_427_reg_29__58_ ( .D(n4479), .CLK(n4109), .Q(n_T_427[122]) );
  DFFX1_LVT u_T_427_reg_29__57_ ( .D(n4478), .CLK(n4109), .Q(n_T_427[121]) );
  DFFX1_LVT u_T_427_reg_29__56_ ( .D(n4473), .CLK(n4109), .Q(n_T_427[120]) );
  DFFX1_LVT u_T_427_reg_29__55_ ( .D(n4472), .CLK(n4109), .Q(n_T_427[119]) );
  DFFX1_LVT u_T_427_reg_29__54_ ( .D(n4467), .CLK(n4109), .Q(n_T_427[118]) );
  DFFX1_LVT u_T_427_reg_29__53_ ( .D(n4466), .CLK(n4109), .Q(n_T_427[117]) );
  DFFX1_LVT u_T_427_reg_29__52_ ( .D(n4461), .CLK(n4109), .Q(n_T_427[116]) );
  DFFX1_LVT u_T_427_reg_29__51_ ( .D(n4458), .CLK(n4109), .Q(n_T_427[115]) );
  DFFX1_LVT u_T_427_reg_29__50_ ( .D(n4457), .CLK(n4109), .Q(n_T_427[114]) );
  DFFX1_LVT u_T_427_reg_29__49_ ( .D(n4452), .CLK(n4109), .Q(n_T_427[113]) );
  DFFX1_LVT u_T_427_reg_29__48_ ( .D(n4451), .CLK(n4109), .Q(n_T_427[112]) );
  DFFX1_LVT u_T_427_reg_29__47_ ( .D(n4448), .CLK(n4108), .Q(n_T_427[111]) );
  DFFX1_LVT u_T_427_reg_29__46_ ( .D(n4445), .CLK(n4108), .Q(n_T_427[110]), 
        .QN(n3176) );
  DFFX1_LVT u_T_427_reg_29__45_ ( .D(n4440), .CLK(n4108), .Q(n_T_427[109]) );
  DFFX1_LVT u_T_427_reg_29__44_ ( .D(n4439), .CLK(n4108), .Q(n_T_427[108]) );
  DFFX1_LVT u_T_427_reg_29__43_ ( .D(n4434), .CLK(n4108), .Q(n_T_427[107]) );
  DFFX1_LVT u_T_427_reg_29__42_ ( .D(n4431), .CLK(n4108), .Q(n_T_427[106]) );
  DFFX1_LVT u_T_427_reg_29__41_ ( .D(n4428), .CLK(n4108), .Q(n_T_427[105]) );
  DFFX1_LVT u_T_427_reg_29__40_ ( .D(n4427), .CLK(n4108), .Q(n_T_427[104]) );
  DFFX1_LVT u_T_427_reg_29__39_ ( .D(n4424), .CLK(n4108), .Q(n_T_427[103]) );
  DFFX1_LVT u_T_427_reg_29__38_ ( .D(n4421), .CLK(n4108), .Q(n_T_427[102]) );
  DFFX1_LVT u_T_427_reg_29__37_ ( .D(n4419), .CLK(n4108), .Q(n_T_427[101]) );
  DFFX1_LVT u_T_427_reg_29__36_ ( .D(n4414), .CLK(n4108), .Q(n_T_427[100]) );
  DFFX1_LVT u_T_427_reg_29__35_ ( .D(n4413), .CLK(n4107), .Q(n_T_427[99]) );
  DFFX1_LVT u_T_427_reg_29__34_ ( .D(n4411), .CLK(n4107), .Q(n_T_427[98]) );
  DFFX1_LVT u_T_427_reg_29__33_ ( .D(n4408), .CLK(n4107), .Q(n_T_427[97]) );
  DFFX1_LVT u_T_427_reg_29__32_ ( .D(n4406), .CLK(n4107), .Q(n_T_427[96]) );
  DFFX1_LVT u_T_427_reg_29__31_ ( .D(n4403), .CLK(n4107), .Q(n_T_427[95]) );
  DFFX1_LVT u_T_427_reg_29__30_ ( .D(n4399), .CLK(n4107), .Q(n_T_427[94]) );
  DFFX1_LVT u_T_427_reg_29__29_ ( .D(n4396), .CLK(n4107), .Q(n_T_427[93]) );
  DFFX1_LVT u_T_427_reg_29__28_ ( .D(n4395), .CLK(n4107), .Q(n_T_427[92]) );
  DFFX1_LVT u_T_427_reg_29__27_ ( .D(n4393), .CLK(n4107), .Q(n_T_427[91]) );
  DFFX1_LVT u_T_427_reg_29__26_ ( .D(n4390), .CLK(n4107), .Q(n_T_427[90]) );
  DFFX1_LVT u_T_427_reg_29__25_ ( .D(n4388), .CLK(n4107), .Q(n_T_427[89]) );
  DFFX1_LVT u_T_427_reg_29__24_ ( .D(n4384), .CLK(n4107), .Q(n_T_427[88]) );
  DFFX1_LVT u_T_427_reg_29__23_ ( .D(n4383), .CLK(n4106), .Q(n_T_427[87]) );
  DFFX1_LVT u_T_427_reg_29__22_ ( .D(n4380), .CLK(n4106), .Q(n_T_427[86]) );
  DFFX1_LVT u_T_427_reg_29__21_ ( .D(n4378), .CLK(n4106), .Q(n_T_427[85]) );
  DFFX1_LVT u_T_427_reg_29__20_ ( .D(n4374), .CLK(n4106), .Q(n_T_427[84]) );
  DFFX1_LVT u_T_427_reg_29__19_ ( .D(n4371), .CLK(n4106), .Q(n_T_427[83]) );
  DFFX1_LVT u_T_427_reg_29__18_ ( .D(n4368), .CLK(n4106), .Q(n_T_427[82]) );
  DFFX1_LVT u_T_427_reg_29__17_ ( .D(n4367), .CLK(n4106), .Q(n_T_427[81]) );
  DFFX1_LVT u_T_427_reg_29__16_ ( .D(n4364), .CLK(n4106), .Q(n_T_427[80]), 
        .QN(n3175) );
  DFFX1_LVT u_T_427_reg_29__15_ ( .D(n4361), .CLK(n4106), .Q(n_T_427[79]) );
  DFFX1_LVT u_T_427_reg_29__14_ ( .D(n4359), .CLK(n4106), .Q(n_T_427[78]) );
  DFFX1_LVT u_T_427_reg_29__13_ ( .D(n4356), .CLK(n4106), .Q(n_T_427[77]) );
  DFFX1_LVT u_T_427_reg_29__12_ ( .D(n4354), .CLK(n4106), .Q(n_T_427[76]) );
  DFFX1_LVT u_T_427_reg_29__11_ ( .D(n4349), .CLK(n4105), .Q(n_T_427[75]) );
  DFFX1_LVT u_T_427_reg_29__10_ ( .D(n4348), .CLK(n4105), .Q(n_T_427[74]) );
  DFFX1_LVT u_T_427_reg_29__9_ ( .D(n4345), .CLK(n4105), .Q(n_T_427[73]) );
  DFFX1_LVT u_T_427_reg_29__8_ ( .D(n4342), .CLK(n4105), .Q(n_T_427[72]) );
  DFFX1_LVT u_T_427_reg_29__7_ ( .D(n4339), .CLK(n4105), .Q(n_T_427[71]) );
  DFFX1_LVT u_T_427_reg_29__6_ ( .D(n4336), .CLK(n4105), .Q(n_T_427[70]) );
  DFFX1_LVT u_T_427_reg_29__5_ ( .D(n4333), .CLK(n4105), .Q(n_T_427[69]) );
  DFFX1_LVT u_T_427_reg_29__4_ ( .D(n4330), .CLK(n4105), .Q(n_T_427[68]) );
  DFFX1_LVT u_T_427_reg_29__3_ ( .D(n4327), .CLK(n4105), .Q(n_T_427[67]) );
  DFFX1_LVT u_T_427_reg_29__2_ ( .D(n4324), .CLK(n4105), .Q(n_T_427[66]) );
  DFFX1_LVT u_T_427_reg_29__1_ ( .D(n4319), .CLK(n4105), .Q(n_T_427[65]) );
  DFFX1_LVT u_T_427_reg_29__0_ ( .D(n4316), .CLK(n4105), .Q(n_T_427[64]) );
  DFFX1_LVT u_T_427_reg_30__63_ ( .D(n4496), .CLK(n4104), .Q(n_T_427[63]) );
  DFFX1_LVT u_T_427_reg_30__62_ ( .D(n4493), .CLK(n4104), .Q(n_T_427[62]) );
  DFFX1_LVT u_T_427_reg_30__61_ ( .D(n4490), .CLK(n4104), .Q(n_T_427[61]) );
  DFFX1_LVT u_T_427_reg_30__60_ ( .D(n4487), .CLK(n4104), .Q(n_T_427[60]) );
  DFFX1_LVT u_T_427_reg_30__59_ ( .D(n4484), .CLK(n4103), .Q(n_T_427[59]) );
  DFFX1_LVT u_T_427_reg_30__58_ ( .D(n4479), .CLK(n4103), .Q(n_T_427[58]) );
  DFFX1_LVT u_T_427_reg_30__57_ ( .D(n4478), .CLK(n4103), .Q(n_T_427[57]) );
  DFFX1_LVT u_T_427_reg_30__56_ ( .D(n4473), .CLK(n4103), .Q(n_T_427[56]) );
  DFFX1_LVT u_T_427_reg_30__55_ ( .D(n4472), .CLK(n4103), .Q(n_T_427[55]) );
  DFFX1_LVT u_T_427_reg_30__54_ ( .D(n4467), .CLK(n4103), .Q(n_T_427[54]) );
  DFFX1_LVT u_T_427_reg_30__53_ ( .D(n4466), .CLK(n4103), .Q(n_T_427[53]) );
  DFFX1_LVT u_T_427_reg_30__52_ ( .D(n4461), .CLK(n4103), .Q(n_T_427[52]) );
  DFFX1_LVT u_T_427_reg_30__51_ ( .D(n4458), .CLK(n4103), .Q(n_T_427[51]) );
  DFFX1_LVT u_T_427_reg_30__50_ ( .D(n4457), .CLK(n4103), .Q(n_T_427[50]) );
  DFFX1_LVT u_T_427_reg_30__49_ ( .D(n4452), .CLK(n4103), .Q(n_T_427[49]) );
  DFFX1_LVT u_T_427_reg_30__48_ ( .D(n4451), .CLK(n4103), .Q(n_T_427[48]) );
  DFFX1_LVT u_T_427_reg_30__47_ ( .D(n4448), .CLK(n4102), .Q(n_T_427[47]) );
  DFFX1_LVT u_T_427_reg_30__46_ ( .D(n4445), .CLK(n4102), .Q(n_T_427[46]) );
  DFFX1_LVT u_T_427_reg_30__45_ ( .D(n4440), .CLK(n4102), .Q(n_T_427[45]) );
  DFFX1_LVT u_T_427_reg_30__44_ ( .D(n4439), .CLK(n4102), .Q(n_T_427[44]) );
  DFFX1_LVT u_T_427_reg_30__43_ ( .D(n4434), .CLK(n4102), .Q(n_T_427[43]) );
  DFFX1_LVT u_T_427_reg_30__42_ ( .D(n4431), .CLK(n4102), .Q(n_T_427[42]) );
  DFFX1_LVT u_T_427_reg_30__41_ ( .D(n4428), .CLK(n4102), .Q(n_T_427[41]) );
  DFFX1_LVT u_T_427_reg_30__40_ ( .D(n4427), .CLK(n4102), .Q(n_T_427[40]) );
  DFFX1_LVT u_T_427_reg_30__39_ ( .D(n4424), .CLK(n4102), .Q(n_T_427[39]) );
  DFFX1_LVT u_T_427_reg_30__38_ ( .D(n4421), .CLK(n4102), .Q(n_T_427[38]) );
  DFFX1_LVT u_T_427_reg_30__37_ ( .D(n4419), .CLK(n4102), .Q(n_T_427[37]) );
  DFFX1_LVT u_T_427_reg_30__36_ ( .D(n4414), .CLK(n4102), .Q(n_T_427[36]) );
  DFFX1_LVT u_T_427_reg_30__35_ ( .D(n4413), .CLK(n4101), .Q(n_T_427[35]) );
  DFFX1_LVT u_T_427_reg_30__34_ ( .D(n4411), .CLK(n4101), .Q(n_T_427[34]) );
  DFFX1_LVT u_T_427_reg_30__33_ ( .D(n4408), .CLK(n4101), .Q(n_T_427[33]) );
  DFFX1_LVT u_T_427_reg_30__32_ ( .D(n4406), .CLK(n4101), .Q(n_T_427[32]) );
  DFFX1_LVT u_T_427_reg_30__31_ ( .D(n4403), .CLK(n4101), .Q(n_T_427[31]) );
  DFFX1_LVT u_T_427_reg_30__30_ ( .D(n4399), .CLK(n4101), .Q(n_T_427[30]) );
  DFFX1_LVT u_T_427_reg_30__29_ ( .D(n4396), .CLK(n4101), .Q(n_T_427[29]) );
  DFFX1_LVT u_T_427_reg_30__28_ ( .D(n4395), .CLK(n4101), .Q(n_T_427[28]) );
  DFFX1_LVT u_T_427_reg_30__27_ ( .D(n4393), .CLK(n4101), .Q(n_T_427[27]) );
  DFFX1_LVT u_T_427_reg_30__26_ ( .D(n4390), .CLK(n4101), .Q(n_T_427[26]) );
  DFFX1_LVT u_T_427_reg_30__25_ ( .D(n4388), .CLK(n4101), .Q(n_T_427[25]) );
  DFFX1_LVT u_T_427_reg_30__24_ ( .D(n4384), .CLK(n4101), .Q(n_T_427[24]) );
  DFFX1_LVT u_T_427_reg_30__23_ ( .D(n4383), .CLK(n4100), .Q(n_T_427[23]), 
        .QN(n3177) );
  DFFX1_LVT u_T_427_reg_30__22_ ( .D(n4380), .CLK(n4100), .Q(n_T_427[22]) );
  DFFX1_LVT u_T_427_reg_30__21_ ( .D(n4378), .CLK(n4100), .Q(n_T_427[21]) );
  DFFX1_LVT u_T_427_reg_30__20_ ( .D(n4374), .CLK(n4100), .Q(n_T_427[20]) );
  DFFX1_LVT u_T_427_reg_30__19_ ( .D(n4371), .CLK(n4100), .Q(n_T_427[19]) );
  DFFX1_LVT u_T_427_reg_30__18_ ( .D(n4368), .CLK(n4100), .Q(n_T_427[18]) );
  DFFX1_LVT u_T_427_reg_30__17_ ( .D(n4367), .CLK(n4100), .Q(n_T_427[17]) );
  DFFX1_LVT u_T_427_reg_30__16_ ( .D(n4364), .CLK(n4100), .Q(n_T_427[16]) );
  DFFX1_LVT u_T_427_reg_30__15_ ( .D(n4361), .CLK(n4100), .Q(n_T_427[15]) );
  DFFX1_LVT u_T_427_reg_30__14_ ( .D(n4359), .CLK(n4100), .Q(n_T_427[14]) );
  DFFX1_LVT u_T_427_reg_30__13_ ( .D(n4356), .CLK(n4100), .Q(n_T_427[13]) );
  DFFX1_LVT u_T_427_reg_30__12_ ( .D(n4354), .CLK(n4100), .Q(n_T_427[12]) );
  DFFX1_LVT u_T_427_reg_30__11_ ( .D(n4349), .CLK(n4099), .Q(n_T_427[11]) );
  DFFX1_LVT u_T_427_reg_30__10_ ( .D(n4348), .CLK(n4099), .Q(n_T_427[10]) );
  DFFX1_LVT u_T_427_reg_30__9_ ( .D(n4345), .CLK(n4099), .Q(n_T_427[9]) );
  DFFX1_LVT u_T_427_reg_30__8_ ( .D(n4342), .CLK(n4099), .Q(n_T_427[8]) );
  DFFX1_LVT u_T_427_reg_30__7_ ( .D(n4339), .CLK(n4099), .Q(n_T_427[7]) );
  DFFX1_LVT u_T_427_reg_30__6_ ( .D(n4336), .CLK(n4099), .Q(n_T_427[6]) );
  DFFX1_LVT u_T_427_reg_30__5_ ( .D(n4333), .CLK(n4099), .Q(n_T_427[5]) );
  DFFX1_LVT u_T_427_reg_30__4_ ( .D(n4330), .CLK(n4099), .Q(n_T_427[4]) );
  DFFX1_LVT u_T_427_reg_30__3_ ( .D(n4327), .CLK(n4099), .Q(n_T_427[3]) );
  DFFX1_LVT u_T_427_reg_30__2_ ( .D(n4324), .CLK(n4099), .Q(n_T_427[2]) );
  DFFX1_LVT u_T_427_reg_30__1_ ( .D(n4319), .CLK(n4099), .Q(n_T_427[1]) );
  DFFX1_LVT u_T_427_reg_30__0_ ( .D(n4316), .CLK(n4099), .Q(n_T_427[0]) );
  DFFX1_LVT u_T_1185_reg_31_ ( .D(N777), .CLK(n4071), .Q(n_T_1187[31]), .QN(
        n3267) );
  DFFX1_LVT u_T_1185_reg_30_ ( .D(N776), .CLK(n4071), .Q(n_T_1187[30]) );
  DFFX1_LVT u_T_1185_reg_29_ ( .D(N775), .CLK(n4071), .Q(n_T_1187[29]), .QN(
        n3131) );
  DFFX1_LVT u_T_1185_reg_28_ ( .D(N774), .CLK(n4071), .Q(n_T_1187[28]), .QN(
        n3274) );
  DFFX1_LVT u_T_1185_reg_26_ ( .D(N772), .CLK(n4071), .Q(n_T_1187[26]), .QN(
        n3265) );
  DFFX1_LVT u_T_1185_reg_25_ ( .D(N771), .CLK(n4071), .Q(n_T_1187[25]), .QN(
        n3089) );
  DFFX1_LVT u_T_1185_reg_24_ ( .D(N770), .CLK(n4071), .Q(n_T_1187[24]), .QN(
        n3275) );
  DFFX1_LVT u_T_1185_reg_23_ ( .D(N769), .CLK(n4071), .Q(n_T_1187[23]), .QN(
        n3268) );
  DFFX1_LVT u_T_1185_reg_22_ ( .D(N768), .CLK(n4071), .Q(n_T_1187[22]) );
  DFFX1_LVT u_T_1185_reg_21_ ( .D(N767), .CLK(n4071), .Q(n_T_1187[21]), .QN(
        n3130) );
  DFFX1_LVT u_T_1185_reg_20_ ( .D(N766), .CLK(n4071), .Q(n_T_1187[20]), .QN(
        n3273) );
  DFFX1_LVT u_T_1185_reg_19_ ( .D(N765), .CLK(n4072), .Q(n_T_1187[19]), .QN(
        n3258) );
  DFFX1_LVT u_T_1185_reg_18_ ( .D(N764), .CLK(n4072), .Q(n_T_1187[18]), .QN(
        n3263) );
  DFFX1_LVT u_T_1185_reg_17_ ( .D(N763), .CLK(n4072), .Q(n_T_1187[17]), .QN(
        n3113) );
  DFFX1_LVT u_T_1185_reg_16_ ( .D(N762), .CLK(n4072), .Q(n_T_1187[16]), .QN(
        n3261) );
  DFFX1_LVT u_T_1185_reg_15_ ( .D(N761), .CLK(n4072), .Q(n_T_1187[15]), .QN(
        n3266) );
  DFFX1_LVT u_T_1185_reg_14_ ( .D(N760), .CLK(n4072), .Q(n_T_1187[14]), .QN(
        n3127) );
  DFFX1_LVT u_T_1185_reg_13_ ( .D(N759), .CLK(n4072), .Q(n_T_1187[13]), .QN(
        n3272) );
  DFFX1_LVT u_T_1185_reg_12_ ( .D(N758), .CLK(n4072), .Q(n_T_1187[12]), .QN(
        n3260) );
  DFFX1_LVT u_T_1185_reg_11_ ( .D(N757), .CLK(n4072), .Q(n_T_1187[11]), .QN(
        n3259) );
  DFFX1_LVT u_T_1185_reg_10_ ( .D(N756), .CLK(n4072), .Q(n_T_1187[10]), .QN(
        n3129) );
  DFFX1_LVT u_T_1185_reg_9_ ( .D(N755), .CLK(n4072), .Q(n_T_1187[9]), .QN(
        n3133) );
  DFFX1_LVT u_T_1185_reg_8_ ( .D(N754), .CLK(n4072), .Q(n_T_1187[8]), .QN(
        n3134) );
  DFFX1_LVT u_T_1185_reg_7_ ( .D(N753), .CLK(n4073), .Q(n_T_1187[7]), .QN(
        n3270) );
  DFFX1_LVT u_T_1185_reg_6_ ( .D(N752), .CLK(n4073), .Q(n_T_1187[6]), .QN(
        n3136) );
  DFFX1_LVT u_T_1185_reg_5_ ( .D(N751), .CLK(n4073), .Q(n_T_1187[5]), .QN(
        n3271) );
  DFFX1_LVT u_T_1185_reg_4_ ( .D(N750), .CLK(n4073), .Q(n_T_1187[4]), .QN(
        n3132) );
  DFFX1_LVT u_T_1185_reg_3_ ( .D(N749), .CLK(n4073), .Q(n_T_1187[3]), .QN(
        n3269) );
  DFFX1_LVT u_T_1185_reg_2_ ( .D(N748), .CLK(n4073), .Q(n_T_1187[2]), .QN(
        n3264) );
  DFFX1_LVT u_T_1185_reg_1_ ( .D(N747), .CLK(n4073), .Q(n_T_1187[1]), .QN(
        n3128) );
  DFFX1_LVT u_T_1298_reg_31_ ( .D(N810), .CLK(n4068), .Q(n_T_1298[31]), .QN(
        n3241) );
  DFFX1_LVT u_T_1298_reg_30_ ( .D(N809), .CLK(n4068), .Q(n_T_1298[30]), .QN(
        n3118) );
  DFFX1_LVT u_T_1298_reg_29_ ( .D(N808), .CLK(n4068), .Q(n_T_1298[29]), .QN(
        n3084) );
  DFFX1_LVT u_T_1298_reg_28_ ( .D(N807), .CLK(n4068), .Q(n_T_1298[28]), .QN(
        n3123) );
  DFFX1_LVT u_T_1298_reg_27_ ( .D(N806), .CLK(n4068), .Q(n_T_1298[27]), .QN(
        n3085) );
  DFFX1_LVT u_T_1298_reg_26_ ( .D(N805), .CLK(n4068), .Q(n_T_1298[26]), .QN(
        n3232) );
  DFFX1_LVT u_T_1298_reg_25_ ( .D(N804), .CLK(n4068), .Q(n_T_1298[25]), .QN(
        n3116) );
  DFFX1_LVT u_T_1298_reg_24_ ( .D(N803), .CLK(n4068), .Q(n_T_1298[24]), .QN(
        n3237) );
  DFFX1_LVT u_T_1298_reg_23_ ( .D(N802), .CLK(n4068), .Q(n_T_1298[23]), .QN(
        n3239) );
  DFFX1_LVT u_T_1298_reg_22_ ( .D(N801), .CLK(n4068), .Q(n_T_1298[22]), .QN(
        n3117) );
  DFFX1_LVT u_T_1298_reg_21_ ( .D(N800), .CLK(n4068), .Q(n_T_1298[21]), .QN(
        n3114) );
  DFFX1_LVT u_T_1298_reg_20_ ( .D(N799), .CLK(n4068), .Q(n_T_1298[20]), .QN(
        n3238) );
  DFFX1_LVT u_T_1298_reg_19_ ( .D(N798), .CLK(n4069), .Q(n_T_1298[19]), .QN(
        n3126) );
  DFFX1_LVT u_T_1298_reg_18_ ( .D(N797), .CLK(n4069), .Q(n_T_1298[18]), .QN(
        n3250) );
  DFFX1_LVT u_T_1298_reg_17_ ( .D(N796), .CLK(n4069), .Q(n_T_1298[17]), .QN(
        n3087) );
  DFFX1_LVT u_T_1298_reg_16_ ( .D(N795), .CLK(n4069), .Q(n_T_1298[16]), .QN(
        n3252) );
  DFFX1_LVT u_T_1298_reg_15_ ( .D(N794), .CLK(n4069), .Q(n_T_1298[15]), .QN(
        n3236) );
  DFFX1_LVT u_T_1298_reg_14_ ( .D(N793), .CLK(n4069), .Q(n_T_1298[14]), .QN(
        n3121) );
  DFFX1_LVT u_T_1298_reg_13_ ( .D(N792), .CLK(n4069), .Q(n_T_1298[13]), .QN(
        n3120) );
  DFFX1_LVT u_T_1298_reg_12_ ( .D(N791), .CLK(n4069), .Q(n_T_1298[12]), .QN(
        n3235) );
  DFFX1_LVT u_T_1298_reg_11_ ( .D(N790), .CLK(n4069), .Q(n_T_1298[11]), .QN(
        n3240) );
  DFFX1_LVT u_T_1298_reg_10_ ( .D(N789), .CLK(n4069), .Q(n_T_1298[10]), .QN(
        n3115) );
  DFFX1_LVT u_T_1298_reg_9_ ( .D(N788), .CLK(n4069), .Q(n_T_1298[9]), .QN(
        n3119) );
  DFFX1_LVT u_T_1298_reg_8_ ( .D(N787), .CLK(n4069), .Q(n_T_1298[8]), .QN(
        n3242) );
  DFFX1_LVT u_T_1298_reg_7_ ( .D(N786), .CLK(n4070), .Q(n_T_1298[7]), .QN(
        n3125) );
  DFFX1_LVT u_T_1298_reg_6_ ( .D(N785), .CLK(n4070), .Q(n_T_1298[6]), .QN(
        n3248) );
  DFFX1_LVT u_T_1298_reg_5_ ( .D(N784), .CLK(n4070), .Q(n_T_1298[5]), .QN(
        n3088) );
  DFFX1_LVT u_T_1298_reg_4_ ( .D(N783), .CLK(n4070), .Q(n_T_1298[4]), .QN(
        n3253) );
  DFFX1_LVT u_T_1298_reg_3_ ( .D(N782), .CLK(n4070), .Q(n_T_1298[3]), .QN(
        n3124) );
  DFFX1_LVT u_T_1298_reg_2_ ( .D(N781), .CLK(n4070), .Q(n_T_1298[2]), .QN(
        n3247) );
  DFFX1_LVT u_T_1298_reg_1_ ( .D(N780), .CLK(n4070), .Q(n_T_1298[1]), .QN(
        n3086) );
  DFFX1_LVT u_T_1298_reg_0_ ( .D(N779), .CLK(n4070), .Q(n_T_1298[0]), .QN(
        n3254) );
  AO22X1_LVT U613 ( .A1(csr_io_pc[0]), .A2(n4062), .A3(1'b0), .A4(n4065), .Y(
        io_imem_req_bits_pc[0]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_61_ ( .D(N743), .CLK(n4085), .Q(n_T_628[63])
         );
  DFFX1_LVT ex_reg_mem_size_reg_1_ ( .D(N370), .CLK(n4314), .Q(
        io_dmem_req_bits_size[1]), .QN(n586) );
  DFFX1_LVT u_T_427_reg_0__50_ ( .D(n4455), .CLK(n4283), .QN(n3277) );
  DFFX1_LVT u_T_427_reg_0__32_ ( .D(n4404), .CLK(n4281), .QN(n3276) );
  DFFX1_LVT u_T_427_reg_19__34_ ( .D(n4410), .CLK(n4167), .QN(n3141) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_39_ ( .D(N721), .CLK(n4083), .Q(n_T_628[41])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_53_ ( .D(N735), .CLK(n4084), .Q(n_T_628[55])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_33_ ( .D(N715), .CLK(n4082), .Q(n_T_628[35])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_56_ ( .D(N738), .CLK(n4084), .Q(n_T_628[58])
         );
  DFFX1_LVT u_T_427_reg_0__55_ ( .D(n4470), .CLK(n4283), .Q(n_T_427[1934]), 
        .QN(n3563) );
  DFFX1_LVT u_T_427_reg_0__53_ ( .D(n4464), .CLK(n4283), .Q(n_T_427[1932]), 
        .QN(n3561) );
  DFFX1_LVT u_T_427_reg_0__48_ ( .D(n4449), .CLK(n4283), .Q(n_T_427[1928]), 
        .QN(n3557) );
  DFFX1_LVT u_T_427_reg_0__47_ ( .D(n4446), .CLK(n4282), .Q(n_T_427[1927]), 
        .QN(n3556) );
  DFFX1_LVT u_T_427_reg_0__40_ ( .D(n4425), .CLK(n4282), .Q(n_T_427[1920]), 
        .QN(n3551) );
  DFFX1_LVT u_T_427_reg_0__37_ ( .D(n4417), .CLK(n4282), .Q(n_T_427[1917]), 
        .QN(n3550) );
  DFFX1_LVT u_T_427_reg_3__17_ ( .D(n4365), .CLK(n4262), .Q(n_T_427[1744]), 
        .QN(n3541) );
  DFFX1_LVT u_T_427_reg_0__17_ ( .D(n4365), .CLK(n4280), .Q(n_T_427[1898]), 
        .QN(n3540) );
  DFFX1_LVT u_T_427_reg_0__15_ ( .D(n4360), .CLK(n4280), .Q(n_T_427[1896]), 
        .QN(n3539) );
  DFFX1_LVT u_T_427_reg_0__13_ ( .D(n4355), .CLK(n4280), .Q(n_T_427[1894]), 
        .QN(n3538) );
  DFFX1_LVT u_T_427_reg_0__12_ ( .D(n4352), .CLK(n4280), .Q(n_T_427[1893]), 
        .QN(n3537) );
  DFFX1_LVT u_T_427_reg_0__10_ ( .D(n4346), .CLK(n4279), .Q(n_T_427[1891]), 
        .QN(n3536) );
  DFFX1_LVT u_T_427_reg_0__9_ ( .D(n4343), .CLK(n4279), .Q(n_T_427[1890]), 
        .QN(n3535) );
  DFFX1_LVT u_T_427_reg_0__8_ ( .D(n4340), .CLK(n4279), .Q(n_T_427[1889]), 
        .QN(n3534) );
  DFFX1_LVT u_T_427_reg_0__7_ ( .D(n4337), .CLK(n4279), .Q(n_T_427[1888]), 
        .QN(n3533) );
  DFFX1_LVT u_T_427_reg_0__6_ ( .D(n4334), .CLK(n4279), .Q(n_T_427[1887]), 
        .QN(n3532) );
  DFFX1_LVT u_T_427_reg_0__3_ ( .D(n4325), .CLK(n4279), .QN(n3531) );
  DFFX1_LVT u_T_427_reg_0__1_ ( .D(n4319), .CLK(n4279), .Q(n_T_427[1883]), 
        .QN(n3530) );
  DFFX1_LVT u_T_427_reg_4__59_ ( .D(n4482), .CLK(n4259), .Q(n_T_427[1722]), 
        .QN(n3518) );
  DFFX1_LVT u_T_427_reg_3__59_ ( .D(n4482), .CLK(n4265), .Q(n_T_427[1786]), 
        .QN(n3517) );
  DFFX1_LVT u_T_427_reg_3__57_ ( .D(n4476), .CLK(n4265), .Q(n_T_427[1784]), 
        .QN(n3515) );
  DFFX1_LVT u_T_427_reg_4__55_ ( .D(n4470), .CLK(n4259), .Q(n_T_427[1718]), 
        .QN(n3513) );
  DFFX1_LVT u_T_427_reg_3__55_ ( .D(n4470), .CLK(n4265), .Q(n_T_427[1782]), 
        .QN(n3512) );
  DFFX1_LVT u_T_427_reg_3__53_ ( .D(n4464), .CLK(n4265), .Q(n_T_427[1780]), 
        .QN(n3510) );
  DFFX1_LVT u_T_427_reg_3__50_ ( .D(n4455), .CLK(n4265), .Q(n_T_427[1777]), 
        .QN(n3507) );
  DFFX1_LVT u_T_427_reg_3__48_ ( .D(n4449), .CLK(n4265), .Q(n_T_427[1775]), 
        .QN(n3505) );
  DFFX1_LVT u_T_427_reg_3__47_ ( .D(n4446), .CLK(n4264), .Q(n_T_427[1774]), 
        .QN(n3504) );
  DFFX1_LVT u_T_427_reg_3__40_ ( .D(n4425), .CLK(n4264), .Q(n_T_427[1767]), 
        .QN(n3499) );
  DFFX1_LVT u_T_427_reg_3__37_ ( .D(n4417), .CLK(n4264), .Q(n_T_427[1764]), 
        .QN(n3498) );
  DFFX1_LVT u_T_427_reg_4__32_ ( .D(n4404), .CLK(n4257), .Q(n_T_427[1695]), 
        .QN(n3496) );
  DFFX1_LVT u_T_427_reg_3__32_ ( .D(n4404), .CLK(n4263), .Q(n_T_427[1759]), 
        .QN(n3495) );
  DFFX1_LVT u_T_427_reg_4__17_ ( .D(n4365), .CLK(n4256), .Q(n_T_427[1680]), 
        .QN(n3494) );
  DFFX1_LVT u_T_427_reg_0__59_ ( .D(n4482), .CLK(n4283), .Q(n_T_427[1938]), 
        .QN(n3493) );
  DFFX1_LVT u_T_427_reg_0__57_ ( .D(n4476), .CLK(n4283), .Q(n_T_427[1936]), 
        .QN(n3491) );
  DFFX1_LVT u_T_427_reg_20__47_ ( .D(n4447), .CLK(n4162), .Q(n_T_427[687]), 
        .QN(n3482) );
  DFFX1_LVT u_T_427_reg_1__38_ ( .D(n4420), .CLK(n4276), .Q(n_T_427[1877]), 
        .QN(n3481) );
  DFFX1_LVT u_T_427_reg_1__35_ ( .D(n4412), .CLK(n4275), .Q(n_T_427[1876]), 
        .QN(n3480) );
  DFFX1_LVT u_T_427_reg_1__33_ ( .D(n4407), .CLK(n4275), .Q(n_T_427[1874]), 
        .QN(n3479) );
  DFFX1_LVT u_T_427_reg_1__31_ ( .D(n4402), .CLK(n4275), .Q(n_T_427[1873]), 
        .QN(n3376) );
  DFFX1_LVT u_T_427_reg_1__28_ ( .D(n4394), .CLK(n4275), .Q(n_T_427[1871]), 
        .QN(n3374) );
  DFFX1_LVT u_T_427_reg_1__26_ ( .D(n4389), .CLK(n4275), .Q(n_T_427[1869]), 
        .QN(n3373) );
  DFFX1_LVT u_T_427_reg_1__25_ ( .D(n4387), .CLK(n4275), .Q(n_T_427[1868]), 
        .QN(n3372) );
  DFFX1_LVT u_T_427_reg_1__22_ ( .D(n4379), .CLK(n4274), .QN(n3371) );
  DFFX1_LVT u_T_427_reg_1__21_ ( .D(n4377), .CLK(n4274), .Q(n_T_427[1866]), 
        .QN(n3370) );
  DFFX1_LVT u_T_427_reg_4__38_ ( .D(n4420), .CLK(n4258), .Q(n_T_427[1701]), 
        .QN(n3685) );
  DFFX1_LVT u_T_427_reg_4__33_ ( .D(n4407), .CLK(n4257), .Q(n_T_427[1696]), 
        .QN(n3655) );
  DFFX1_LVT u_T_427_reg_2__47_ ( .D(n4446), .CLK(n4270), .Q(n_T_427[1835]), 
        .QN(n3477) );
  DFFX1_LVT u_T_427_reg_2__50_ ( .D(n4455), .CLK(n4271), .Q(n_T_427[1838]), 
        .QN(n3476) );
  DFFX1_LVT u_T_427_reg_2__57_ ( .D(n4476), .CLK(n4271), .Q(n_T_427[1844]), 
        .QN(n3473) );
  DFFX1_LVT u_T_427_reg_2__53_ ( .D(n4464), .CLK(n4271), .Q(n_T_427[1841]), 
        .QN(n3470) );
  DFFX1_LVT u_T_427_reg_2__46_ ( .D(n4443), .CLK(n4270), .Q(n_T_427[1834]), 
        .QN(n3467) );
  DFFX1_LVT u_T_427_reg_1__46_ ( .D(n4443), .CLK(n4276), .Q(n_T_427[1880]), 
        .QN(n3466) );
  DFFX1_LVT u_T_427_reg_1__44_ ( .D(n4437), .CLK(n4276), .Q(n_T_427[1879]), 
        .QN(n3465) );
  DFFX1_LVT u_T_427_reg_19__40_ ( .D(n4426), .CLK(n4168), .Q(n_T_427[743]), 
        .QN(n3461) );
  DFFX1_LVT u_T_427_reg_2__40_ ( .D(n4425), .CLK(n4270), .Q(n_T_427[1828]), 
        .QN(n3460) );
  DFFX1_LVT u_T_427_reg_7__39_ ( .D(n4422), .CLK(n4240), .Q(n_T_427[1510]), 
        .QN(n3459) );
  DFFX1_LVT u_T_427_reg_2__39_ ( .D(n4422), .CLK(n4270), .Q(n_T_427[1827]), 
        .QN(n3458) );
  DFFX1_LVT u_T_427_reg_1__39_ ( .D(n4422), .CLK(n4276), .Q(n_T_427[1878]), 
        .QN(n3457) );
  DFFX1_LVT u_T_427_reg_2__37_ ( .D(n4417), .CLK(n4270), .Q(n_T_427[1825]), 
        .QN(n3456) );
  DFFX1_LVT u_T_427_reg_2__34_ ( .D(n4409), .CLK(n4269), .Q(n_T_427[1822]), 
        .QN(n3453) );
  DFFX1_LVT u_T_427_reg_1__34_ ( .D(n4409), .CLK(n4275), .Q(n_T_427[1875]), 
        .QN(n3452) );
  DFFX1_LVT u_T_427_reg_2__23_ ( .D(n4381), .CLK(n4268), .Q(n_T_427[1812]), 
        .QN(n3448) );
  DFFX1_LVT u_T_427_reg_2__16_ ( .D(n4362), .CLK(n4268), .Q(n_T_427[1806]), 
        .QN(n3444) );
  DFFX1_LVT u_T_427_reg_12__15_ ( .D(n4360), .CLK(n4208), .Q(n_T_427[1166]), 
        .QN(n3443) );
  DFFX1_LVT u_T_427_reg_7__15_ ( .D(n4360), .CLK(n4238), .Q(n_T_427[1486]), 
        .QN(n3442) );
  DFFX1_LVT u_T_427_reg_12__14_ ( .D(n4358), .CLK(n4208), .Q(n_T_427[1165]), 
        .QN(n3441) );
  DFFX1_LVT u_T_427_reg_7__14_ ( .D(n4357), .CLK(n4238), .Q(n_T_427[1485]), 
        .QN(n3440) );
  DFFX1_LVT u_T_427_reg_12__13_ ( .D(n4355), .CLK(n4208), .Q(n_T_427[1164]), 
        .QN(n3439) );
  DFFX1_LVT u_T_427_reg_7__13_ ( .D(n4355), .CLK(n4238), .Q(n_T_427[1484]), 
        .QN(n3438) );
  DFFX1_LVT u_T_427_reg_12__12_ ( .D(n4353), .CLK(n4208), .Q(n_T_427[1163]), 
        .QN(n3437) );
  DFFX1_LVT u_T_427_reg_7__12_ ( .D(n4352), .CLK(n4238), .Q(n_T_427[1483]), 
        .QN(n3436) );
  DFFX1_LVT u_T_427_reg_12__10_ ( .D(n4347), .CLK(n4207), .Q(n_T_427[1161]), 
        .QN(n3434) );
  DFFX1_LVT u_T_427_reg_7__10_ ( .D(n4346), .CLK(n4237), .Q(n_T_427[1481]), 
        .QN(n3433) );
  DFFX1_LVT u_T_427_reg_12__9_ ( .D(n4344), .CLK(n4207), .Q(n_T_427[1160]), 
        .QN(n3432) );
  DFFX1_LVT u_T_427_reg_7__9_ ( .D(n4343), .CLK(n4237), .Q(n_T_427[1480]), 
        .QN(n3431) );
  DFFX1_LVT u_T_427_reg_12__8_ ( .D(n4341), .CLK(n4207), .Q(n_T_427[1159]), 
        .QN(n3430) );
  DFFX1_LVT u_T_427_reg_7__8_ ( .D(n4340), .CLK(n4237), .Q(n_T_427[1479]), 
        .QN(n3429) );
  DFFX1_LVT u_T_427_reg_12__7_ ( .D(n4338), .CLK(n4207), .Q(n_T_427[1158]), 
        .QN(n3428) );
  DFFX1_LVT u_T_427_reg_7__7_ ( .D(n4337), .CLK(n4237), .Q(n_T_427[1478]), 
        .QN(n3427) );
  DFFX1_LVT u_T_427_reg_12__6_ ( .D(n4335), .CLK(n4207), .Q(n_T_427[1157]), 
        .QN(n3426) );
  DFFX1_LVT u_T_427_reg_7__6_ ( .D(n4334), .CLK(n4237), .Q(n_T_427[1477]), 
        .QN(n3425) );
  DFFX1_LVT u_T_427_reg_12__5_ ( .D(n4332), .CLK(n4207), .Q(n_T_427[1156]), 
        .QN(n3424) );
  DFFX1_LVT u_T_427_reg_7__5_ ( .D(n4331), .CLK(n4237), .Q(n_T_427[1476]), 
        .QN(n3423) );
  DFFX1_LVT u_T_427_reg_12__4_ ( .D(n4329), .CLK(n4207), .Q(n_T_427[1155]) );
  DFFX1_LVT u_T_427_reg_7__4_ ( .D(n4328), .CLK(n4237), .Q(n_T_427[1475]), 
        .QN(n3422) );
  DFFX1_LVT u_T_427_reg_12__3_ ( .D(n4326), .CLK(n4207), .Q(n_T_427[1154]), 
        .QN(n3421) );
  DFFX1_LVT u_T_427_reg_7__3_ ( .D(n4325), .CLK(n4237), .Q(n_T_427[1474]), 
        .QN(n3420) );
  DFFX1_LVT u_T_427_reg_12__2_ ( .D(n4323), .CLK(n4207), .Q(n_T_427[1153]), 
        .QN(n3419) );
  DFFX1_LVT u_T_427_reg_7__2_ ( .D(n4322), .CLK(n4237), .Q(n_T_427[1473]), 
        .QN(n3418) );
  DFFX1_LVT u_T_427_reg_2__44_ ( .D(n4437), .CLK(n4270), .Q(n_T_427[1832]), 
        .QN(n3415) );
  DFFX1_LVT u_T_427_reg_2__48_ ( .D(n4449), .CLK(n4271), .Q(n_T_427[1836]), 
        .QN(n3414) );
  DFFX1_LVT u_T_427_reg_14__59_ ( .D(n4483), .CLK(n4199), .Q(n_T_427[1082]), 
        .QN(n3368) );
  DFFX1_LVT u_T_427_reg_12__59_ ( .D(n4483), .CLK(n4211), .Q(n_T_427[1210]), 
        .QN(n3367) );
  DFFX1_LVT u_T_427_reg_14__57_ ( .D(n4477), .CLK(n4199), .Q(n_T_427[1080]), 
        .QN(n3364) );
  DFFX1_LVT u_T_427_reg_12__57_ ( .D(n4477), .CLK(n4211), .Q(n_T_427[1208]), 
        .QN(n3363) );
  DFFX1_LVT u_T_427_reg_12__55_ ( .D(n4471), .CLK(n4211), .Q(n_T_427[1206]), 
        .QN(n3361) );
  DFFX1_LVT u_T_427_reg_12__53_ ( .D(n4465), .CLK(n4211), .Q(n_T_427[1204]), 
        .QN(n3358) );
  DFFX1_LVT u_T_427_reg_14__53_ ( .D(n4465), .CLK(n4199), .Q(n_T_427[1076]), 
        .QN(n3357) );
  DFFX1_LVT u_T_427_reg_12__50_ ( .D(n4456), .CLK(n4211), .Q(n_T_427[1201]), 
        .QN(n3352) );
  DFFX1_LVT u_T_427_reg_14__50_ ( .D(n4456), .CLK(n4199), .Q(n_T_427[1073]), 
        .QN(n3351) );
  DFFX1_LVT u_T_427_reg_12__48_ ( .D(n4450), .CLK(n4211), .Q(n_T_427[1199]), 
        .QN(n3348) );
  DFFX1_LVT u_T_427_reg_14__47_ ( .D(n4447), .CLK(n4198), .Q(n_T_427[1070]), 
        .QN(n3347) );
  DFFX1_LVT u_T_427_reg_12__47_ ( .D(n4447), .CLK(n4210), .Q(n_T_427[1198]), 
        .QN(n3346) );
  DFFX1_LVT u_T_427_reg_12__46_ ( .D(n4444), .CLK(n4210), .Q(n_T_427[1197]), 
        .QN(n3345) );
  DFFX1_LVT u_T_427_reg_12__44_ ( .D(n4438), .CLK(n4210), .Q(n_T_427[1195]), 
        .QN(n3342) );
  DFFX1_LVT u_T_427_reg_14__40_ ( .D(n4426), .CLK(n4198), .Q(n_T_427[1063]), 
        .QN(n3338) );
  DFFX1_LVT u_T_427_reg_12__40_ ( .D(n4426), .CLK(n4210), .Q(n_T_427[1191]), 
        .QN(n3337) );
  DFFX1_LVT u_T_427_reg_12__37_ ( .D(n4418), .CLK(n4210), .Q(n_T_427[1188]), 
        .QN(n3336) );
  DFFX1_LVT u_T_427_reg_12__34_ ( .D(n4410), .CLK(n4209), .Q(n_T_427[1185]), 
        .QN(n3335) );
  DFFX1_LVT u_T_427_reg_12__32_ ( .D(n4405), .CLK(n4209), .Q(n_T_427[1183]), 
        .QN(n3334) );
  DFFX1_LVT u_T_427_reg_14__32_ ( .D(n4405), .CLK(n4197), .Q(n_T_427[1055]), 
        .QN(n3333) );
  DFFX1_LVT u_T_427_reg_1__23_ ( .D(n4381), .CLK(n4274), .Q(n_T_427[1867]), 
        .QN(n3325) );
  DFFX1_LVT u_T_427_reg_14__23_ ( .D(n4382), .CLK(n4196), .Q(n_T_427[1046]), 
        .QN(n3324) );
  DFFX1_LVT u_T_427_reg_12__23_ ( .D(n4382), .CLK(n4208), .Q(n_T_427[1174]), 
        .QN(n3323) );
  DFFX1_LVT u_T_427_reg_12__17_ ( .D(n4366), .CLK(n4208), .Q(n_T_427[1168]), 
        .QN(n3313) );
  DFFX1_LVT u_T_427_reg_12__16_ ( .D(n4363), .CLK(n4208), .Q(n_T_427[1167]), 
        .QN(n3312) );
  DFFX1_LVT u_T_427_reg_20__39_ ( .D(n4423), .CLK(n4162), .Q(n_T_427[679]), 
        .QN(n3179) );
  DFFX1_LVT u_T_427_reg_0__16_ ( .D(n4362), .CLK(n4280), .Q(n_T_427[1897]), 
        .QN(n3524) );
  DFFX1_LVT u_T_427_reg_19__50_ ( .D(n4456), .CLK(n4169), .Q(n_T_427[753]), 
        .QN(n3407) );
  DFFX1_LVT u_T_427_reg_19__46_ ( .D(n4444), .CLK(n4168), .Q(n_T_427[749]), 
        .QN(n3406) );
  DFFX1_LVT u_T_427_reg_7__38_ ( .D(n4420), .CLK(n4240), .Q(n_T_427[1509]), 
        .QN(n3403) );
  DFFX1_LVT u_T_427_reg_2__38_ ( .D(n4420), .CLK(n4270), .Q(n_T_427[1826]), 
        .QN(n3402) );
  DFFX1_LVT u_T_427_reg_2__35_ ( .D(n4412), .CLK(n4269), .Q(n_T_427[1823]), 
        .QN(n3401) );
  DFFX1_LVT u_T_427_reg_19__35_ ( .D(n4412), .CLK(n4167), .Q(n_T_427[738]), 
        .QN(n3400) );
  DFFX1_LVT u_T_427_reg_2__33_ ( .D(n4407), .CLK(n4269), .Q(n_T_427[1821]), 
        .QN(n3399) );
  DFFX1_LVT u_T_427_reg_19__32_ ( .D(n4405), .CLK(n4167), .Q(n_T_427[736]), 
        .QN(n3398) );
  DFFX1_LVT u_T_427_reg_2__31_ ( .D(n4402), .CLK(n4269), .Q(n_T_427[1820]), 
        .QN(n3397) );
  DFFX1_LVT u_T_427_reg_2__28_ ( .D(n4394), .CLK(n4269), .Q(n_T_427[1817]), 
        .QN(n3395) );
  DFFX1_LVT u_T_427_reg_2__26_ ( .D(n4389), .CLK(n4269), .Q(n_T_427[1815]), 
        .QN(n3394) );
  DFFX1_LVT u_T_427_reg_2__25_ ( .D(n4387), .CLK(n4269), .Q(n_T_427[1814]), 
        .QN(n3393) );
  DFFX1_LVT u_T_427_reg_2__22_ ( .D(n4379), .CLK(n4268), .Q(n_T_427[1811]), 
        .QN(n3392) );
  DFFX1_LVT u_T_427_reg_2__21_ ( .D(n4377), .CLK(n4268), .Q(n_T_427[1810]), 
        .QN(n3391) );
  DFFX1_LVT u_T_427_reg_4__15_ ( .D(n4360), .CLK(n4256), .Q(n_T_427[1678]), 
        .QN(n3390) );
  DFFX1_LVT u_T_427_reg_4__14_ ( .D(n4357), .CLK(n4256), .Q(n_T_427[1677]), 
        .QN(n3389) );
  DFFX1_LVT u_T_427_reg_4__13_ ( .D(n4355), .CLK(n4256), .Q(n_T_427[1676]), 
        .QN(n3388) );
  DFFX1_LVT u_T_427_reg_4__12_ ( .D(n4352), .CLK(n4256), .Q(n_T_427[1675]), 
        .QN(n3387) );
  DFFX1_LVT u_T_427_reg_12__11_ ( .D(n4350), .CLK(n4207), .Q(n_T_427[1162]) );
  DFFX1_LVT u_T_427_reg_7__11_ ( .D(n4350), .CLK(n4237), .Q(n_T_427[1482]), 
        .QN(n3386) );
  DFFX1_LVT u_T_427_reg_4__10_ ( .D(n4346), .CLK(n4255), .Q(n_T_427[1673]), 
        .QN(n3385) );
  DFFX1_LVT u_T_427_reg_4__9_ ( .D(n4343), .CLK(n4255), .Q(n_T_427[1672]), 
        .QN(n3384) );
  DFFX1_LVT u_T_427_reg_4__8_ ( .D(n4340), .CLK(n4255), .Q(n_T_427[1671]), 
        .QN(n3383) );
  DFFX1_LVT u_T_427_reg_4__7_ ( .D(n4337), .CLK(n4255), .Q(n_T_427[1670]), 
        .QN(n3382) );
  DFFX1_LVT u_T_427_reg_4__6_ ( .D(n4334), .CLK(n4255), .Q(n_T_427[1669]), 
        .QN(n3381) );
  DFFX1_LVT u_T_427_reg_4__5_ ( .D(n4331), .CLK(n4255), .Q(n_T_427[1668]), 
        .QN(n3380) );
  DFFX1_LVT u_T_427_reg_4__4_ ( .D(n4328), .CLK(n4255), .Q(n_T_427[1667]), 
        .QN(n3379) );
  DFFX1_LVT u_T_427_reg_4__3_ ( .D(n4325), .CLK(n4255), .Q(n_T_427[1666]), 
        .QN(n3378) );
  DFFX1_LVT u_T_427_reg_4__2_ ( .D(n4322), .CLK(n4255), .Q(n_T_427[1665]), 
        .QN(n3377) );
  DFFX1_LVT u_T_427_reg_19__57_ ( .D(n4477), .CLK(n4169), .Q(n_T_427[760]), 
        .QN(n3302) );
  DFFX1_LVT u_T_427_reg_19__55_ ( .D(n4471), .CLK(n4169), .Q(n_T_427[758]), 
        .QN(n3301) );
  DFFX1_LVT u_T_427_reg_14__46_ ( .D(n4444), .CLK(n4198), .Q(n_T_427[1069]), 
        .QN(n3300) );
  DFFX1_LVT u_T_427_reg_12__35_ ( .D(n4412), .CLK(n4209), .Q(n_T_427[1186]), 
        .QN(n3299) );
  DFFX1_LVT u_T_427_reg_12__33_ ( .D(n4407), .CLK(n4209), .Q(n_T_427[1184]), 
        .QN(n3298) );
  DFFX1_LVT u_T_427_reg_14__31_ ( .D(n4402), .CLK(n4197), .Q(n_T_427[1054]), 
        .QN(n3297) );
  DFFX1_LVT u_T_427_reg_12__31_ ( .D(n4402), .CLK(n4209), .Q(n_T_427[1182]), 
        .QN(n3296) );
  DFFX1_LVT u_T_427_reg_14__28_ ( .D(n4394), .CLK(n4197), .Q(n_T_427[1051]), 
        .QN(n3293) );
  DFFX1_LVT u_T_427_reg_12__28_ ( .D(n4394), .CLK(n4209), .Q(n_T_427[1179]), 
        .QN(n3292) );
  DFFX1_LVT u_T_427_reg_14__26_ ( .D(n4389), .CLK(n4197), .Q(n_T_427[1049]), 
        .QN(n3291) );
  DFFX1_LVT u_T_427_reg_12__26_ ( .D(n4389), .CLK(n4209), .Q(n_T_427[1177]), 
        .QN(n3290) );
  DFFX1_LVT u_T_427_reg_14__25_ ( .D(n4387), .CLK(n4197), .Q(n_T_427[1048]), 
        .QN(n3289) );
  DFFX1_LVT u_T_427_reg_12__25_ ( .D(n4387), .CLK(n4209), .Q(n_T_427[1176]), 
        .QN(n3288) );
  DFFX1_LVT u_T_427_reg_14__22_ ( .D(n4379), .CLK(n4196), .Q(n_T_427[1045]), 
        .QN(n3287) );
  DFFX1_LVT u_T_427_reg_12__22_ ( .D(n4379), .CLK(n4208), .Q(n_T_427[1173]), 
        .QN(n3286) );
  DFFX1_LVT u_T_427_reg_14__21_ ( .D(n4377), .CLK(n4196), .Q(n_T_427[1044]), 
        .QN(n3285) );
  DFFX1_LVT u_T_427_reg_12__21_ ( .D(n4377), .CLK(n4208), .Q(n_T_427[1172]), 
        .QN(n3284) );
  DFFX1_LVT u_T_427_reg_14__17_ ( .D(n4366), .CLK(n4196), .Q(n_T_427[1040]), 
        .QN(n3283) );
  DFFX1_LVT u_T_427_reg_14__16_ ( .D(n4363), .CLK(n4196), .Q(n_T_427[1039]), 
        .QN(n3282) );
  DFFX1_LVT u_T_427_reg_20__35_ ( .D(n4413), .CLK(n4161), .Q(n_T_427[675]), 
        .QN(n3369) );
  DFFX1_LVT u_T_427_reg_20__4_ ( .D(n4329), .CLK(n4159), .Q(n_T_427[644]), 
        .QN(n3174) );
  DFFX1_LVT u_T_427_reg_20__2_ ( .D(n4323), .CLK(n4159), .Q(n_T_427[642]), 
        .QN(n3173) );
  DFFX2_LVT ex_ctrl_alu_fn_reg_2_ ( .D(N283), .CLK(n4313), .Q(alu_io_fn[2]) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_50_ ( .D(N732), .CLK(net34650), .Q(n_T_628[52]) );
  DFFX1_LVT mem_reg_sfence_reg ( .D(n2525), .CLK(clock), .Q(n326), .QN(
        mem_reg_sfence) );
  DFFX1_LVT u_T_1057_reg ( .D(n2524), .CLK(n4499), .Q(n_T_1057) );
  DFFASX1_LVT imem_might_request_reg_reg ( .D(N271), .CLK(clock), .SETB(1'b1), 
        .Q(io_imem_might_request) );
  DFFASX1_LVT wb_reg_inst_reg_8_ ( .D(n_T_849[1]), .CLK(n4311), .SETB(1'b1), 
        .Q(wb_waddr[1]), .QN(n3103) );
  OA21X1_LVT wb_reg_cause_reg_63__U2 ( .A1(mem_reg_xcpt_interrupt), .A2(
        mem_reg_xcpt), .A3(mem_reg_cause[63]), .Y(n2521) );
  DFFASX1_LVT wb_reg_cause_reg_63_ ( .D(n2521), .CLK(n4311), .SETB(1'b1), .Q(
        wb_reg_cause[63]) );
  DFFASX1_LVT mem_reg_cause_reg_63_ ( .D(n308), .CLK(net34480), .SETB(1'b1), 
        .QN(mem_reg_cause[63]) );
  OA21X1_LVT wb_reg_cause_reg_1__U2 ( .A1(n5168), .A2(n63), .A3(n1281), .Y(
        n2518) );
  DFFASX1_LVT wb_reg_cause_reg_1_ ( .D(n2518), .CLK(n4300), .SETB(1'b1), .QN(
        wb_reg_cause[1]) );
  INVX0_LVT mem_reg_slow_bypass_reg_U4 ( .A(io_dmem_req_bits_size[1]), .Y(
        n2515) );
  DFFX1_LVT mem_reg_slow_bypass_reg ( .D(n2516), .CLK(n4285), .Q(
        mem_reg_slow_bypass) );
  OA21X1_LVT mem_reg_flush_pipe_reg_U2 ( .A1(n2495), .A2(n9516), .A3(n309), 
        .Y(n2514) );
  DFFX1_LVT mem_reg_flush_pipe_reg ( .D(n2514), .CLK(n4285), .Q(n64), .QN(
        mem_reg_flush_pipe) );
  DFFSSRX1_LVT ex_reg_rvc_reg ( .D(n9430), .SETB(1'b1), .RSTB(n4497), .CLK(
        net34469), .Q(n3215), .QN(ex_reg_rvc) );
  DFFSSRX1_LVT ex_ctrl_fp_reg ( .D(1'b0), .SETB(1'b0), .RSTB(n2512), .CLK(
        n4312), .Q(n322), .QN(io_dmem_req_bits_tag[0]) );
  DFFSSRX1_LVT ex_ctrl_mem_reg ( .D(1'b0), .SETB(1'b0), .RSTB(n2510), .CLK(
        n4312), .Q(n312), .QN(ex_ctrl_mem) );
  DFFX1_LVT ex_reg_cause_reg_63_ ( .D(csr_io_interrupt), .CLK(net34640), .QN(
        n308) );
  DFFSSRX1_LVT wb_reg_valid_reg ( .D(io_dmem_s1_kill), .SETB(n9425), .RSTB(
        1'b1), .CLK(n4499), .Q(n3203), .QN(wb_reg_valid) );
  DFFSSRX1_LVT ex_ctrl_mem_cmd_reg_1_ ( .D(n9520), .SETB(n9435), .RSTB(n1853), 
        .CLK(net34469), .Q(io_dmem_req_bits_cmd[1]), .QN(n559) );
  DFFASX1_LVT ex_reg_cause_reg_3_ ( .D(n2507), .CLK(net34640), .SETB(1'b1), 
        .Q(n75) );
  DFFSSRX1_LVT u_T_1185_reg_27_ ( .D(n5310), .SETB(1'b1), .RSTB(n5309), .CLK(
        net34660), .Q(n3135), .QN(n_T_1187[27]) );
  DFFSSRX1_LVT wb_reg_flush_pipe_reg ( .D(n64), .SETB(n1829), .RSTB(1'b1), 
        .CLK(clock), .QN(wb_reg_flush_pipe) );
  DFFSSRX1_LVT ex_reg_rs_bypass_0_reg ( .D(n9412), .SETB(1'b1), .RSTB(n1262), 
        .CLK(net34469), .Q(n3101), .QN(n2493) );
  DFFSSRX1_LVT ex_ctrl_mem_cmd_reg_3_ ( .D(1'b0), .SETB(n3578), .RSTB(n5138), 
        .CLK(net34469), .Q(io_dmem_req_bits_cmd[3]), .QN(n3122) );
  DFFSSRX1_LVT ex_ctrl_sel_alu1_reg_1_ ( .D(1'b0), .SETB(n2675), .RSTB(n9100), 
        .CLK(net34469), .Q(n561) );
  DFFSSRX1_LVT mem_reg_xcpt_reg ( .D(n2501), .SETB(n98), .RSTB(n407), .CLK(
        clock), .Q(mem_reg_xcpt), .QN(n3251) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_38_ ( .D(N720), .CLK(n4083), .Q(n_T_628[40])
         );
  DFFSSRX1_LVT ex_reg_xcpt_reg ( .D(n2874), .SETB(n1431), .RSTB(1'b1), .CLK(
        n4499), .QN(n2501) );
  DFFX1_LVT ex_reg_rs_msb_0_reg_59_ ( .D(N741), .CLK(n4084), .Q(n_T_628[61])
         );
  DFFX1_LVT ex_reg_rs_msb_0_reg_32_ ( .D(N714), .CLK(n4082), .Q(n_T_628[34])
         );
  AO221X1_LVT U2645 ( .A1(1'b1), .A2(n2234), .A3(n9158), .A4(n_T_642[3]), .A5(
        n2236), .Y(alu_io_in2[3]) );
  OA221X1_LVT U2646 ( .A1(1'b0), .A2(n1628), .A3(n9090), .A4(n2238), .A5(n2239), .Y(n2241) );
  OA221X1_LVT U2647 ( .A1(1'b0), .A2(n2199), .A3(n9512), .A4(n_T_698[1]), .A5(
        n2200), .Y(n2202) );
  OA221X1_LVT U2648 ( .A1(1'b0), .A2(n2208), .A3(n_T_698[13]), .A4(n9500), 
        .A5(n2209), .Y(n2210) );
  OA221X1_LVT U2649 ( .A1(1'b0), .A2(n2196), .A3(n9488), .A4(n_T_698[23]), 
        .A5(n2210), .Y(n2211) );
  OA21X1_LVT U2650 ( .A1(n3195), .A2(n3596), .A3(n2035), .Y(n2337) );
  IBUFFX2_LVT U2651 ( .A(n9517), .Y(n9434) );
  NAND3X4_LVT U2652 ( .A1(n3078), .A2(n9519), .A3(n9434), .Y(n5072) );
  AND2X1_LVT U2653 ( .A1(n3573), .A2(n3572), .Y(n1832) );
  AND2X1_LVT U2654 ( .A1(n6914), .A2(n1832), .Y(n6965) );
  AND2X1_LVT U2655 ( .A1(n6906), .A2(n1832), .Y(n5124) );
  AND4X1_LVT U2656 ( .A1(n2623), .A2(n2624), .A3(n5161), .A4(n5162), .Y(n2170)
         );
  NAND3X0_LVT U2657 ( .A1(n5147), .A2(n5173), .A3(n1833), .Y(n5162) );
  NAND3X0_LVT U2658 ( .A1(n5145), .A2(n3079), .A3(n1834), .Y(n1833) );
  AO21X1_LVT U2659 ( .A1(n2528), .A2(n9434), .A3(n5143), .Y(n1834) );
  NAND2X0_LVT U2660 ( .A1(n2138), .A2(n1835), .Y(n5174) );
  INVX1_LVT U2661 ( .A(io_fpu_inst[28]), .Y(n1835) );
  NOR2X0_LVT U2662 ( .A1(n3783), .A2(n2139), .Y(n2138) );
  NAND3X0_LVT U2663 ( .A1(n5107), .A2(n1837), .A3(n5106), .Y(n5108) );
  OR2X1_LVT U2664 ( .A1(n1836), .A2(n1431), .Y(n9229) );
  OR2X1_LVT U2665 ( .A1(n1837), .A2(n9092), .Y(n1836) );
  AND2X1_LVT U2666 ( .A1(io_fpu_inst[5]), .A2(n9522), .Y(n1837) );
  NAND2X0_LVT U2667 ( .A1(n1838), .A2(n5173), .Y(n5135) );
  INVX1_LVT U2668 ( .A(io_fpu_inst[13]), .Y(n1838) );
  OA22X1_LVT U2669 ( .A1(n9079), .A2(n1839), .A3(n3079), .A4(n5133), .Y(n2642)
         );
  INVX1_LVT U2670 ( .A(n5173), .Y(n1839) );
  AND2X1_LVT U2671 ( .A1(n9105), .A2(n3593), .Y(n5173) );
  OA21X1_LVT U2672 ( .A1(n4504), .A2(n1840), .A3(n4506), .Y(n4512) );
  OR3X1_LVT U2673 ( .A1(n2553), .A2(n5099), .A3(n4509), .Y(n1840) );
  AOI22X1_LVT U2674 ( .A1(n2648), .A2(n2649), .A3(n5173), .A4(n2647), .Y(n2658) );
  NAND4X0_LVT U2675 ( .A1(n3723), .A2(n3724), .A3(n8914), .A4(n1841), .Y(n8924) );
  AND2X1_LVT U2676 ( .A1(n8913), .A2(n8912), .Y(n1841) );
  AND3X1_LVT U2677 ( .A1(n3590), .A2(io_fpu_inst[6]), .A3(n9529), .Y(n2649) );
  INVX0_LVT U2678 ( .A(n9113), .Y(n3582) );
  AND3X1_LVT U2679 ( .A1(n5075), .A2(io_fpu_inst[5]), .A3(n3597), .Y(n5119) );
  IBUFFX2_LVT U2680 ( .A(n3708), .Y(n3771) );
  NAND2X1_LVT U2681 ( .A1(n3771), .A2(n_T_427[763]), .Y(n8910) );
  NAND3X1_LVT U2682 ( .A1(n7105), .A2(n7104), .A3(n7103), .Y(n7106) );
  NAND3X0_LVT U2683 ( .A1(n2166), .A2(n8125), .A3(n1842), .Y(N718) );
  AND3X1_LVT U2684 ( .A1(n2165), .A2(n8126), .A3(n8124), .Y(n1842) );
  NAND3X1_LVT U2685 ( .A1(n7087), .A2(n7086), .A3(n7085), .Y(n7109) );
  AND2X1_LVT U2686 ( .A1(n2552), .A2(n3590), .Y(n5074) );
  AOI22X2_LVT U2687 ( .A1(n1844), .A2(n1843), .A3(n_T_427[1016]), .A4(n3755), 
        .Y(n1855) );
  IBUFFX2_LVT U2688 ( .A(n3364), .Y(n1843) );
  IBUFFX2_LVT U2689 ( .A(n4013), .Y(n1844) );
  NAND2X1_LVT U2690 ( .A1(n2882), .A2(n_T_427[1916]), .Y(n8046) );
  NAND3X1_LVT U2691 ( .A1(n7083), .A2(n7082), .A3(n7081), .Y(n7110) );
  NAND2X4_LVT U2692 ( .A1(n9105), .A2(n3593), .Y(n3039) );
  NAND4X1_LVT U2693 ( .A1(n8312), .A2(n8310), .A3(n8311), .A4(n2608), .Y(n8313) );
  NOR2X0_LVT U2694 ( .A1(n8314), .A2(n8313), .Y(n3035) );
  NAND3X0_LVT U2695 ( .A1(n8051), .A2(n8049), .A3(n8050), .Y(n8080) );
  OA21X1_LVT U2696 ( .A1(n2657), .A2(n2637), .A3(n2633), .Y(n5110) );
  NAND2X0_LVT U2697 ( .A1(n2169), .A2(n2170), .Y(n2144) );
  NAND4X0_LVT U2698 ( .A1(n2894), .A2(n1892), .A3(n2893), .A4(n1845), .Y(N689)
         );
  AND3X1_LVT U2699 ( .A1(n2937), .A2(n1900), .A3(n1846), .Y(n1845) );
  AND2X1_LVT U2700 ( .A1(n7245), .A2(n7244), .Y(n1846) );
  NAND2X0_LVT U2701 ( .A1(n_T_427[1650]), .A2(n3652), .Y(n8596) );
  AND2X1_LVT U2702 ( .A1(n2933), .A2(n2934), .Y(n1888) );
  NAND2X0_LVT U2703 ( .A1(n_T_427[1662]), .A2(n3643), .Y(n9023) );
  NBUFFX2_LVT U2704 ( .A(n5116), .Y(n1847) );
  NAND2X0_LVT U2705 ( .A1(n_T_427[810]), .A2(n9056), .Y(n8323) );
  NAND2X0_LVT U2706 ( .A1(n_T_427[826]), .A2(n9056), .Y(n8884) );
  IBUFFX32_LVT U2707 ( .A(n3137), .Y(n1848) );
  NAND2X0_LVT U2708 ( .A1(n1848), .A2(n3692), .Y(n3569) );
  NAND2X0_LVT U2709 ( .A1(n_T_427[1400]), .A2(n3610), .Y(n8781) );
  IBUFFX2_LVT U2710 ( .A(n9095), .Y(n2570) );
  NAND3X4_LVT U2711 ( .A1(n5101), .A2(n2570), .A3(n9097), .Y(n5104) );
  AND2X1_LVT U2712 ( .A1(n2561), .A2(n3765), .Y(n3772) );
  AND3X1_LVT U2713 ( .A1(n4511), .A2(n4513), .A3(n4512), .Y(n9432) );
  NAND4X0_LVT U2714 ( .A1(n2917), .A2(n2916), .A3(n2958), .A4(n1849), .Y(N693)
         );
  AND2X1_LVT U2715 ( .A1(n2959), .A2(n2960), .Y(n1849) );
  AND2X4_LVT U2716 ( .A1(n7911), .A2(n7910), .Y(n8105) );
  IBUFFX2_LVT U2717 ( .A(n2984), .Y(n4013) );
  IBUFFX4_LVT U2718 ( .A(n4013), .Y(n1875) );
  OA21X1_LVT U2719 ( .A1(n3163), .A2(n3987), .A3(n8781), .Y(n8784) );
  NOR2X0_LVT U2720 ( .A1(io_fpu_inst[6]), .A2(n3590), .Y(n5164) );
  AND3X1_LVT U2721 ( .A1(n8896), .A2(n8894), .A3(n1850), .Y(n8899) );
  OA21X1_LVT U2722 ( .A1(n3409), .A2(n2969), .A3(n8895), .Y(n1850) );
  NAND2X0_LVT U2723 ( .A1(n9529), .A2(n5071), .Y(n4504) );
  AND2X1_LVT U2724 ( .A1(n3590), .A2(n9524), .Y(n5071) );
  AND3X1_LVT U2725 ( .A1(n8590), .A2(n8589), .A3(n1851), .Y(n3725) );
  AOI22X1_LVT U2726 ( .A1(n_T_427[1010]), .A2(n3759), .A3(n1875), .A4(n1884), 
        .Y(n1851) );
  NAND3X0_LVT U2727 ( .A1(n2571), .A2(n3587), .A3(n1852), .Y(n4500) );
  AND3X1_LVT U2728 ( .A1(n3590), .A2(n9445), .A3(n9435), .Y(n1852) );
  NBUFFX2_LVT U2729 ( .A(n3077), .Y(n1853) );
  NBUFFX2_LVT U2730 ( .A(n3078), .Y(io_fpu_inst[30]) );
  NAND3X2_LVT U2731 ( .A1(n3773), .A2(n6954), .A3(n2068), .Y(n9014) );
  NAND3X0_LVT U2732 ( .A1(n8796), .A2(n8795), .A3(n1855), .Y(n8797) );
  NAND3X0_LVT U2733 ( .A1(n8194), .A2(n8195), .A3(n1856), .Y(n8196) );
  OA21X1_LVT U2734 ( .A1(n3460), .A2(n3751), .A3(n8193), .Y(n1856) );
  NBUFFX2_LVT U2735 ( .A(n3076), .Y(io_fpu_inst[3]) );
  NOR4X1_LVT U2736 ( .A1(n8797), .A2(n8789), .A3(n8790), .A4(n8798), .Y(n2365)
         );
  NAND4X1_LVT U2737 ( .A1(n9061), .A2(n9060), .A3(n2619), .A4(n9057), .Y(n2600) );
  NOR3X2_LVT U2738 ( .A1(n2600), .A2(n9063), .A3(n9062), .Y(n3750) );
  NAND3X2_LVT U2739 ( .A1(n5109), .A2(n5110), .A3(n9432), .Y(n6906) );
  AND2X1_LVT U2740 ( .A1(n3593), .A2(io_fpu_inst[4]), .Y(n3597) );
  OR3X1_LVT U2741 ( .A1(n7106), .A2(n1858), .A3(n7107), .Y(n7108) );
  NAND4X0_LVT U2742 ( .A1(n7102), .A2(n2587), .A3(n2588), .A4(n7101), .Y(n1858) );
  NBUFFX2_LVT U2743 ( .A(ibuf_io_inst_0_bits_raw[30]), .Y(n1859) );
  IBUFFX2_LVT U2744 ( .A(io_fpu_inst[31]), .Y(n2139) );
  AOI22X2_LVT U2745 ( .A1(n1861), .A2(n1860), .A3(n3606), .A4(n_T_427[1379]), 
        .Y(n8054) );
  IBUFFX2_LVT U2746 ( .A(n9006), .Y(n1860) );
  IBUFFX2_LVT U2747 ( .A(n3145), .Y(n1861) );
  AND3X1_LVT U2748 ( .A1(n4510), .A2(n2620), .A3(n5149), .Y(n2145) );
  NAND2X0_LVT U2749 ( .A1(n3582), .A2(n1862), .Y(n4506) );
  AND2X1_LVT U2750 ( .A1(n4505), .A2(n5086), .Y(n1862) );
  NBUFFX2_LVT U2751 ( .A(n2553), .Y(n1863) );
  AND3X2_LVT U2752 ( .A1(n2988), .A2(n2989), .A3(n8946), .Y(n1883) );
  NAND4X1_LVT U2753 ( .A1(n3634), .A2(n1883), .A3(n2530), .A4(n2987), .Y(N741)
         );
  IBUFFX32_LVT U2754 ( .A(n_T_427[1187]), .Y(n1864) );
  OR2X1_LVT U2755 ( .A1(n3663), .A2(n1864), .Y(n8076) );
  IBUFFX2_LVT U2756 ( .A(n3783), .Y(n2553) );
  NAND3X0_LVT U2757 ( .A1(n3766), .A2(n2925), .A3(n1865), .Y(N714) );
  AND3X1_LVT U2758 ( .A1(n3762), .A2(n2923), .A3(n2924), .Y(n1865) );
  AND3X1_LVT U2759 ( .A1(n2911), .A2(n8729), .A3(n1866), .Y(n2581) );
  AND2X1_LVT U2760 ( .A1(n8727), .A2(n8728), .Y(n1866) );
  IBUFFX2_LVT U2761 ( .A(n3692), .Y(n3987) );
  NAND2X0_LVT U2762 ( .A1(n2602), .A2(n8220), .Y(n2601) );
  OA22X1_LVT U2763 ( .A1(n2641), .A2(n2642), .A3(n5158), .A4(n5141), .Y(n2623)
         );
  NBUFFX2_LVT U2764 ( .A(n9104), .Y(n1867) );
  NAND2X0_LVT U2765 ( .A1(n8848), .A2(n1868), .Y(n2147) );
  NAND2X0_LVT U2766 ( .A1(n_T_427[825]), .A2(n9056), .Y(n1868) );
  NBUFFX2_LVT U2767 ( .A(n9022), .Y(n3643) );
  AND3X1_LVT U2768 ( .A1(n6966), .A2(n6965), .A3(n2548), .Y(n7911) );
  NBUFFX2_LVT U2769 ( .A(n9022), .Y(n3649) );
  NAND2X0_LVT U2770 ( .A1(n_T_427[228]), .A2(n3745), .Y(n8048) );
  NOR2X0_LVT U2771 ( .A1(n1869), .A2(n7974), .Y(n2129) );
  NAND3X0_LVT U2772 ( .A1(n7971), .A2(n7973), .A3(n7972), .Y(n1869) );
  AND2X1_LVT U2773 ( .A1(n7248), .A2(n1870), .Y(n1893) );
  NAND2X0_LVT U2774 ( .A1(n_T_427[1352]), .A2(n3603), .Y(n1870) );
  NAND2X0_LVT U2775 ( .A1(n_T_427[1717]), .A2(n3689), .Y(n8697) );
  AOI22X1_LVT U2776 ( .A1(n1872), .A2(n1871), .A3(n3628), .A4(n_T_427[1420]), 
        .Y(n7360) );
  INVX1_LVT U2777 ( .A(n2090), .Y(n1871) );
  INVX1_LVT U2778 ( .A(n3092), .Y(n1872) );
  NAND3X0_LVT U2779 ( .A1(n2884), .A2(n2898), .A3(n1873), .Y(N672) );
  AND3X1_LVT U2780 ( .A1(n2883), .A2(n2900), .A3(n2899), .Y(n1873) );
  NAND3X1_LVT U2781 ( .A1(n5075), .A2(io_fpu_inst[5]), .A3(n3597), .Y(n5076)
         );
  NAND2X0_LVT U2782 ( .A1(n_T_427[1647]), .A2(n3643), .Y(n8493) );
  AOI22X2_LVT U2783 ( .A1(n1875), .A2(n1874), .A3(n3761), .A4(n_T_427[989]), 
        .Y(n7859) );
  IBUFFX2_LVT U2784 ( .A(n3332), .Y(n1874) );
  NAND2X0_LVT U2785 ( .A1(n_T_427[298]), .A2(n3789), .Y(n8289) );
  NOR3X0_LVT U2786 ( .A1(n3076), .A2(n9111), .A3(io_fpu_inst[11]), .Y(n4503)
         );
  NAND2X0_LVT U2787 ( .A1(n_T_427[1657]), .A2(n3649), .Y(n8829) );
  NBUFFX2_LVT U2788 ( .A(n9522), .Y(io_fpu_inst[25]) );
  NAND4X0_LVT U2789 ( .A1(n2892), .A2(n2584), .A3(n2891), .A4(n1877), .Y(N690)
         );
  AND2X1_LVT U2790 ( .A1(n7273), .A2(n2936), .Y(n1877) );
  NAND3X0_LVT U2791 ( .A1(n2905), .A2(n2971), .A3(n1878), .Y(N694) );
  AND3X1_LVT U2792 ( .A1(n2970), .A2(n2972), .A3(n2904), .Y(n1878) );
  NAND2X0_LVT U2793 ( .A1(n5119), .A2(n1879), .Y(n5111) );
  AND2X1_LVT U2794 ( .A1(n9089), .A2(csr_io_decode_0_write_illegal), .Y(n1879)
         );
  NAND4X0_LVT U2795 ( .A1(n3008), .A2(n3071), .A3(n3007), .A4(n1880), .Y(N698)
         );
  AND2X1_LVT U2796 ( .A1(n3070), .A2(n3069), .Y(n1880) );
  NAND3X0_LVT U2797 ( .A1(n2907), .A2(n2976), .A3(n1881), .Y(N686) );
  AND3X1_LVT U2798 ( .A1(n2975), .A2(n2906), .A3(n2977), .Y(n1881) );
  NBUFFX2_LVT U2799 ( .A(n9525), .Y(io_fpu_inst[6]) );
  NBUFFX2_LVT U2800 ( .A(n9528), .Y(n3077) );
  OR4X2_LVT U2801 ( .A1(n5099), .A2(n3077), .A3(n2537), .A4(io_fpu_inst[6]), 
        .Y(n2634) );
  IBUFFX2_LVT U2802 ( .A(n9528), .Y(n3578) );
  NAND4X0_LVT U2803 ( .A1(n8834), .A2(n8832), .A3(n8833), .A4(n1882), .Y(n8835) );
  OR2X1_LVT U2804 ( .A1(n3366), .A2(n4011), .Y(n1882) );
  AND2X1_LVT U2805 ( .A1(n3765), .A2(n6923), .Y(n2983) );
  NAND2X0_LVT U2806 ( .A1(n_T_427[1641]), .A2(n3649), .Y(n8272) );
  IBUFFX2_LVT U2807 ( .A(n3353), .Y(n1884) );
  OA21X1_LVT U2808 ( .A1(n3584), .A2(n1885), .A3(n5076), .Y(n3072) );
  AND2X1_LVT U2809 ( .A1(n9076), .A2(n3585), .Y(n1885) );
  NAND3X0_LVT U2810 ( .A1(n3014), .A2(n3694), .A3(n1886), .Y(N705) );
  AND3X1_LVT U2811 ( .A1(n3013), .A2(n3693), .A3(n3695), .Y(n1886) );
  NAND3X0_LVT U2812 ( .A1(n3016), .A2(n3699), .A3(n1887), .Y(N706) );
  AND3X1_LVT U2813 ( .A1(n3015), .A2(n3698), .A3(n3700), .Y(n1887) );
  NBUFFX2_LVT U2814 ( .A(n9528), .Y(n3076) );
  NAND4X1_LVT U2815 ( .A1(n2167), .A2(n2168), .A3(n2932), .A4(n1888), .Y(N722)
         );
  NAND4X0_LVT U2816 ( .A1(n2896), .A2(n2942), .A3(n2895), .A4(n1889), .Y(N683)
         );
  AND2X1_LVT U2817 ( .A1(n2943), .A2(n2944), .Y(n1889) );
  NAND4X0_LVT U2818 ( .A1(n2890), .A2(n2939), .A3(n2889), .A4(n1890), .Y(N692)
         );
  AND2X1_LVT U2819 ( .A1(n2941), .A2(n2940), .Y(n1890) );
  NBUFFX2_LVT U2820 ( .A(n3593), .Y(n1891) );
  AND2X1_LVT U2821 ( .A1(n2561), .A2(n6922), .Y(n3709) );
  AND3X1_LVT U2822 ( .A1(n7247), .A2(n7246), .A3(n1893), .Y(n1892) );
  OA21X1_LVT U2823 ( .A1(n3305), .A2(n1894), .A3(n8955), .Y(n8958) );
  IBUFFX4_LVT U2824 ( .A(n3768), .Y(n1894) );
  OA21X1_LVT U2825 ( .A1(n3339), .A2(n1894), .A3(n8250), .Y(n8253) );
  OA21X1_LVT U2826 ( .A1(n3346), .A2(n1894), .A3(n8446), .Y(n8449) );
  OA21X1_LVT U2827 ( .A1(n3365), .A2(n1894), .A3(n8828), .Y(n8831) );
  OA21X2_LVT U2828 ( .A1(n3349), .A2(n1894), .A3(n8510), .Y(n8513) );
  AND3X1_LVT U2829 ( .A1(n2962), .A2(n2961), .A3(n1895), .Y(n2945) );
  AND3X1_LVT U2830 ( .A1(n8480), .A2(n8479), .A3(n1896), .Y(n1895) );
  AOI22X1_LVT U2831 ( .A1(n_T_427[1135]), .A2(n3668), .A3(n3635), .A4(
        n_T_427[1263]), .Y(n1896) );
  AND4X1_LVT U2832 ( .A1(n7132), .A2(n1899), .A3(n7134), .A4(n7133), .Y(n1898)
         );
  IBUFFX32_LVT U2833 ( .A(n3424), .Y(n1897) );
  AND2X1_LVT U2834 ( .A1(n3599), .A2(n1898), .Y(n1901) );
  NAND2X0_LVT U2835 ( .A1(n1897), .A2(n3768), .Y(n1899) );
  IBUFFX4_LVT U2836 ( .A(n3768), .Y(n4010) );
  OA22X1_LVT U2837 ( .A1(n3189), .A2(n4016), .A3(n3432), .A4(n2081), .Y(n1900)
         );
  NAND4X0_LVT U2838 ( .A1(n2886), .A2(n2885), .A3(n3598), .A4(n1901), .Y(N685)
         );
  NAND2X0_LVT U2839 ( .A1(n1902), .A2(n2909), .Y(N682) );
  AND3X1_LVT U2840 ( .A1(n2978), .A2(n2908), .A3(n1903), .Y(n1902) );
  AND3X1_LVT U2841 ( .A1(n2979), .A2(n7044), .A3(n1904), .Y(n1903) );
  AND2X1_LVT U2842 ( .A1(n7046), .A2(n1905), .Y(n1904) );
  OA21X1_LVT U2843 ( .A1(n3419), .A2(n3663), .A3(n7045), .Y(n1905) );
  NAND4X0_LVT U2844 ( .A1(n3778), .A2(n1907), .A3(n2949), .A4(n1906), .Y(N721)
         );
  AND2X1_LVT U2845 ( .A1(n2948), .A2(n3754), .Y(n1906) );
  AND4X1_LVT U2846 ( .A1(n1909), .A2(n8255), .A3(n1908), .A4(n8256), .Y(n1907)
         );
  AND2X1_LVT U2847 ( .A1(n8254), .A2(n8252), .Y(n1908) );
  AND2X1_LVT U2848 ( .A1(n8251), .A2(n8253), .Y(n1909) );
  NAND4X0_LVT U2849 ( .A1(n2888), .A2(n2887), .A3(n2938), .A4(n1910), .Y(N695)
         );
  AND2X1_LVT U2850 ( .A1(n1912), .A2(n1911), .Y(n1910) );
  AND4X1_LVT U2851 ( .A1(n7411), .A2(n1913), .A3(n7414), .A4(n7412), .Y(n1911)
         );
  AND3X1_LVT U2852 ( .A1(n7416), .A2(n7415), .A3(n7413), .Y(n1912) );
  OA22X1_LVT U2853 ( .A1(n4016), .A2(n3093), .A3(n3443), .A4(n4009), .Y(n1913)
         );
  AND3X2_LVT U2854 ( .A1(n2677), .A2(io_fpu_inst[14]), .A3(n9231), .Y(n9087)
         );
  AND3X2_LVT U2855 ( .A1(n9412), .A2(n9099), .A3(n5167), .Y(n2677) );
  NAND4X0_LVT U2856 ( .A1(n4765), .A2(n6924), .A3(n4764), .A4(n4763), .Y(n4766) );
  NAND3X0_LVT U2857 ( .A1(n1914), .A2(n1915), .A3(n1916), .Y(n4852) );
  OR4X1_LVT U2858 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .Y(n1914)
         );
  OR4X1_LVT U2859 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .Y(n1915)
         );
  AND4X1_LVT U2860 ( .A1(n4780), .A2(io_fpu_dec_ren1), .A3(n4779), .A4(n9286), 
        .Y(n1916) );
  NAND4X1_LVT U2861 ( .A1(n4954), .A2(n4955), .A3(n4953), .A4(n4952), .Y(n1917) );
  NBUFFX2_LVT U2862 ( .A(n6810), .Y(n1918) );
  NBUFFX2_LVT U2863 ( .A(n6810), .Y(n1919) );
  AND2X1_LVT U2864 ( .A1(n2981), .A2(n3864), .Y(n6829) );
  OR2X2_LVT U2865 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(
        ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n4814) );
  OA22X1_LVT U2866 ( .A1(n3162), .A2(n1994), .A3(n3514), .A4(n3800), .Y(n6676)
         );
  AND4X1_LVT U2867 ( .A1(n1920), .A2(n1921), .A3(n1922), .A4(n1923), .Y(n6458)
         );
  AOI22X2_LVT U2868 ( .A1(n3829), .A2(n_T_427[1835]), .A3(n_T_427[1710]), .A4(
        n3825), .Y(n1920) );
  AOI22X2_LVT U2869 ( .A1(n3893), .A2(n_T_427[1582]), .A3(n_T_427[1646]), .A4(
        n3887), .Y(n1921) );
  AOI22X2_LVT U2870 ( .A1(n3925), .A2(n_T_427[1518]), .A3(n_T_427[1390]), .A4(
        n3919), .Y(n1922) );
  AOI22X2_LVT U2871 ( .A1(n3935), .A2(n_T_427[1454]), .A3(n_T_427[1326]), .A4(
        n3930), .Y(n1923) );
  AND4X1_LVT U2872 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .Y(n6317)
         );
  AOI22X2_LVT U2873 ( .A1(n3830), .A2(n_T_427[1829]), .A3(n_T_427[1704]), .A4(
        n3825), .Y(n1924) );
  AOI22X2_LVT U2874 ( .A1(n3892), .A2(n_T_427[1576]), .A3(n_T_427[1640]), .A4(
        n3887), .Y(n1925) );
  AOI22X2_LVT U2875 ( .A1(n3925), .A2(n_T_427[1512]), .A3(n_T_427[1384]), .A4(
        n3919), .Y(n1926) );
  AOI22X2_LVT U2876 ( .A1(n3935), .A2(n_T_427[1448]), .A3(n_T_427[1320]), .A4(
        n3929), .Y(n1927) );
  AND4X1_LVT U2877 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .Y(n6204)
         );
  AOI22X2_LVT U2878 ( .A1(n3829), .A2(n_T_427[1824]), .A3(n_T_427[1699]), .A4(
        n3825), .Y(n1928) );
  AOI22X1_LVT U2879 ( .A1(n3892), .A2(n_T_427[1571]), .A3(n_T_427[1635]), .A4(
        n3886), .Y(n1929) );
  AOI22X1_LVT U2880 ( .A1(n3924), .A2(n_T_427[1507]), .A3(n_T_427[1379]), .A4(
        n3919), .Y(n1930) );
  AOI22X1_LVT U2881 ( .A1(n3934), .A2(n_T_427[1443]), .A3(n_T_427[1315]), .A4(
        n3929), .Y(n1931) );
  AND4X1_LVT U2882 ( .A1(n1932), .A2(n1933), .A3(n1934), .A4(n1935), .Y(n6409)
         );
  AOI22X2_LVT U2883 ( .A1(n3830), .A2(n_T_427[1833]), .A3(n_T_427[1708]), .A4(
        n3825), .Y(n1932) );
  AOI22X2_LVT U2884 ( .A1(n3893), .A2(n_T_427[1580]), .A3(n_T_427[1644]), .A4(
        n3888), .Y(n1933) );
  AOI22X2_LVT U2885 ( .A1(n3925), .A2(n_T_427[1516]), .A3(n_T_427[1388]), .A4(
        n3919), .Y(n1934) );
  AOI22X2_LVT U2886 ( .A1(n3935), .A2(n_T_427[1452]), .A3(n_T_427[1324]), .A4(
        n3930), .Y(n1935) );
  AND4X1_LVT U2887 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .Y(n6363)
         );
  AOI22X2_LVT U2888 ( .A1(n3829), .A2(n_T_427[1831]), .A3(n_T_427[1706]), .A4(
        n3825), .Y(n1936) );
  AOI22X2_LVT U2889 ( .A1(n3893), .A2(n_T_427[1578]), .A3(n_T_427[1642]), .A4(
        n3887), .Y(n1937) );
  AOI22X2_LVT U2890 ( .A1(n3925), .A2(n_T_427[1514]), .A3(n_T_427[1386]), .A4(
        n3920), .Y(n1938) );
  AOI22X2_LVT U2891 ( .A1(n3935), .A2(n_T_427[1450]), .A3(n_T_427[1322]), .A4(
        n3929), .Y(n1939) );
  AND4X1_LVT U2892 ( .A1(n1940), .A2(n1941), .A3(n1942), .A4(n1943), .Y(n6225)
         );
  AOI22X2_LVT U2893 ( .A1(n3829), .A2(n_T_427[1825]), .A3(n_T_427[1700]), .A4(
        n3825), .Y(n1940) );
  AOI22X2_LVT U2894 ( .A1(n3892), .A2(n_T_427[1572]), .A3(n_T_427[1636]), .A4(
        n3887), .Y(n1941) );
  AOI22X1_LVT U2895 ( .A1(n3924), .A2(n_T_427[1508]), .A3(n_T_427[1380]), .A4(
        n3919), .Y(n1942) );
  AOI22X1_LVT U2896 ( .A1(n3934), .A2(n_T_427[1444]), .A3(n_T_427[1316]), .A4(
        n3929), .Y(n1943) );
  AOI22X1_LVT U2897 ( .A1(n3801), .A2(n_T_427[1864]), .A3(n_T_427[1746]), .A4(
        n2866), .Y(n1988) );
  AND4X1_LVT U2898 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(n1947), .Y(n6012)
         );
  AOI22X1_LVT U2899 ( .A1(n1918), .A2(n_T_427[347]), .A3(n_T_427[539]), .A4(
        n3819), .Y(n1944) );
  AOI22X1_LVT U2900 ( .A1(n3912), .A2(n_T_427[475]), .A3(n_T_427[922]), .A4(
        n3896), .Y(n1945) );
  AOI22X1_LVT U2901 ( .A1(n3914), .A2(n_T_427[27]), .A3(n_T_427[155]), .A4(
        n2863), .Y(n1946) );
  AND3X1_LVT U2902 ( .A1(n6005), .A2(n6004), .A3(n6003), .Y(n1947) );
  AND4X1_LVT U2903 ( .A1(n1948), .A2(n1949), .A3(n1950), .A4(n1951), .Y(n6532)
         );
  AOI22X1_LVT U2904 ( .A1(n2765), .A2(n_T_427[1838]), .A3(n_T_427[1713]), .A4(
        n3824), .Y(n1948) );
  AOI22X2_LVT U2905 ( .A1(n3893), .A2(n_T_427[1585]), .A3(n_T_427[1649]), .A4(
        n3887), .Y(n1949) );
  AOI22X2_LVT U2906 ( .A1(n3925), .A2(n_T_427[1521]), .A3(n_T_427[1393]), .A4(
        n3920), .Y(n1950) );
  AOI22X2_LVT U2907 ( .A1(n3935), .A2(n_T_427[1457]), .A3(n_T_427[1329]), .A4(
        n3929), .Y(n1951) );
  AND4X1_LVT U2908 ( .A1(n1952), .A2(n1953), .A3(n1954), .A4(n1955), .Y(n6609)
         );
  AOI22X1_LVT U2909 ( .A1(n2765), .A2(n_T_427[1841]), .A3(n_T_427[1716]), .A4(
        n3824), .Y(n1952) );
  AOI22X2_LVT U2910 ( .A1(n3893), .A2(n_T_427[1588]), .A3(n_T_427[1652]), .A4(
        n3888), .Y(n1953) );
  AOI22X2_LVT U2911 ( .A1(n3926), .A2(n_T_427[1524]), .A3(n_T_427[1396]), .A4(
        n3920), .Y(n1954) );
  AOI22X2_LVT U2912 ( .A1(n3936), .A2(n_T_427[1460]), .A3(n_T_427[1332]), .A4(
        n3930), .Y(n1955) );
  AND4X1_LVT U2913 ( .A1(n1956), .A2(n1957), .A3(n1958), .A4(n1959), .Y(n6702)
         );
  AOI22X1_LVT U2914 ( .A1(n2765), .A2(n_T_427[1844]), .A3(n_T_427[1720]), .A4(
        n3824), .Y(n1956) );
  AOI22X2_LVT U2915 ( .A1(n3893), .A2(n_T_427[1592]), .A3(n_T_427[1656]), .A4(
        n3888), .Y(n1957) );
  AOI22X2_LVT U2916 ( .A1(n3926), .A2(n_T_427[1528]), .A3(n_T_427[1400]), .A4(
        n3921), .Y(n1958) );
  AOI22X2_LVT U2917 ( .A1(n3936), .A2(n_T_427[1464]), .A3(n_T_427[1336]), .A4(
        n3930), .Y(n1959) );
  AND4X1_LVT U2918 ( .A1(n1960), .A2(n1961), .A3(n1962), .A4(n1963), .Y(n6850)
         );
  AOI22X1_LVT U2919 ( .A1(n2765), .A2(n_T_427[1847]), .A3(n_T_427[1725]), .A4(
        n3827), .Y(n1960) );
  AOI22X2_LVT U2920 ( .A1(n3894), .A2(n_T_427[1597]), .A3(n_T_427[1661]), .A4(
        n3888), .Y(n1961) );
  AOI22X2_LVT U2921 ( .A1(n3926), .A2(n_T_427[1533]), .A3(n_T_427[1405]), .A4(
        n3920), .Y(n1962) );
  AOI22X2_LVT U2922 ( .A1(n3936), .A2(n_T_427[1469]), .A3(n_T_427[1341]), .A4(
        n3929), .Y(n1963) );
  AND4X1_LVT U2923 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .Y(n5947)
         );
  AOI22X1_LVT U2924 ( .A1(n2765), .A2(n_T_427[1813]), .A3(n_T_427[1687]), .A4(
        n3826), .Y(n1964) );
  AOI22X2_LVT U2925 ( .A1(n3892), .A2(n_T_427[1559]), .A3(n_T_427[1623]), .A4(
        n3887), .Y(n1965) );
  AOI22X2_LVT U2926 ( .A1(n3924), .A2(n_T_427[1495]), .A3(n_T_427[1367]), .A4(
        n3918), .Y(n1966) );
  AOI22X2_LVT U2927 ( .A1(n3934), .A2(n_T_427[1431]), .A3(n_T_427[1303]), .A4(
        n3928), .Y(n1967) );
  AND4X1_LVT U2928 ( .A1(n1968), .A2(n1969), .A3(n1970), .A4(n1971), .Y(n6292)
         );
  AOI22X1_LVT U2929 ( .A1(n2765), .A2(n_T_427[1828]), .A3(n_T_427[1703]), .A4(
        n3825), .Y(n1968) );
  AOI22X2_LVT U2930 ( .A1(n3892), .A2(n_T_427[1575]), .A3(n_T_427[1639]), .A4(
        n3887), .Y(n1969) );
  AOI22X2_LVT U2931 ( .A1(n3925), .A2(n_T_427[1511]), .A3(n_T_427[1383]), .A4(
        n3919), .Y(n1970) );
  AOI22X2_LVT U2932 ( .A1(n3935), .A2(n_T_427[1447]), .A3(n_T_427[1319]), .A4(
        n3929), .Y(n1971) );
  AND4X1_LVT U2933 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .Y(n6629)
         );
  AOI22X1_LVT U2934 ( .A1(n2765), .A2(n_T_427[1842]), .A3(n_T_427[1717]), .A4(
        n3824), .Y(n1972) );
  AOI22X2_LVT U2935 ( .A1(n3893), .A2(n_T_427[1589]), .A3(n_T_427[1653]), .A4(
        n3888), .Y(n1973) );
  AOI22X2_LVT U2936 ( .A1(n3926), .A2(n_T_427[1525]), .A3(n_T_427[1397]), .A4(
        n3921), .Y(n1974) );
  AOI22X2_LVT U2937 ( .A1(n3936), .A2(n_T_427[1461]), .A3(n_T_427[1333]), .A4(
        n3930), .Y(n1975) );
  AND4X1_LVT U2938 ( .A1(n1976), .A2(n1977), .A3(n1978), .A4(n1979), .Y(n6342)
         );
  AOI22X1_LVT U2939 ( .A1(n2765), .A2(n_T_427[1830]), .A3(n_T_427[1705]), .A4(
        n3825), .Y(n1976) );
  AOI22X2_LVT U2940 ( .A1(n3893), .A2(n_T_427[1577]), .A3(n_T_427[1641]), .A4(
        n3887), .Y(n1977) );
  AOI22X2_LVT U2941 ( .A1(n3925), .A2(n_T_427[1513]), .A3(n_T_427[1385]), .A4(
        n3920), .Y(n1978) );
  AOI22X2_LVT U2942 ( .A1(n3935), .A2(n_T_427[1449]), .A3(n_T_427[1321]), .A4(
        n3929), .Y(n1979) );
  AND4X1_LVT U2943 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .Y(n5923)
         );
  AOI22X1_LVT U2944 ( .A1(n2028), .A2(n_T_427[1867]), .A3(n_T_427[1750]), .A4(
        n2868), .Y(n1980) );
  AOI22X1_LVT U2945 ( .A1(n2765), .A2(n_T_427[1812]), .A3(n_T_427[1686]), .A4(
        n3825), .Y(n1981) );
  AOI22X1_LVT U2946 ( .A1(n3891), .A2(n_T_427[1558]), .A3(n_T_427[1622]), .A4(
        n3886), .Y(n1982) );
  AOI22X2_LVT U2947 ( .A1(n5911), .A2(n6877), .A3(n_T_427[1904]), .A4(n3884), 
        .Y(n1983) );
  AND4X1_LVT U2948 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .Y(n5724)
         );
  AOI22X2_LVT U2949 ( .A1(n6764), .A2(n_T_427[1859]), .A3(n_T_427[1740]), .A4(
        n2866), .Y(n1984) );
  AOI22X2_LVT U2950 ( .A1(n3828), .A2(n_T_427[1803]), .A3(n_T_427[1676]), .A4(
        n3827), .Y(n1985) );
  AOI22X1_LVT U2951 ( .A1(n3891), .A2(n_T_427[1548]), .A3(n_T_427[1612]), .A4(
        n3885), .Y(n1986) );
  AOI22X2_LVT U2952 ( .A1(n3923), .A2(n_T_427[1484]), .A3(n_T_427[1356]), .A4(
        n3918), .Y(n1987) );
  AND4X1_LVT U2953 ( .A1(n1988), .A2(n1989), .A3(n1990), .A4(n1991), .Y(n2429)
         );
  AOI22X1_LVT U2954 ( .A1(n2765), .A2(n_T_427[1808]), .A3(n_T_427[1682]), .A4(
        n3825), .Y(n1989) );
  AOI22X2_LVT U2955 ( .A1(n3886), .A2(n_T_427[1618]), .A3(n_T_427[1554]), .A4(
        n3891), .Y(n1990) );
  AOI22X2_LVT U2956 ( .A1(n3918), .A2(n_T_427[1362]), .A3(n_T_427[1490]), .A4(
        n3924), .Y(n1991) );
  INVX1_LVT U2957 ( .A(n3586), .Y(n1992) );
  NBUFFX2_LVT U2958 ( .A(n3877), .Y(n1993) );
  AND2X1_LVT U2959 ( .A1(n5434), .A2(n6238), .Y(n2981) );
  NBUFFX2_LVT U2960 ( .A(n2875), .Y(n1994) );
  NBUFFX2_LVT U2961 ( .A(n2875), .Y(n3080) );
  AND4X1_LVT U2962 ( .A1(n1995), .A2(n1996), .A3(n1997), .A4(n1998), .Y(n6096)
         );
  AOI22X2_LVT U2963 ( .A1(n2866), .A2(n_T_427[1758]), .A3(n_T_427[1820]), .A4(
        n3830), .Y(n1995) );
  AOI22X1_LVT U2964 ( .A1(n_T_427[1873]), .A2(n3801), .A3(n3884), .A4(
        n_T_427[1912]), .Y(n1996) );
  AOI22X1_LVT U2965 ( .A1(n3826), .A2(n_T_427[1694]), .A3(n_T_427[1566]), .A4(
        n3890), .Y(n1997) );
  AOI22X1_LVT U2966 ( .A1(n3889), .A2(n_T_427[1630]), .A3(n_T_427[1502]), .A4(
        n3922), .Y(n1998) );
  AND4X1_LVT U2967 ( .A1(n1999), .A2(n2000), .A3(n2001), .A4(n2002), .Y(n5876)
         );
  AOI22X1_LVT U2968 ( .A1(n2868), .A2(n_T_427[1748]), .A3(n_T_427[1810]), .A4(
        n3829), .Y(n1999) );
  AOI22X1_LVT U2969 ( .A1(n_T_427[1866]), .A2(n6764), .A3(n3884), .A4(
        n_T_427[1902]), .Y(n2000) );
  AOI22X1_LVT U2970 ( .A1(n3827), .A2(n_T_427[1684]), .A3(n_T_427[1556]), .A4(
        n3890), .Y(n2001) );
  AOI22X2_LVT U2971 ( .A1(n3888), .A2(n_T_427[1620]), .A3(n_T_427[1492]), .A4(
        n3922), .Y(n2002) );
  AND4X1_LVT U2972 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .Y(n5991)
         );
  AOI22X2_LVT U2973 ( .A1(n2866), .A2(n_T_427[1753]), .A3(n_T_427[1815]), .A4(
        n3830), .Y(n2003) );
  AOI22X1_LVT U2974 ( .A1(n3802), .A2(n_T_427[1869]), .A3(n3884), .A4(
        n_T_427[1907]), .Y(n2004) );
  AOI22X1_LVT U2975 ( .A1(n3827), .A2(n_T_427[1689]), .A3(n_T_427[1561]), .A4(
        n3890), .Y(n2005) );
  AOI22X1_LVT U2976 ( .A1(n3889), .A2(n_T_427[1625]), .A3(n_T_427[1497]), .A4(
        n3922), .Y(n2006) );
  AND4X1_LVT U2977 ( .A1(n2007), .A2(n2008), .A3(n2009), .A4(n2010), .Y(n5763)
         );
  AOI22X1_LVT U2978 ( .A1(n3801), .A2(n_T_427[1861]), .A3(n_T_427[1742]), .A4(
        n2868), .Y(n2007) );
  AOI22X1_LVT U2979 ( .A1(n2765), .A2(n_T_427[1805]), .A3(n_T_427[1678]), .A4(
        n3824), .Y(n2008) );
  AOI22X1_LVT U2980 ( .A1(n3892), .A2(n_T_427[1550]), .A3(n_T_427[1614]), .A4(
        n3886), .Y(n2009) );
  AOI22X2_LVT U2981 ( .A1(n3924), .A2(n_T_427[1486]), .A3(n_T_427[1358]), .A4(
        n3918), .Y(n2010) );
  AND4X1_LVT U2982 ( .A1(n2011), .A2(n2012), .A3(n2013), .A4(n2014), .Y(n2290)
         );
  AOI22X2_LVT U2983 ( .A1(n2866), .A2(n_T_427[1755]), .A3(n_T_427[1817]), .A4(
        n2765), .Y(n2011) );
  AOI22X1_LVT U2984 ( .A1(n_T_427[1871]), .A2(n6764), .A3(n3884), .A4(
        n_T_427[1909]), .Y(n2012) );
  AOI22X1_LVT U2985 ( .A1(n3827), .A2(n_T_427[1691]), .A3(n_T_427[1563]), .A4(
        n3890), .Y(n2013) );
  AOI22X2_LVT U2986 ( .A1(n3922), .A2(n_T_427[1499]), .A3(n_T_427[1627]), .A4(
        n3887), .Y(n2014) );
  AND4X1_LVT U2987 ( .A1(n2015), .A2(n2016), .A3(n2017), .A4(n2018), .Y(n2229)
         );
  AOI22X1_LVT U2988 ( .A1(n3802), .A2(n_T_427[1850]), .A3(n_T_427[1731]), .A4(
        n3798), .Y(n2015) );
  AOI22X1_LVT U2989 ( .A1(n2765), .A2(n_T_427[1794]), .A3(n_T_427[1667]), .A4(
        n3826), .Y(n2016) );
  AOI22X1_LVT U2990 ( .A1(n3891), .A2(n_T_427[1539]), .A3(n_T_427[1603]), .A4(
        n3885), .Y(n2017) );
  AOI22X1_LVT U2991 ( .A1(n5534), .A2(n1992), .A3(n_T_427[1885]), .A4(n3884), 
        .Y(n2018) );
  AND4X1_LVT U2992 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .Y(n2249)
         );
  AOI22X2_LVT U2993 ( .A1(n2866), .A2(n_T_427[1765]), .A3(n_T_427[1826]), .A4(
        n2765), .Y(n2019) );
  AOI22X1_LVT U2994 ( .A1(n_T_427[1877]), .A2(n3802), .A3(n3884), .A4(
        n_T_427[1918]), .Y(n2020) );
  AOI22X1_LVT U2995 ( .A1(n3827), .A2(n_T_427[1701]), .A3(n_T_427[1573]), .A4(
        n3890), .Y(n2021) );
  AOI22X2_LVT U2996 ( .A1(n3922), .A2(n_T_427[1509]), .A3(n_T_427[1637]), .A4(
        n3889), .Y(n2022) );
  AND4X1_LVT U2997 ( .A1(n2023), .A2(n2024), .A3(n2025), .A4(n2026), .Y(n6158)
         );
  AOI22X1_LVT U2998 ( .A1(n3802), .A2(n_T_427[1875]), .A3(n_T_427[1761]), .A4(
        n2868), .Y(n2023) );
  AOI22X1_LVT U2999 ( .A1(n6146), .A2(n6877), .A3(n3884), .A4(n_T_427[1914]), 
        .Y(n2024) );
  AOI22X2_LVT U3000 ( .A1(n3829), .A2(n_T_427[1822]), .A3(n_T_427[1697]), .A4(
        n3825), .Y(n2025) );
  AOI22X1_LVT U3001 ( .A1(n3892), .A2(n_T_427[1569]), .A3(n_T_427[1633]), .A4(
        n3886), .Y(n2026) );
  NBUFFX2_LVT U3002 ( .A(n2875), .Y(n2027) );
  INVX1_LVT U3003 ( .A(n2875), .Y(n2028) );
  IBUFFX2_LVT U3004 ( .A(io_dmem_resp_bits_tag[0]), .Y(n2029) );
  NBUFFX2_LVT U3005 ( .A(io_dmem_resp_valid), .Y(n2030) );
  NAND3X0_LVT U3006 ( .A1(n9390), .A2(n2152), .A3(n2573), .Y(n9395) );
  IBUFFX2_LVT U3007 ( .A(n3883), .Y(n3881) );
  IBUFFX2_LVT U3008 ( .A(n3883), .Y(n3882) );
  AOI22X2_LVT U3009 ( .A1(n3828), .A2(n_T_427[1809]), .A3(n_T_427[1683]), .A4(
        n3827), .Y(n2800) );
  IBUFFX2_LVT U3010 ( .A(n3082), .Y(n3824) );
  IBUFFX2_LVT U3011 ( .A(n3082), .Y(n3827) );
  IBUFFX2_LVT U3012 ( .A(n4969), .Y(n4748) );
  NAND2X4_LVT U3013 ( .A1(n6238), .A2(n3579), .Y(n3803) );
  AND3X1_LVT U3014 ( .A1(n2031), .A2(n2032), .A3(n2033), .Y(n2035) );
  AOI22X1_LVT U3015 ( .A1(n3891), .A2(n_T_427[1549]), .A3(n_T_427[1613]), .A4(
        n3886), .Y(n2031) );
  AOI22X2_LVT U3016 ( .A1(n1992), .A2(n5736), .A3(n_T_427[1895]), .A4(n3884), 
        .Y(n2032) );
  AOI22X1_LVT U3017 ( .A1(n2765), .A2(n_T_427[1804]), .A3(n_T_427[1677]), .A4(
        n3826), .Y(n2033) );
  NBUFFX2_LVT U3018 ( .A(n5453), .Y(n2034) );
  AND2X1_LVT U3019 ( .A1(n4901), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5453) );
  IBUFFX2_LVT U3020 ( .A(n6898), .Y(n3596) );
  IBUFFX2_LVT U3021 ( .A(n3195), .Y(n4359) );
  AOI21X2_LVT U3022 ( .A1(n3843), .A2(csr_io_rw_rdata[14]), .A3(n5731), .Y(
        n3195) );
  AND2X4_LVT U3023 ( .A1(n4970), .A2(n4752), .Y(n6948) );
  AND2X4_LVT U3024 ( .A1(n6948), .A2(n6956), .Y(n9041) );
  AND2X4_LVT U3025 ( .A1(n6948), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n9039) );
  OR2X2_LVT U3026 ( .A1(n2877), .A2(ibuf_io_inst_0_bits_inst_rs1[0]), .Y(n4969) );
  OR2X2_LVT U3027 ( .A1(ibuf_io_inst_0_bits_inst_rs2[3]), .A2(n4880), .Y(n6423) );
  NBUFFX2_LVT U3028 ( .A(n3040), .Y(n2036) );
  AND2X4_LVT U3029 ( .A1(n2036), .A2(n2061), .Y(n9389) );
  AND2X4_LVT U3030 ( .A1(n2036), .A2(n3042), .Y(n9393) );
  IBUFFX2_LVT U3031 ( .A(n3042), .Y(n2037) );
  DELLN3X2_LVT U3032 ( .A(n2037), .Y(n2061) );
  NBUFFX2_LVT U3033 ( .A(ibuf_io_inst_0_bits_inst_rs1[2]), .Y(n2038) );
  AND2X4_LVT U3034 ( .A1(n4748), .A2(n4752), .Y(n6957) );
  AND3X1_LVT U3035 ( .A1(n2039), .A2(n2040), .A3(n2041), .Y(n2108) );
  AND4X1_LVT U3036 ( .A1(n8184), .A2(n8182), .A3(n8183), .A4(n2612), .Y(n2039)
         );
  AND2X1_LVT U3037 ( .A1(n8170), .A2(n8169), .Y(n2040) );
  AND3X1_LVT U3038 ( .A1(n8181), .A2(n8180), .A3(n8179), .Y(n2041) );
  OA21X1_LVT U3039 ( .A1(n3144), .A2(n2120), .A3(n7935), .Y(n7936) );
  AND3X1_LVT U3040 ( .A1(n2042), .A2(n2043), .A3(n2044), .Y(n3743) );
  AND3X1_LVT U3041 ( .A1(n8458), .A2(n2589), .A3(n8459), .Y(n2042) );
  AND3X1_LVT U3042 ( .A1(n8465), .A2(n8464), .A3(n8463), .Y(n2043) );
  AND2X1_LVT U3043 ( .A1(n8461), .A2(n8460), .Y(n2044) );
  OA21X1_LVT U3044 ( .A1(n3146), .A2(n3767), .A3(n8101), .Y(n8104) );
  NAND3X0_LVT U3045 ( .A1(n2045), .A2(n2046), .A3(n2047), .Y(N696) );
  AND3X1_LVT U3046 ( .A1(n2086), .A2(n2087), .A3(n2088), .Y(n2045) );
  AND3X1_LVT U3047 ( .A1(n7420), .A2(n7419), .A3(n7418), .Y(n2046) );
  AND3X1_LVT U3048 ( .A1(n7424), .A2(n7423), .A3(n7422), .Y(n2047) );
  AND2X1_LVT U3049 ( .A1(n8994), .A2(n_T_427[122]), .Y(n2149) );
  NAND3X2_LVT U3050 ( .A1(n4497), .A2(n6916), .A3(n6915), .Y(n2627) );
  AND3X1_LVT U3051 ( .A1(n2048), .A2(n2049), .A3(n2050), .Y(n2173) );
  AND4X1_LVT U3052 ( .A1(n8564), .A2(n8562), .A3(n2603), .A4(n2593), .Y(n2048)
         );
  AND3X1_LVT U3053 ( .A1(n8560), .A2(n8559), .A3(n8558), .Y(n2049) );
  AND3X1_LVT U3054 ( .A1(n8554), .A2(n8555), .A3(n8556), .Y(n2050) );
  AND2X1_LVT U3055 ( .A1(n2051), .A2(n2052), .Y(n2160) );
  AND3X1_LVT U3056 ( .A1(n8381), .A2(n8380), .A3(n8379), .Y(n2051) );
  AND3X1_LVT U3057 ( .A1(n8384), .A2(n8382), .A3(n2604), .Y(n2052) );
  AND2X1_LVT U3058 ( .A1(n2053), .A2(n2054), .Y(n2543) );
  AND3X1_LVT U3059 ( .A1(n8365), .A2(n8364), .A3(n8363), .Y(n2053) );
  AND3X1_LVT U3060 ( .A1(n8361), .A2(n8360), .A3(n8359), .Y(n2054) );
  NAND3X1_LVT U3061 ( .A1(n4497), .A2(n6915), .A3(n6916), .Y(n6962) );
  NAND3X0_LVT U3062 ( .A1(n5166), .A2(n3049), .A3(n5110), .Y(n3075) );
  AND2X1_LVT U3063 ( .A1(n1612), .A2(n3049), .Y(n2510) );
  OA21X1_LVT U3064 ( .A1(n3480), .A2(n3767), .A3(n8027), .Y(n8030) );
  AND2X1_LVT U3065 ( .A1(n2055), .A2(n2056), .Y(n2096) );
  AND3X1_LVT U3066 ( .A1(n7188), .A2(n7189), .A3(n2622), .Y(n2055) );
  AND4X1_LVT U3067 ( .A1(n7191), .A2(n7193), .A3(n7192), .A4(n2597), .Y(n2056)
         );
  OA21X1_LVT U3068 ( .A1(n3479), .A2(n2120), .A3(n7959), .Y(n7962) );
  AND4X1_LVT U3069 ( .A1(n2057), .A2(n2058), .A3(n2059), .A4(n2060), .Y(n2166)
         );
  AND2X1_LVT U3070 ( .A1(n8136), .A2(n8135), .Y(n2057) );
  AND4X1_LVT U3071 ( .A1(n8150), .A2(n8148), .A3(n8149), .A4(n2614), .Y(n2058)
         );
  AND3X1_LVT U3072 ( .A1(n8134), .A2(n8133), .A3(n8132), .Y(n2059) );
  AND3X1_LVT U3073 ( .A1(n8130), .A2(n8129), .A3(n8128), .Y(n2060) );
  AND3X1_LVT U3074 ( .A1(n2133), .A2(n2574), .A3(n2061), .Y(n2150) );
  AND3X1_LVT U3075 ( .A1(n2062), .A2(n2063), .A3(n2064), .Y(n3740) );
  AND3X1_LVT U3076 ( .A1(n8529), .A2(n8530), .A3(n8531), .Y(n2062) );
  AND2X1_LVT U3077 ( .A1(n8526), .A2(n8525), .Y(n2063) );
  AND3X1_LVT U3078 ( .A1(n8524), .A2(n8523), .A3(n8522), .Y(n2064) );
  NAND3X0_LVT U3079 ( .A1(n2065), .A2(n2066), .A3(n2067), .Y(N691) );
  AND3X1_LVT U3080 ( .A1(n2111), .A2(n2112), .A3(n2113), .Y(n2065) );
  AND3X1_LVT U3081 ( .A1(n7285), .A2(n7284), .A3(n7283), .Y(n2066) );
  AND3X1_LVT U3082 ( .A1(n7281), .A2(n7280), .A3(n7279), .Y(n2067) );
  AND2X1_LVT U3083 ( .A1(n2143), .A2(n6917), .Y(n2068) );
  NAND3X2_LVT U3084 ( .A1(n6940), .A2(n6972), .A3(n3772), .Y(n2069) );
  NAND2X4_LVT U3085 ( .A1(n5446), .A2(n5451), .Y(n3081) );
  AND2X1_LVT U3086 ( .A1(n2070), .A2(n2071), .Y(n2557) );
  AND3X1_LVT U3087 ( .A1(n8112), .A2(n8111), .A3(n8110), .Y(n2070) );
  AND3X1_LVT U3088 ( .A1(n8116), .A2(n8115), .A3(n8114), .Y(n2071) );
  NBUFFX2_LVT U3089 ( .A(ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n2072) );
  AND2X1_LVT U3090 ( .A1(n2073), .A2(n2074), .Y(n2109) );
  AND3X1_LVT U3091 ( .A1(n8168), .A2(n8167), .A3(n8166), .Y(n2073) );
  AND3X1_LVT U3092 ( .A1(n8164), .A2(n8163), .A3(n8162), .Y(n2074) );
  AND2X1_LVT U3093 ( .A1(n2075), .A2(n2076), .Y(n2095) );
  AND4X1_LVT U3094 ( .A1(n7174), .A2(n7172), .A3(n7173), .A4(n2586), .Y(n2075)
         );
  AND3X1_LVT U3095 ( .A1(n7187), .A2(n7186), .A3(n7185), .Y(n2076) );
  AND2X1_LVT U3096 ( .A1(n2077), .A2(n2078), .Y(n3742) );
  AND3X1_LVT U3097 ( .A1(n8452), .A2(n8450), .A3(n2579), .Y(n2077) );
  AND3X1_LVT U3098 ( .A1(n8449), .A2(n8448), .A3(n8447), .Y(n2078) );
  AND2X1_LVT U3099 ( .A1(n2079), .A2(n2080), .Y(n3739) );
  AND3X1_LVT U3100 ( .A1(n8516), .A2(n8514), .A3(n2580), .Y(n2079) );
  AND3X1_LVT U3101 ( .A1(n8513), .A2(n8512), .A3(n8511), .Y(n2080) );
  DELLN1X2_LVT U3102 ( .A(n8105), .Y(n2135) );
  NAND4X1_LVT U3103 ( .A1(n4954), .A2(n4955), .A3(n4953), .A4(n4952), .Y(n9282) );
  AND3X2_LVT U3104 ( .A1(n6940), .A2(n6972), .A3(n3772), .Y(n3689) );
  IBUFFX2_LVT U3105 ( .A(n3768), .Y(n2081) );
  AND2X1_LVT U3106 ( .A1(n2082), .A2(n2083), .Y(n3736) );
  AND3X1_LVT U3107 ( .A1(n8619), .A2(n8617), .A3(n2578), .Y(n2082) );
  AND3X1_LVT U3108 ( .A1(n8616), .A2(n8615), .A3(n8614), .Y(n2083) );
  AND2X1_LVT U3109 ( .A1(n2084), .A2(n2085), .Y(n2159) );
  AND3X1_LVT U3110 ( .A1(n8373), .A2(n8372), .A3(n8371), .Y(n2084) );
  AND3X1_LVT U3111 ( .A1(n8377), .A2(n8376), .A3(n8375), .Y(n2085) );
  OA21X2_LVT U3112 ( .A1(n2657), .A2(n2637), .A3(n2633), .Y(n2130) );
  AND3X1_LVT U3113 ( .A1(n7427), .A2(n7425), .A3(n2610), .Y(n2086) );
  AND3X1_LVT U3114 ( .A1(n7429), .A2(n7428), .A3(n3568), .Y(n2087) );
  AND3X1_LVT U3115 ( .A1(n7442), .A2(n7441), .A3(n7440), .Y(n2088) );
  IBUFFX2_LVT U3116 ( .A(n9036), .Y(n2089) );
  IBUFFX2_LVT U3117 ( .A(n9036), .Y(n2090) );
  AND2X4_LVT U3118 ( .A1(n6939), .A2(n6938), .Y(n9036) );
  NBUFFX2_LVT U3119 ( .A(n9016), .Y(n2091) );
  NBUFFX2_LVT U3120 ( .A(n9016), .Y(n2092) );
  NBUFFX2_LVT U3121 ( .A(n3613), .Y(n3610) );
  NBUFFX2_LVT U3122 ( .A(n9015), .Y(n2093) );
  NBUFFX2_LVT U3123 ( .A(n9015), .Y(n2094) );
  NAND3X0_LVT U3124 ( .A1(n2095), .A2(n2096), .A3(n2097), .Y(N687) );
  AND3X1_LVT U3125 ( .A1(n7171), .A2(n7170), .A3(n7169), .Y(n2097) );
  NBUFFX2_LVT U3126 ( .A(ibuf_io_inst_0_bits_inst_rs1[0]), .Y(n2098) );
  AND3X2_LVT U3127 ( .A1(n6940), .A2(n6926), .A3(n2983), .Y(n9016) );
  NAND3X0_LVT U3128 ( .A1(n2099), .A2(n2100), .A3(n2101), .Y(N726) );
  AND3X1_LVT U3129 ( .A1(n2124), .A2(n2125), .A3(n2126), .Y(n2099) );
  AND3X1_LVT U3130 ( .A1(n8408), .A2(n8407), .A3(n8406), .Y(n2100) );
  AND3X1_LVT U3131 ( .A1(n2117), .A2(n2118), .A3(n2119), .Y(n2101) );
  NAND3X0_LVT U3132 ( .A1(n2102), .A2(n2103), .A3(n2104), .Y(N742) );
  AND3X1_LVT U3133 ( .A1(n2114), .A2(n2115), .A3(n2116), .Y(n2102) );
  AND3X1_LVT U3134 ( .A1(n8974), .A2(n8973), .A3(n8972), .Y(n2103) );
  AND3X1_LVT U3135 ( .A1(n2162), .A2(n2163), .A3(n2164), .Y(n2104) );
  NAND3X0_LVT U3136 ( .A1(n2107), .A2(n2106), .A3(n2105), .Y(n2140) );
  AND2X1_LVT U3137 ( .A1(n3569), .A2(n2142), .Y(n2105) );
  AND4X1_LVT U3138 ( .A1(n7670), .A2(n7683), .A3(n7669), .A4(n2141), .Y(n2106)
         );
  AND3X1_LVT U3139 ( .A1(n7668), .A2(n2592), .A3(n7672), .Y(n2107) );
  AND3X2_LVT U3140 ( .A1(n3773), .A2(n6957), .A3(n6973), .Y(n3712) );
  AND3X2_LVT U3141 ( .A1(n6973), .A2(n6946), .A3(n2983), .Y(n9007) );
  AND3X2_LVT U3142 ( .A1(n6973), .A2(n6974), .A3(n3772), .Y(n2984) );
  AND2X4_LVT U3143 ( .A1(n2144), .A2(n6924), .Y(n6973) );
  NBUFFX2_LVT U3144 ( .A(n9026), .Y(n3760) );
  NBUFFX2_LVT U3145 ( .A(n9026), .Y(n3761) );
  AND3X2_LVT U3146 ( .A1(n6973), .A2(n6957), .A3(n2983), .Y(n9026) );
  NAND3X0_LVT U3147 ( .A1(n2108), .A2(n2109), .A3(n2110), .Y(N719) );
  AND3X1_LVT U3148 ( .A1(n8160), .A2(n8159), .A3(n8158), .Y(n2110) );
  AND3X1_LVT U3149 ( .A1(n7301), .A2(n7300), .A3(n7299), .Y(n2111) );
  AND4X1_LVT U3150 ( .A1(n2595), .A2(n7302), .A3(n7303), .A4(n7304), .Y(n2112)
         );
  AND3X1_LVT U3151 ( .A1(n7298), .A2(n7297), .A3(n7296), .Y(n2113) );
  AND3X1_LVT U3152 ( .A1(n8970), .A2(n8969), .A3(n8968), .Y(n2114) );
  AND3X1_LVT U3153 ( .A1(n8978), .A2(n8977), .A3(n8976), .Y(n2115) );
  AND4X1_LVT U3154 ( .A1(n8979), .A2(n2175), .A3(n2176), .A4(n2177), .Y(n2116)
         );
  AND3X1_LVT U3155 ( .A1(n8412), .A2(n8411), .A3(n8410), .Y(n2117) );
  AND3X1_LVT U3156 ( .A1(n8419), .A2(n8417), .A3(n2605), .Y(n2118) );
  AND3X1_LVT U3157 ( .A1(n8416), .A2(n8415), .A3(n8414), .Y(n2119) );
  NBUFFX2_LVT U3158 ( .A(n9006), .Y(n2120) );
  OR2X4_LVT U3159 ( .A1(n3140), .A2(n2120), .Y(n2668) );
  NBUFFX2_LVT U3160 ( .A(n9030), .Y(n3667) );
  NAND3X0_LVT U3161 ( .A1(n2121), .A2(n2122), .A3(n2123), .Y(N733) );
  AND3X1_LVT U3162 ( .A1(n8643), .A2(n8642), .A3(n8641), .Y(n2121) );
  AND4X1_LVT U3163 ( .A1(n3721), .A2(n3722), .A3(n8655), .A4(n8656), .Y(n2122)
         );
  NOR2X0_LVT U3164 ( .A1(n8670), .A2(n8669), .Y(n2123) );
  DELLN1X2_LVT U3165 ( .A(n5119), .Y(n2134) );
  AND3X1_LVT U3166 ( .A1(n8425), .A2(n8426), .A3(n8427), .Y(n2124) );
  AND3X1_LVT U3167 ( .A1(n8432), .A2(n8433), .A3(n8431), .Y(n2125) );
  AND2X1_LVT U3168 ( .A1(n8428), .A2(n8429), .Y(n2126) );
  AND3X1_LVT U3169 ( .A1(n4511), .A2(n4512), .A3(n4513), .Y(n3049) );
  AND3X2_LVT U3170 ( .A1(n2130), .A2(n5166), .A3(n9432), .Y(n2169) );
  OR2X2_LVT U3171 ( .A1(n3322), .A2(n2969), .Y(n2664) );
  OR2X2_LVT U3172 ( .A1(n3370), .A2(n3989), .Y(n2656) );
  NBUFFX2_LVT U3173 ( .A(n9026), .Y(n3758) );
  NBUFFX2_LVT U3174 ( .A(n9026), .Y(n3756) );
  NBUFFX2_LVT U3175 ( .A(n9026), .Y(n3759) );
  NBUFFX2_LVT U3176 ( .A(n9026), .Y(n3757) );
  NAND3X0_LVT U3177 ( .A1(n2127), .A2(n2128), .A3(n2129), .Y(N713) );
  AND3X1_LVT U3178 ( .A1(n7965), .A2(n7964), .A3(n7963), .Y(n2127) );
  AND3X1_LVT U3179 ( .A1(n2963), .A2(n2964), .A3(n2965), .Y(n2128) );
  AND2X4_LVT U3180 ( .A1(n5403), .A2(n5402), .Y(div_io_resp_ready) );
  DELLN2X2_LVT U3181 ( .A(n9381), .Y(n3046) );
  NAND3X2_LVT U3182 ( .A1(n9436), .A2(n2635), .A3(n5154), .Y(n5066) );
  NAND4X1_LVT U3183 ( .A1(n9075), .A2(n5164), .A3(io_fpu_inst[4]), .A4(n9104), 
        .Y(n2632) );
  AND2X4_LVT U3184 ( .A1(io_fpu_inst[5]), .A2(n9522), .Y(n3575) );
  AND3X4_LVT U3185 ( .A1(n3590), .A2(n3577), .A3(io_fpu_inst[6]), .Y(n5102) );
  OR3X2_LVT U3186 ( .A1(io_fpu_inst[23]), .A2(io_fpu_inst[24]), .A3(
        io_fpu_inst[22]), .Y(n5144) );
  IBUFFX2_LVT U3187 ( .A(ibuf_io_inst_0_bits_inst_rs2[4]), .Y(n5434) );
  AO21X2_LVT U3188 ( .A1(n9076), .A2(n3585), .A3(n3584), .Y(n2131) );
  NBUFFX2_LVT U3189 ( .A(n5423), .Y(n2132) );
  NBUFFX2_LVT U3190 ( .A(n9390), .Y(n2133) );
  NOR2X4_LVT U3191 ( .A1(n5306), .A2(n2132), .Y(n5356) );
  IBUFFX2_LVT U3192 ( .A(n9390), .Y(n9392) );
  AND3X2_LVT U3193 ( .A1(n3046), .A2(n2132), .A3(n5427), .Y(n5379) );
  AND2X4_LVT U3194 ( .A1(n5423), .A2(n5306), .Y(n5339) );
  DELLN1X2_LVT U3195 ( .A(n9022), .Y(n3642) );
  OR3X1_LVT U3196 ( .A1(n2461), .A2(n8078), .A3(n8080), .Y(N716) );
  AND3X1_LVT U3197 ( .A1(n7681), .A2(n7671), .A3(n7682), .Y(n2141) );
  AND2X4_LVT U3198 ( .A1(n2981), .A2(n3796), .Y(n6889) );
  AND2X4_LVT U3199 ( .A1(n2981), .A2(n3868), .Y(n6811) );
  AO21X2_LVT U3200 ( .A1(wb_ctrl_wxd), .A2(csr_io_retire), .A3(n9381), .Y(
        n9397) );
  NAND2X2_LVT U3201 ( .A1(n5415), .A2(n5403), .Y(n9381) );
  IBUFFX2_LVT U3202 ( .A(n5119), .Y(n2547) );
  NBUFFX2_LVT U3203 ( .A(n9519), .Y(io_fpu_inst[29]) );
  NBUFFX2_LVT U3204 ( .A(n2546), .Y(n2137) );
  IBUFFX4_LVT U3205 ( .A(n2546), .Y(n2537) );
  NAND2X0_LVT U3206 ( .A1(n9439), .A2(n2137), .Y(n2568) );
  NOR2X1_LVT U3207 ( .A1(n9517), .A2(n9519), .Y(n2546) );
  AO21X2_LVT U3208 ( .A1(io_fpu_inst[28]), .A2(n2138), .A3(n3039), .Y(n4843)
         );
  OR3X1_LVT U3209 ( .A1(n7684), .A2(n2140), .A3(n7685), .Y(N704) );
  OR2X2_LVT U3210 ( .A1(n9028), .A2(n3327), .Y(n2142) );
  AND3X1_LVT U3211 ( .A1(n2137), .A2(n9447), .A3(n2174), .Y(n4502) );
  NBUFFX2_LVT U3212 ( .A(n9029), .Y(n3637) );
  NAND3X2_LVT U3213 ( .A1(n5008), .A2(n5007), .A3(n5006), .Y(n3048) );
  OA21X2_LVT U3214 ( .A1(n9089), .A2(n9288), .A3(n2134), .Y(n5088) );
  NAND3X1_LVT U3215 ( .A1(n9107), .A2(n1891), .A3(io_fpu_inst[14]), .Y(n9088)
         );
  NAND3X1_LVT U3216 ( .A1(n4918), .A2(csr_io_decode_0_fp_csr), .A3(n2134), .Y(
        n4929) );
  NAND3X2_LVT U3217 ( .A1(n9288), .A2(csr_io_decode_0_write_illegal), .A3(
        n5119), .Y(n5120) );
  NAND3X2_LVT U3218 ( .A1(n5154), .A2(n3593), .A3(n9436), .Y(n5069) );
  OR2X4_LVT U3219 ( .A1(io_fpu_inst[14]), .A2(n3593), .Y(n4509) );
  DELLN1X2_LVT U3220 ( .A(n8932), .Y(n2859) );
  AND2X4_LVT U3221 ( .A1(n4749), .A2(n4752), .Y(n6974) );
  OR2X2_LVT U3222 ( .A1(n4752), .A2(n4969), .Y(n6955) );
  NAND2X0_LVT U3223 ( .A1(n2169), .A2(n2170), .Y(n2143) );
  NAND3X2_LVT U3224 ( .A1(n2533), .A2(n2532), .A3(n9388), .Y(n6935) );
  AND2X4_LVT U3225 ( .A1(n6972), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n9037) );
  AND2X4_LVT U3226 ( .A1(n6972), .A2(n6956), .Y(n8932) );
  AO21X2_LVT U3227 ( .A1(n7068), .A2(n7067), .A3(n3612), .Y(n7069) );
  AO21X2_LVT U3228 ( .A1(n7040), .A2(n7039), .A3(n3612), .Y(n7041) );
  AO21X2_LVT U3229 ( .A1(n7097), .A2(n7096), .A3(n3612), .Y(n7098) );
  AO21X2_LVT U3230 ( .A1(n6968), .A2(n6967), .A3(n3612), .Y(n6969) );
  AO21X2_LVT U3231 ( .A1(n7008), .A2(n7007), .A3(n3612), .Y(n7009) );
  NOR2X4_LVT U3232 ( .A1(n4040), .A2(n3612), .Y(n8939) );
  NOR2X4_LVT U3233 ( .A1(n3184), .A2(n9047), .Y(n8873) );
  NAND2X0_LVT U3234 ( .A1(n2145), .A2(n2146), .Y(n4511) );
  NOR3X4_LVT U3235 ( .A1(n2552), .A2(n4509), .A3(n4508), .Y(n2146) );
  NAND3X1_LVT U3236 ( .A1(n2677), .A2(n1863), .A3(io_fpu_inst[3]), .Y(n_GEN_9)
         );
  OA21X2_LVT U3237 ( .A1(n9438), .A2(n5129), .A3(n3076), .Y(n5068) );
  OR3X1_LVT U3238 ( .A1(n2147), .A2(n2148), .A3(n2149), .Y(n8849) );
  AND2X1_LVT U3239 ( .A1(n_T_427[186]), .A2(n3791), .Y(n2148) );
  DELLN1X2_LVT U3240 ( .A(n9056), .Y(n3600) );
  NBUFFX2_LVT U3241 ( .A(n9517), .Y(io_fpu_inst[31]) );
  AND3X4_LVT U3242 ( .A1(n9412), .A2(n9448), .A3(n9242), .Y(n9116) );
  NAND3X2_LVT U3243 ( .A1(n9412), .A2(n9099), .A3(n5167), .Y(n1431) );
  IBUFFX2_LVT U3244 ( .A(n3040), .Y(n2152) );
  AND2X1_LVT U3245 ( .A1(io_dmem_resp_valid), .A2(io_dmem_resp_bits_has_data), 
        .Y(n2153) );
  NOR2X4_LVT U3246 ( .A1(n9412), .A2(ibuf_io_inst_0_bits_rvc), .Y(n2529) );
  AND2X2_LVT U3247 ( .A1(n6939), .A2(n6936), .Y(n9412) );
  IBUFFX2_LVT U3248 ( .A(n3683), .Y(n2154) );
  IBUFFX2_LVT U3249 ( .A(n3683), .Y(n2155) );
  OA21X2_LVT U3250 ( .A1(n3407), .A2(n3691), .A3(n8561), .Y(n2603) );
  OA21X2_LVT U3251 ( .A1(n3405), .A2(n3708), .A3(n8323), .Y(n8326) );
  NAND3X0_LVT U3252 ( .A1(n2156), .A2(n2157), .A3(n2158), .Y(n8776) );
  AND3X1_LVT U3253 ( .A1(n8753), .A2(n8752), .A3(n2591), .Y(n2156) );
  AND4X1_LVT U3254 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n2638), .Y(n2157)
         );
  AND2X1_LVT U3255 ( .A1(n8755), .A2(n8754), .Y(n2158) );
  AO21X2_LVT U3256 ( .A1(n7588), .A2(n7587), .A3(n9047), .Y(n7589) );
  AO21X2_LVT U3257 ( .A1(n7467), .A2(n7466), .A3(n3631), .Y(n7468) );
  OR2X4_LVT U3258 ( .A1(n8457), .A2(n3612), .Y(n8458) );
  NAND3X0_LVT U3259 ( .A1(n2159), .A2(n2160), .A3(n2161), .Y(N725) );
  NOR3X0_LVT U3260 ( .A1(n8400), .A2(n8399), .A3(n8398), .Y(n2161) );
  AND3X1_LVT U3261 ( .A1(n8990), .A2(n8989), .A3(n8988), .Y(n2162) );
  AND2X1_LVT U3262 ( .A1(n8993), .A2(n8992), .Y(n2163) );
  AND3X1_LVT U3263 ( .A1(n8999), .A2(n8998), .A3(n8997), .Y(n2164) );
  AND3X1_LVT U3264 ( .A1(n8147), .A2(n8146), .A3(n8145), .Y(n2165) );
  AND3X1_LVT U3265 ( .A1(n8266), .A2(n8265), .A3(n8264), .Y(n2167) );
  NOR2X0_LVT U3266 ( .A1(n8276), .A2(n8275), .Y(n2168) );
  NAND2X0_LVT U3267 ( .A1(n2169), .A2(n2170), .Y(n6966) );
  AND3X2_LVT U3268 ( .A1(n5163), .A2(n9434), .A3(n2615), .Y(n5156) );
  NAND3X0_LVT U3269 ( .A1(n2171), .A2(n2172), .A3(n2173), .Y(N730) );
  AND3X1_LVT U3270 ( .A1(n8539), .A2(n8538), .A3(n8537), .Y(n2171) );
  AND3X1_LVT U3271 ( .A1(n8552), .A2(n8551), .A3(n8550), .Y(n2172) );
  NAND3X1_LVT U3272 ( .A1(n2553), .A2(n3079), .A3(n9434), .Y(n5114) );
  IBUFFX2_LVT U3273 ( .A(n9075), .Y(n2639) );
  AND2X1_LVT U3274 ( .A1(n2621), .A2(n6964), .Y(n2561) );
  OR3X1_LVT U3275 ( .A1(n9529), .A2(n9440), .A3(io_fpu_inst[27]), .Y(n4501) );
  OA21X1_LVT U3276 ( .A1(n3148), .A2(n3989), .A3(n8242), .Y(n8245) );
  NAND2X0_LVT U3277 ( .A1(n2527), .A2(n_T_427[447]), .Y(n2619) );
  IBUFFX2_LVT U3278 ( .A(n3715), .Y(n3994) );
  IBUFFX2_LVT U3279 ( .A(n5163), .Y(n9090) );
  OA21X1_LVT U3280 ( .A1(n3170), .A2(n2969), .A3(n9005), .Y(n9011) );
  NAND2X0_LVT U3281 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[17]), .Y(n7470)
         );
  OA21X1_LVT U3282 ( .A1(n3159), .A2(n2969), .A3(n8675), .Y(n8678) );
  NBUFFX2_LVT U3283 ( .A(n9523), .Y(io_fpu_inst[14]) );
  INVX1_LVT U3284 ( .A(n9516), .Y(io_ptw_status_debug) );
  OR2X1_LVT U3285 ( .A1(n9111), .A2(n9445), .Y(n9112) );
  IBUFFX2_LVT U3286 ( .A(io_fpu_inst[8]), .Y(n2174) );
  NAND2X0_LVT U3287 ( .A1(n_T_427[1149]), .A2(n3670), .Y(n2175) );
  OR2X1_LVT U3288 ( .A1(n4011), .A2(n3307), .Y(n2176) );
  NAND2X0_LVT U3289 ( .A1(n_T_427[1277]), .A2(n3641), .Y(n2177) );
  AO22X1_LVT U3290 ( .A1(io_fpu_dmem_resp_data[4]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[4]), .A4(n9065), .Y(n2178) );
  AO22X1_LVT U3291 ( .A1(n_T_628[4]), .A2(n2497), .A3(n_T_918[4]), .A4(n9066), 
        .Y(n2179) );
  OR2X1_LVT U3292 ( .A1(n2178), .A2(n2179), .Y(io_fpu_fromint_data[4]) );
  INVX0_LVT U3293 ( .A(n9492), .Y(n2180) );
  AO222X1_LVT U3294 ( .A1(n2180), .A2(n4060), .A3(n4063), .A4(csr_io_pc[30]), 
        .A5(csr_io_evec[30]), .A6(n4066), .Y(io_imem_req_bits_pc[30]) );
  AND4X1_LVT U3295 ( .A1(n3122), .A2(n3245), .A3(io_dmem_req_bits_cmd[1]), 
        .A4(io_dmem_req_bits_cmd[0]), .Y(n2181) );
  AO21X1_LVT U3296 ( .A1(io_dmem_req_bits_cmd[2]), .A2(n2181), .A3(n2515), .Y(
        n2516) );
  AND2X1_LVT U3297 ( .A1(n2572), .A2(n_T_1187[21]), .Y(n2182) );
  NAND2X0_LVT U3298 ( .A1(n5328), .A2(n5385), .Y(n2183) );
  AO22X1_LVT U3299 ( .A1(n5383), .A2(n5325), .A3(n2182), .A4(n2183), .Y(N767)
         );
  NAND4X0_LVT U3300 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .Y(n2184) );
  AO22X1_LVT U3301 ( .A1(n6813), .A2(n_T_427[832]), .A3(n_T_427[768]), .A4(
        n3906), .Y(n2185) );
  OA22X1_LVT U3302 ( .A1(n3081), .A2(n3138), .A3(n3530), .A4(n3880), .Y(n2186)
         );
  NAND2X0_LVT U3303 ( .A1(n4321), .A2(n3958), .Y(n2187) );
  NAND2X0_LVT U3304 ( .A1(n5479), .A2(n1992), .Y(n2188) );
  NAND4X0_LVT U3305 ( .A1(n2186), .A2(n9382), .A3(n2187), .A4(n2188), .Y(n2189) );
  OR3X1_LVT U3306 ( .A1(n2184), .A2(n2185), .A3(n2189), .Y(n2190) );
  NAND4X0_LVT U3307 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .Y(n2191) );
  INVX0_LVT U3308 ( .A(n5480), .Y(n2192) );
  OA21X1_LVT U3309 ( .A1(n2190), .A2(n2191), .A3(n2192), .Y(N679) );
  AOI22X1_LVT U3310 ( .A1(n_T_918[48]), .A2(n6855), .A3(io_fpu_toint_data[48]), 
        .A4(n6856), .Y(n2193) );
  NAND2X0_LVT U3311 ( .A1(n6857), .A2(n2193), .Y(N646) );
  INVX0_LVT U3312 ( .A(n9356), .Y(n2194) );
  INVX0_LVT U3313 ( .A(n123), .Y(n2195) );
  OA22X1_LVT U3314 ( .A1(n_T_698[18]), .A2(n9496), .A3(n_T_698[12]), .A4(n9491), .Y(n2196) );
  NAND2X0_LVT U3315 ( .A1(n9451), .A2(n9450), .Y(n2197) );
  NAND4X0_LVT U3316 ( .A1(n9453), .A2(n9471), .A3(n9472), .A4(n9452), .Y(n2198) );
  NOR4X0_LVT U3317 ( .A1(n_T_698[0]), .A2(n4599), .A3(n2197), .A4(n2198), .Y(
        n2199) );
  HADDX1_LVT U3318 ( .A0(n9334), .B0(n137), .SO(n2200) );
  OA21X1_LVT U3320 ( .A1(n_T_698[3]), .A2(n9503), .A3(n2202), .Y(n2203) );
  OA21X1_LVT U3321 ( .A1(n9495), .A2(n_T_698[4]), .A3(n2203), .Y(n2204) );
  OA21X1_LVT U3322 ( .A1(n9499), .A2(n_T_698[7]), .A3(n2204), .Y(n2205) );
  OA21X1_LVT U3323 ( .A1(n_T_698[6]), .A2(n9485), .A3(n2205), .Y(n2206) );
  OA21X1_LVT U3324 ( .A1(n_T_698[9]), .A2(n9507), .A3(n2206), .Y(n2207) );
  OA21X1_LVT U3325 ( .A1(n_T_698[8]), .A2(n9511), .A3(n2207), .Y(n2208) );
  OA22X1_LVT U3326 ( .A1(n_T_698[10]), .A2(n9509), .A3(n_T_698[14]), .A4(n9506), .Y(n2209) );
  OA221X1_LVT U3327 ( .A1(n9356), .A2(n123), .A3(n2194), .A4(n2195), .A5(n2211), .Y(n4600) );
  AO22X1_LVT U3328 ( .A1(io_fpu_dmem_resp_data[5]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[5]), .A4(n9065), .Y(n2212) );
  AO22X1_LVT U3329 ( .A1(n_T_628[5]), .A2(n2493), .A3(n_T_918[5]), .A4(n9066), 
        .Y(n2213) );
  OR2X1_LVT U3330 ( .A1(n2212), .A2(n2213), .Y(io_fpu_fromint_data[5]) );
  AO222X1_LVT U3331 ( .A1(n4065), .A2(csr_io_evec[39]), .A3(n9377), .A4(n4059), 
        .A5(n4062), .A6(csr_io_pc[39]), .Y(io_imem_req_bits_pc[39]) );
  NAND2X0_LVT U3332 ( .A1(n5357), .A2(n5356), .Y(n2214) );
  AND2X1_LVT U3333 ( .A1(n_T_1187[2]), .A2(n2214), .Y(n2215) );
  AO22X1_LVT U3334 ( .A1(n2572), .A2(n2215), .A3(n5355), .A4(n5374), .Y(N748)
         );
  AND4X1_LVT U3335 ( .A1(n2973), .A2(n7201), .A3(n7199), .A4(n7200), .Y(n2216)
         );
  AND4X1_LVT U3336 ( .A1(n7216), .A2(n7217), .A3(n7195), .A4(n7196), .Y(n2217)
         );
  AND3X1_LVT U3337 ( .A1(n7218), .A2(n7197), .A3(n2217), .Y(n2218) );
  NAND3X0_LVT U3338 ( .A1(n2974), .A2(n2216), .A3(n2218), .Y(N688) );
  AO222X1_LVT U3339 ( .A1(n9293), .A2(n2515), .A3(n_T_702[24]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[56]), .Y(N517) );
  AO22X1_LVT U3340 ( .A1(n2872), .A2(n_T_427[68]), .A3(n_T_427[1027]), .A4(
        n3900), .Y(n2219) );
  AO22X1_LVT U3341 ( .A1(n2865), .A2(n_T_427[388]), .A3(n_T_427[771]), .A4(
        n3907), .Y(n2220) );
  AO22X1_LVT U3342 ( .A1(n3909), .A2(n_T_427[132]), .A3(n_T_427[452]), .A4(
        n3912), .Y(n2221) );
  AO22X1_LVT U3343 ( .A1(n2879), .A2(n_T_427[4]), .A3(n_T_427[516]), .A4(n2851), .Y(n2222) );
  NOR4X0_LVT U3344 ( .A1(n2219), .A2(n2220), .A3(n2221), .A4(n2222), .Y(n2223)
         );
  AO22X1_LVT U3345 ( .A1(n3917), .A2(n_T_427[1347]), .A3(n_T_427[1475]), .A4(
        n3923), .Y(n2224) );
  AO22X1_LVT U3346 ( .A1(n3927), .A2(n_T_427[1283]), .A3(n_T_427[1411]), .A4(
        n3933), .Y(n2225) );
  AO22X1_LVT U3347 ( .A1(n3937), .A2(n_T_427[1219]), .A3(n_T_427[1155]), .A4(
        n3943), .Y(n2226) );
  AO22X1_LVT U3348 ( .A1(n3947), .A2(n_T_427[963]), .A3(n_T_427[1091]), .A4(
        n3953), .Y(n2227) );
  NOR4X0_LVT U3349 ( .A1(n2224), .A2(n2225), .A3(n2226), .A4(n2227), .Y(n2228)
         );
  NAND2X0_LVT U3350 ( .A1(n4330), .A2(n3958), .Y(n2230) );
  NAND4X0_LVT U3351 ( .A1(n2223), .A2(n2228), .A3(n2229), .A4(n2230), .Y(
        id_rs_1[4]) );
  AOI22X1_LVT U3352 ( .A1(n_T_918[49]), .A2(n6855), .A3(io_fpu_toint_data[49]), 
        .A4(n6856), .Y(n2231) );
  NAND2X0_LVT U3353 ( .A1(n6857), .A2(n2231), .Y(N647) );
  INVX0_LVT U3354 ( .A(n_T_728[0]), .Y(n2232) );
  AOI21X1_LVT U3355 ( .A1(n_T_726[1]), .A2(n2232), .A3(n_T_728[1]), .Y(n2233)
         );
  AO221X1_LVT U3356 ( .A1(n9242), .A2(bpu_io_xcpt_if), .A3(n9242), .A4(n2233), 
        .A5(csr_io_interrupt), .Y(n74) );
  OAI22X1_LVT U3357 ( .A1(n589), .A2(n9163), .A3(n159), .A4(n9164), .Y(n2234)
         );
  NAND3X0_LVT U3358 ( .A1(n9157), .A2(n9155), .A3(n9156), .Y(n2235) );
  OA221X1_LVT U3359 ( .A1(n2235), .A2(io_fpu_dmem_resp_data[3]), .A3(n2235), 
        .A4(n9165), .A5(n9227), .Y(n2236) );
  AO222X1_LVT U3361 ( .A1(n4061), .A2(n9373), .A3(n4066), .A4(csr_io_evec[34]), 
        .A5(csr_io_pc[34]), .A6(n4062), .Y(io_imem_req_bits_pc[34]) );
  INVX0_LVT U3362 ( .A(n9230), .Y(n2238) );
  NAND2X0_LVT U3363 ( .A1(n3583), .A2(n5164), .Y(n2239) );
  OA221X1_LVT U3365 ( .A1(n2669), .A2(n5108), .A3(n2669), .A4(n2629), .A5(
        n2241), .Y(n5166) );
  AND2X1_LVT U3366 ( .A1(n_T_1187[24]), .A2(n2572), .Y(n2242) );
  NAND2X0_LVT U3367 ( .A1(n5379), .A2(n5307), .Y(n2243) );
  AO22X1_LVT U3368 ( .A1(n5366), .A2(n5305), .A3(n2242), .A4(n2243), .Y(N770)
         );
  AO222X1_LVT U3369 ( .A1(n_T_702[23]), .A2(n9301), .A3(n_T_702[7]), .A4(n2515), .A5(n4058), .A6(n_T_702[55]), .Y(N516) );
  AO22X1_LVT U3370 ( .A1(n3932), .A2(n_T_427[1445]), .A3(n_T_427[1381]), .A4(
        n3921), .Y(n2244) );
  AO22X1_LVT U3371 ( .A1(n3942), .A2(n_T_427[1189]), .A3(n_T_427[1317]), .A4(
        n3931), .Y(n2245) );
  AO22X1_LVT U3372 ( .A1(n3952), .A2(n_T_427[1125]), .A3(n_T_427[1253]), .A4(
        n3938), .Y(n2246) );
  AO22X1_LVT U3373 ( .A1(n3898), .A2(n_T_427[1061]), .A3(n_T_427[997]), .A4(
        n3948), .Y(n2247) );
  NOR4X0_LVT U3374 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .Y(n2248)
         );
  NOR4X0_LVT U3375 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .Y(n2250)
         );
  NAND3X0_LVT U3376 ( .A1(n2248), .A2(n2249), .A3(n2250), .Y(id_rs_1[38]) );
  AOI22X1_LVT U3377 ( .A1(n_T_918[50]), .A2(n6855), .A3(io_fpu_toint_data[50]), 
        .A4(n6856), .Y(n2251) );
  NAND2X0_LVT U3378 ( .A1(n6857), .A2(n2251), .Y(N648) );
  INVX0_LVT U3379 ( .A(n9448), .Y(n2252) );
  OR3X1_LVT U3380 ( .A1(bpu_io_xcpt_if), .A2(n_T_726[0]), .A3(n_T_728[0]), .Y(
        n2253) );
  OA221X1_LVT U3381 ( .A1(n9448), .A2(csr_io_interrupt_cause[0]), .A3(n2252), 
        .A4(n2253), .A5(n74), .Y(N303) );
  AO22X1_LVT U3382 ( .A1(io_fpu_dmem_resp_data[6]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[6]), .A4(n9065), .Y(n2254) );
  AO22X1_LVT U3383 ( .A1(n_T_628[6]), .A2(n2497), .A3(n_T_918[6]), .A4(n9066), 
        .Y(n2255) );
  OR2X1_LVT U3384 ( .A1(n2254), .A2(n2255), .Y(io_fpu_fromint_data[6]) );
  AO222X1_LVT U3385 ( .A1(n9302), .A2(n2515), .A3(n_T_702[63]), .A4(n4058), 
        .A5(n9301), .A6(n_T_702[31]), .Y(N524) );
  AO22X1_LVT U3386 ( .A1(n3919), .A2(n_T_427[1375]), .A3(n_T_427[1503]), .A4(
        n3924), .Y(n2256) );
  AO22X1_LVT U3387 ( .A1(n3928), .A2(n_T_427[1311]), .A3(n_T_427[1439]), .A4(
        n3934), .Y(n2257) );
  AO22X1_LVT U3388 ( .A1(n3939), .A2(n_T_427[1247]), .A3(n_T_427[1183]), .A4(
        n3944), .Y(n2258) );
  AO22X1_LVT U3389 ( .A1(n3949), .A2(n_T_427[991]), .A3(n_T_427[1119]), .A4(
        n3954), .Y(n2259) );
  NOR4X0_LVT U3390 ( .A1(n2256), .A2(n2257), .A3(n2258), .A4(n2259), .Y(n2260)
         );
  AOI22X1_LVT U3391 ( .A1(n6884), .A2(n_T_427[736]), .A3(n_T_427[96]), .A4(
        n2872), .Y(n2261) );
  AND4X1_LVT U3392 ( .A1(n2261), .A2(n2689), .A3(n2688), .A4(n2687), .Y(n2262)
         );
  AOI22X1_LVT U3393 ( .A1(n3888), .A2(n_T_427[1631]), .A3(n_T_427[1567]), .A4(
        n3894), .Y(n2263) );
  OA22X1_LVT U3394 ( .A1(n3081), .A2(n3143), .A3(n3082), .A4(n3496), .Y(n2264)
         );
  OA22X1_LVT U3395 ( .A1(n3878), .A2(n6110), .A3(n3276), .A4(n3881), .Y(n2265)
         );
  OA22X2_LVT U3396 ( .A1(n3803), .A2(n3144), .A3(n3495), .A4(n3800), .Y(n2266)
         );
  AND4X1_LVT U3397 ( .A1(n2263), .A2(n2264), .A3(n2265), .A4(n2266), .Y(n2267)
         );
  NAND2X0_LVT U3398 ( .A1(n4406), .A2(n3957), .Y(n2268) );
  NAND4X0_LVT U3399 ( .A1(n2260), .A2(n2262), .A3(n2267), .A4(n2268), .Y(
        id_rs_1[32]) );
  AOI22X1_LVT U3400 ( .A1(n_T_918[51]), .A2(n6855), .A3(io_fpu_toint_data[51]), 
        .A4(n6856), .Y(n2269) );
  NAND2X0_LVT U3401 ( .A1(n6857), .A2(n2269), .Y(N649) );
  AOI22X1_LVT U3402 ( .A1(n9500), .A2(ibuf_io_pc[13]), .A3(n9509), .A4(
        ibuf_io_pc[10]), .Y(n2270) );
  OA221X1_LVT U3403 ( .A1(n9500), .A2(ibuf_io_pc[13]), .A3(n9509), .A4(
        ibuf_io_pc[10]), .A5(n2270), .Y(n2271) );
  INVX0_LVT U3404 ( .A(ibuf_io_pc[15]), .Y(n2272) );
  AOI22X1_LVT U3405 ( .A1(n2272), .A2(n9355), .A3(n9490), .A4(ibuf_io_pc[11]), 
        .Y(n2273) );
  OA221X1_LVT U3406 ( .A1(n2272), .A2(n9355), .A3(n9490), .A4(ibuf_io_pc[11]), 
        .A5(n2273), .Y(n2274) );
  AOI22X1_LVT U3407 ( .A1(n9510), .A2(ibuf_io_pc[19]), .A3(n9504), .A4(
        ibuf_io_pc[29]), .Y(n2275) );
  OA221X1_LVT U3408 ( .A1(n9510), .A2(ibuf_io_pc[19]), .A3(n9504), .A4(
        ibuf_io_pc[29]), .A5(n2275), .Y(n2276) );
  INVX0_LVT U3409 ( .A(ibuf_io_pc[21]), .Y(n2277) );
  INVX0_LVT U3410 ( .A(n9361), .Y(n2278) );
  AO22X1_LVT U3411 ( .A1(ibuf_io_pc[21]), .A2(n9361), .A3(n2277), .A4(n2278), 
        .Y(n2279) );
  NAND4X0_LVT U3412 ( .A1(n2271), .A2(n2274), .A3(n2276), .A4(n2279), .Y(n4575) );
  INVX0_LVT U3413 ( .A(n5426), .Y(n2280) );
  AND2X1_LVT U3414 ( .A1(n2280), .A2(n5428), .Y(n5384) );
  AO22X1_LVT U3415 ( .A1(io_fpu_dmem_resp_data[8]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[8]), .A4(n9065), .Y(n2281) );
  AO22X1_LVT U3416 ( .A1(n_T_628[8]), .A2(n2493), .A3(n_T_918[8]), .A4(n9066), 
        .Y(n2282) );
  OR2X1_LVT U3417 ( .A1(n2281), .A2(n2282), .Y(io_fpu_fromint_data[8]) );
  AO22X1_LVT U3418 ( .A1(io_fpu_dmem_resp_data[16]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[16]), .A4(n9065), .Y(n2283) );
  AO22X1_LVT U3419 ( .A1(n_T_628[16]), .A2(n2497), .A3(n_T_918[16]), .A4(n9066), .Y(n2284) );
  OR2X1_LVT U3420 ( .A1(n2283), .A2(n2284), .Y(io_fpu_fromint_data[16]) );
  AO222X1_LVT U3421 ( .A1(n_T_702[22]), .A2(n9301), .A3(n_T_702[6]), .A4(n2515), .A5(n4058), .A6(n_T_702[54]), .Y(N515) );
  AO22X1_LVT U3422 ( .A1(n3932), .A2(n_T_427[1435]), .A3(n_T_427[1371]), .A4(
        n3921), .Y(n2285) );
  AO22X1_LVT U3423 ( .A1(n3942), .A2(n_T_427[1179]), .A3(n_T_427[1307]), .A4(
        n3931), .Y(n2286) );
  AO22X1_LVT U3424 ( .A1(n3952), .A2(n_T_427[1115]), .A3(n_T_427[1243]), .A4(
        n3941), .Y(n2287) );
  AO22X1_LVT U3425 ( .A1(n3898), .A2(n_T_427[1051]), .A3(n_T_427[987]), .A4(
        n3951), .Y(n2288) );
  NOR4X0_LVT U3426 ( .A1(n2285), .A2(n2286), .A3(n2287), .A4(n2288), .Y(n2289)
         );
  NOR4X0_LVT U3427 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .Y(n2291)
         );
  NAND3X0_LVT U3428 ( .A1(n2289), .A2(n2290), .A3(n2291), .Y(id_rs_1[28]) );
  AOI22X1_LVT U3429 ( .A1(n_T_918[52]), .A2(n6855), .A3(io_fpu_toint_data[52]), 
        .A4(n6856), .Y(n2292) );
  NAND2X0_LVT U3430 ( .A1(n6857), .A2(n2292), .Y(N650) );
  AO22X1_LVT U3431 ( .A1(n9510), .A2(n_T_698[19]), .A3(n9501), .A4(n_T_698[22]), .Y(n2293) );
  AO22X1_LVT U3432 ( .A1(n9488), .A2(n_T_698[23]), .A3(n9497), .A4(n_T_698[25]), .Y(n2294) );
  AO22X1_LVT U3433 ( .A1(n9499), .A2(n_T_698[7]), .A3(n9502), .A4(n_T_698[31]), 
        .Y(n2295) );
  AO22X1_LVT U3434 ( .A1(n9512), .A2(n_T_698[1]), .A3(n9495), .A4(n_T_698[4]), 
        .Y(n2296) );
  OR4X1_LVT U3435 ( .A1(n2293), .A2(n2294), .A3(n2295), .A4(n2296), .Y(n4599)
         );
  INVX0_LVT U3436 ( .A(n5423), .Y(n2297) );
  AND2X1_LVT U3437 ( .A1(n2297), .A2(n5306), .Y(n5335) );
  AO22X1_LVT U3438 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[11]), .A3(
        n_T_918[11]), .A4(n6899), .Y(n2298) );
  AO22X1_LVT U3439 ( .A1(n_T_635[11]), .A2(n6901), .A3(
        io_imem_sfence_bits_addr[11]), .A4(n6900), .Y(n2299) );
  OR2X1_LVT U3440 ( .A1(n2298), .A2(n2299), .Y(n_T_702[11]) );
  AO22X1_LVT U3441 ( .A1(io_fpu_dmem_resp_data[9]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[9]), .A4(n9065), .Y(n2300) );
  AO22X1_LVT U3442 ( .A1(n_T_628[9]), .A2(n2497), .A3(n_T_918[9]), .A4(n9066), 
        .Y(n2301) );
  OR2X1_LVT U3443 ( .A1(n2300), .A2(n2301), .Y(io_fpu_fromint_data[9]) );
  AO22X1_LVT U3444 ( .A1(io_fpu_dmem_resp_data[17]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[17]), .A4(n9065), .Y(n2302) );
  AO22X1_LVT U3445 ( .A1(n_T_628[17]), .A2(n2497), .A3(n_T_918[17]), .A4(n9066), .Y(n2303) );
  OR2X1_LVT U3446 ( .A1(n2302), .A2(n2303), .Y(io_fpu_fromint_data[17]) );
  NAND2X0_LVT U3447 ( .A1(n_T_427[1626]), .A2(n3648), .Y(n2304) );
  AND3X1_LVT U3448 ( .A1(n2304), .A2(n7761), .A3(n7762), .Y(n2305) );
  AND4X1_LVT U3449 ( .A1(n7759), .A2(n2305), .A3(n7758), .A4(n7757), .Y(n2306)
         );
  NAND4X0_LVT U3450 ( .A1(n3061), .A2(n2306), .A3(n3062), .A4(n3063), .Y(N707)
         );
  AO222X1_LVT U3451 ( .A1(n9300), .A2(n2515), .A3(n_T_702[30]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[62]), .Y(N523) );
  AO22X1_LVT U3452 ( .A1(n2862), .A2(n_T_427[144]), .A3(n_T_427[464]), .A4(
        n2824), .Y(n2307) );
  AO22X1_LVT U3453 ( .A1(n3810), .A2(n_T_427[272]), .A3(n3820), .A4(
        n_T_427[656]), .Y(n2308) );
  AO22X1_LVT U3454 ( .A1(n3835), .A2(n_T_427[400]), .A3(n3898), .A4(
        n_T_427[1039]), .Y(n2309) );
  AO22X1_LVT U3455 ( .A1(n3903), .A2(n_T_427[720]), .A3(n_T_427[783]), .A4(
        n2860), .Y(n2310) );
  NOR4X0_LVT U3456 ( .A1(n2307), .A2(n2308), .A3(n2309), .A4(n2310), .Y(n2311)
         );
  AO22X1_LVT U3457 ( .A1(n3918), .A2(n_T_427[1359]), .A3(n_T_427[1487]), .A4(
        n3923), .Y(n2312) );
  AO22X1_LVT U3458 ( .A1(n3928), .A2(n_T_427[1295]), .A3(n_T_427[1423]), .A4(
        n3933), .Y(n2313) );
  AO22X1_LVT U3459 ( .A1(n3938), .A2(n_T_427[1231]), .A3(n_T_427[1167]), .A4(
        n3943), .Y(n2314) );
  AO22X1_LVT U3460 ( .A1(n3948), .A2(n_T_427[975]), .A3(n_T_427[1103]), .A4(
        n3953), .Y(n2315) );
  NOR4X0_LVT U3461 ( .A1(n2312), .A2(n2313), .A3(n2314), .A4(n2315), .Y(n2316)
         );
  AOI22X1_LVT U3462 ( .A1(n3886), .A2(n_T_427[1615]), .A3(n_T_427[1551]), .A4(
        n3891), .Y(n2317) );
  AOI22X1_LVT U3463 ( .A1(n3826), .A2(n_T_427[1679]), .A3(n_T_427[1806]), .A4(
        n3830), .Y(n2318) );
  AND4X1_LVT U3464 ( .A1(n2317), .A2(n2755), .A3(n2756), .A4(n2318), .Y(n2319)
         );
  NAND2X0_LVT U3465 ( .A1(n4364), .A2(n3957), .Y(n2320) );
  NAND4X0_LVT U3466 ( .A1(n2311), .A2(n2316), .A3(n2319), .A4(n2320), .Y(
        id_rs_1[16]) );
  AOI22X1_LVT U3467 ( .A1(n_T_918[53]), .A2(n6855), .A3(io_fpu_toint_data[53]), 
        .A4(n6856), .Y(n2321) );
  NAND2X0_LVT U3468 ( .A1(n6857), .A2(n2321), .Y(N651) );
  AO22X1_LVT U3469 ( .A1(n_T_427[252]), .A2(n3986), .A3(n_T_427[636]), .A4(
        n4034), .Y(n2322) );
  AO22X1_LVT U3470 ( .A1(n4052), .A2(n_T_427[60]), .A3(n_T_427[188]), .A4(
        n2859), .Y(n2323) );
  AO22X1_LVT U3471 ( .A1(n_T_427[700]), .A2(n4021), .A3(n_T_427[955]), .A4(
        n4023), .Y(n2324) );
  OR3X1_LVT U3472 ( .A1(n2322), .A2(n2323), .A3(n2324), .Y(n8902) );
  AO22X1_LVT U3473 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[27]), .A3(
        n_T_918[27]), .A4(n6899), .Y(n2325) );
  AO22X1_LVT U3474 ( .A1(n_T_635[27]), .A2(n6901), .A3(
        io_imem_sfence_bits_addr[27]), .A4(n6900), .Y(n2326) );
  OR2X1_LVT U3475 ( .A1(n2325), .A2(n2326), .Y(n_T_702[27]) );
  AO22X1_LVT U3476 ( .A1(n4054), .A2(n_T_698[1]), .A3(n9103), .A4(
        io_fpu_fromint_data[1]), .Y(alu_io_in1[1]) );
  AO22X1_LVT U3477 ( .A1(io_fpu_dmem_resp_data[12]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[12]), .A4(n9065), .Y(n2327) );
  AO22X1_LVT U3478 ( .A1(n_T_628[12]), .A2(n2497), .A3(n_T_918[12]), .A4(n9066), .Y(n2328) );
  OR2X1_LVT U3479 ( .A1(n2327), .A2(n2328), .Y(io_fpu_fromint_data[12]) );
  NOR4X0_LVT U3480 ( .A1(n8197), .A2(n8196), .A3(n8206), .A4(n8205), .Y(n2329)
         );
  NAND2X0_LVT U3481 ( .A1(n3746), .A2(n2329), .Y(N720) );
  AND2X1_LVT U3482 ( .A1(n_T_1187[26]), .A2(n2572), .Y(n2330) );
  NAND2X0_LVT U3483 ( .A1(n5356), .A2(n5307), .Y(n2331) );
  AO22X1_LVT U3484 ( .A1(n5374), .A2(n5305), .A3(n2330), .A4(n2331), .Y(N772)
         );
  AO222X1_LVT U3485 ( .A1(n9299), .A2(n2515), .A3(n_T_702[29]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[61]), .Y(N522) );
  AO22X1_LVT U3486 ( .A1(n3923), .A2(n_T_427[1485]), .A3(n_T_427[1357]), .A4(
        n3918), .Y(n2332) );
  AO22X1_LVT U3487 ( .A1(n3933), .A2(n_T_427[1421]), .A3(n_T_427[1293]), .A4(
        n3928), .Y(n2333) );
  AO22X1_LVT U3488 ( .A1(n3943), .A2(n_T_427[1165]), .A3(n_T_427[1229]), .A4(
        n3938), .Y(n2334) );
  AO22X1_LVT U3489 ( .A1(n3953), .A2(n_T_427[1101]), .A3(n_T_427[973]), .A4(
        n3948), .Y(n2335) );
  NOR4X0_LVT U3490 ( .A1(n2332), .A2(n2333), .A3(n2334), .A4(n2335), .Y(n2336)
         );
  NOR4X0_LVT U3491 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .Y(n2338)
         );
  NAND4X0_LVT U3492 ( .A1(n2336), .A2(n2337), .A3(n2819), .A4(n2338), .Y(
        id_rs_1[14]) );
  AOI22X1_LVT U3493 ( .A1(n_T_918[54]), .A2(n6855), .A3(io_fpu_toint_data[54]), 
        .A4(n6856), .Y(n2339) );
  NAND2X0_LVT U3494 ( .A1(n6857), .A2(n2339), .Y(N652) );
  AO22X1_LVT U3495 ( .A1(n_T_427[48]), .A2(n4051), .A3(n_T_427[176]), .A4(
        n2859), .Y(n2340) );
  AO22X1_LVT U3496 ( .A1(n4027), .A2(n_T_427[879]), .A3(n_T_427[624]), .A4(
        n4035), .Y(n2341) );
  AO22X1_LVT U3497 ( .A1(n_T_427[240]), .A2(n3983), .A3(n_T_427[688]), .A4(
        n4022), .Y(n2342) );
  OR3X1_LVT U3498 ( .A1(n2340), .A2(n2341), .A3(n2342), .Y(n8470) );
  AO22X1_LVT U3499 ( .A1(io_fpu_dmem_resp_data[3]), .A2(n9064), .A3(n9065), 
        .A4(io_imem_sfence_bits_addr[3]), .Y(n2343) );
  AO22X1_LVT U3500 ( .A1(n9066), .A2(n_T_918[3]), .A3(n2497), .A4(n_T_628[3]), 
        .Y(n2344) );
  OR2X1_LVT U3501 ( .A1(n2343), .A2(n2344), .Y(io_fpu_fromint_data[3]) );
  INVX0_LVT U3502 ( .A(n9508), .Y(n2345) );
  AO222X1_LVT U3503 ( .A1(n2345), .A2(n4061), .A3(csr_io_evec[36]), .A4(n4067), 
        .A5(csr_io_pc[36]), .A6(n4062), .Y(io_imem_req_bits_pc[36]) );
  INVX0_LVT U3504 ( .A(N290), .Y(n2346) );
  NAND4X0_LVT U3505 ( .A1(n5090), .A2(io_dmem_req_bits_cmd[2]), .A3(n559), 
        .A4(io_dmem_req_bits_cmd[4]), .Y(n2347) );
  NAND3X0_LVT U3506 ( .A1(n9426), .A2(n5091), .A3(mem_reg_sfence), .Y(n2348)
         );
  OA21X1_LVT U3507 ( .A1(n2346), .A2(n2347), .A3(n2348), .Y(n2525) );
  AND2X1_LVT U3508 ( .A1(n_T_1187[25]), .A2(n2572), .Y(n2349) );
  NAND2X0_LVT U3509 ( .A1(n5339), .A2(n5307), .Y(n2350) );
  AO22X1_LVT U3510 ( .A1(n5383), .A2(n5305), .A3(n2349), .A4(n2350), .Y(N771)
         );
  AO22X1_LVT U3511 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[7]), .A3(n_T_918[7]), .A4(n6899), .Y(n2351) );
  AO22X1_LVT U3512 ( .A1(n_T_635[7]), .A2(n6901), .A3(
        io_imem_sfence_bits_addr[7]), .A4(n6900), .Y(n2352) );
  OR2X1_LVT U3513 ( .A1(n2351), .A2(n2352), .Y(n_T_702[7]) );
  AO222X1_LVT U3514 ( .A1(n9298), .A2(n2515), .A3(n_T_702[28]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[60]), .Y(N521) );
  AO222X1_LVT U3515 ( .A1(n6249), .A2(mem_br_target[11]), .A3(n_T_918[11]), 
        .A4(n6855), .A5(io_fpu_toint_data[11]), .A6(n6856), .Y(N609) );
  AOI22X1_LVT U3516 ( .A1(n_T_918[55]), .A2(n6855), .A3(io_fpu_toint_data[55]), 
        .A4(n6856), .Y(n2353) );
  NAND2X0_LVT U3517 ( .A1(n6857), .A2(n2353), .Y(N653) );
  AO22X1_LVT U3518 ( .A1(n_T_427[748]), .A2(n4048), .A3(n_T_427[812]), .A4(
        n3982), .Y(n2354) );
  NOR4X0_LVT U3519 ( .A1(n8387), .A2(n8386), .A3(n8385), .A4(n2354), .Y(n2355)
         );
  OR2X1_LVT U3520 ( .A1(n3656), .A2(n2355), .Y(n8388) );
  AO222X1_LVT U3521 ( .A1(n3852), .A2(io_dmem_resp_bits_data[22]), .A3(
        div_io_resp_bits_data[22]), .A4(n3855), .A5(n3849), .A6(
        io_imem_sfence_bits_addr[22]), .Y(n2356) );
  AOI21X1_LVT U3522 ( .A1(csr_io_rw_rdata[22]), .A2(n3844), .A3(n2356), .Y(
        n3094) );
  AOI22X1_LVT U3523 ( .A1(n3910), .A2(n_T_427[448]), .A3(n_T_427[320]), .A4(
        n1918), .Y(n2357) );
  AOI22X1_LVT U3524 ( .A1(n6830), .A2(n_T_427[384]), .A3(n_T_427[767]), .A4(
        n3906), .Y(n2358) );
  AND4X1_LVT U3525 ( .A1(n2357), .A2(n2358), .A3(n2881), .A4(n2880), .Y(n5464)
         );
  AO22X1_LVT U3526 ( .A1(io_fpu_dmem_resp_data[2]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[2]), .A4(n9065), .Y(n2359) );
  AO22X1_LVT U3527 ( .A1(n_T_628[2]), .A2(n2493), .A3(n_T_918[2]), .A4(n9066), 
        .Y(n2360) );
  OR2X1_LVT U3528 ( .A1(n2359), .A2(n2360), .Y(io_fpu_fromint_data[2]) );
  AO22X1_LVT U3529 ( .A1(io_fpu_dmem_resp_data[19]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[19]), .A4(n9065), .Y(n2361) );
  AO22X1_LVT U3530 ( .A1(n_T_628[19]), .A2(n2497), .A3(n_T_918[19]), .A4(n9066), .Y(n2362) );
  OR2X1_LVT U3531 ( .A1(n2361), .A2(n2362), .Y(io_fpu_fromint_data[19]) );
  AO22X1_LVT U3532 ( .A1(io_fpu_dmem_resp_data[29]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[29]), .A4(n9065), .Y(n2363) );
  AO22X1_LVT U3533 ( .A1(n_T_628[29]), .A2(n2497), .A3(n_T_918[29]), .A4(n9066), .Y(n2364) );
  OR2X1_LVT U3534 ( .A1(n2363), .A2(n2364), .Y(io_fpu_fromint_data[29]) );
  NAND2X0_LVT U3535 ( .A1(n3734), .A2(n2365), .Y(N737) );
  AO222X1_LVT U3536 ( .A1(n9297), .A2(n2515), .A3(n_T_702[27]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[59]), .Y(N520) );
  AO222X1_LVT U3537 ( .A1(n6249), .A2(mem_br_target[13]), .A3(n_T_918[13]), 
        .A4(n6855), .A5(io_fpu_toint_data[13]), .A6(n6856), .Y(N611) );
  AOI22X1_LVT U3538 ( .A1(n_T_918[56]), .A2(n6855), .A3(io_fpu_toint_data[56]), 
        .A4(n6856), .Y(n2366) );
  NAND2X0_LVT U3539 ( .A1(n6857), .A2(n2366), .Y(N654) );
  NAND3X0_LVT U3540 ( .A1(n5092), .A2(n5093), .A3(n5094), .Y(n2367) );
  AND2X1_LVT U3541 ( .A1(mem_ctrl_mem), .A2(n2367), .Y(n9424) );
  NOR4X0_LVT U3542 ( .A1(n7680), .A2(n7679), .A3(n7678), .A4(n7677), .Y(n2368)
         );
  NOR4X0_LVT U3543 ( .A1(n7676), .A2(n7675), .A3(n7674), .A4(n7673), .Y(n2369)
         );
  AO21X2_LVT U3544 ( .A1(n2368), .A2(n2369), .A3(n3631), .Y(n7681) );
  HADDX1_LVT U3545 ( .A0(n3104), .B0(n5405), .SO(n2370) );
  NAND2X0_LVT U3546 ( .A1(n2370), .A2(n3251), .Y(n5409) );
  INVX0_LVT U3547 ( .A(ibuf_io_pc[37]), .Y(n2371) );
  INVX0_LVT U3548 ( .A(n9494), .Y(n2372) );
  AO22X1_LVT U3549 ( .A1(ibuf_io_pc[37]), .A2(n9494), .A3(n2371), .A4(n2372), 
        .Y(n4577) );
  AO22X1_LVT U3550 ( .A1(io_fpu_dmem_resp_data[30]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[30]), .A4(n9065), .Y(n2373) );
  AO22X1_LVT U3551 ( .A1(n_T_628[30]), .A2(n2493), .A3(n_T_918[30]), .A4(n9066), .Y(n2374) );
  OR2X1_LVT U3552 ( .A1(n2373), .A2(n2374), .Y(io_fpu_fromint_data[30]) );
  AND2X1_LVT U3553 ( .A1(n_T_1187[28]), .A2(n2572), .Y(n2375) );
  NAND2X0_LVT U3554 ( .A1(n5367), .A2(n5314), .Y(n2376) );
  AO22X1_LVT U3555 ( .A1(n5366), .A2(n5317), .A3(n2375), .A4(n2376), .Y(N774)
         );
  AO222X1_LVT U3556 ( .A1(n_T_702[3]), .A2(n2515), .A3(n_T_702[19]), .A4(n9301), .A5(n4058), .A6(n_T_702[51]), .Y(N512) );
  AO222X1_LVT U3557 ( .A1(mem_br_target[12]), .A2(n6249), .A3(n_T_918[12]), 
        .A4(n6855), .A5(io_fpu_toint_data[12]), .A6(n6856), .Y(N610) );
  AOI22X1_LVT U3558 ( .A1(n_T_918[57]), .A2(n6855), .A3(io_fpu_toint_data[57]), 
        .A4(n6856), .Y(n2377) );
  NAND2X0_LVT U3559 ( .A1(n6857), .A2(n2377), .Y(N655) );
  INVX0_LVT U3560 ( .A(n5095), .Y(n2378) );
  AO221X1_LVT U3561 ( .A1(n5064), .A2(io_dmem_s2_nack), .A3(n5064), .A4(
        blocked), .A5(n2378), .Y(n2379) );
  AND2X1_LVT U3562 ( .A1(n5065), .A2(n2379), .Y(N811) );
  INVX0_LVT U3563 ( .A(n5191), .Y(n2380) );
  NAND3X0_LVT U3564 ( .A1(n5185), .A2(n5184), .A3(n2380), .Y(n5280) );
  INVX0_LVT U3565 ( .A(n5428), .Y(n2381) );
  AND2X1_LVT U3566 ( .A1(n2381), .A2(n5426), .Y(n5328) );
  AO22X1_LVT U3567 ( .A1(n3713), .A2(n_T_427[171]), .A3(n_T_427[555]), .A4(
        n3788), .Y(n8328) );
  AO22X1_LVT U3568 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[16]), .A3(n6899), 
        .A4(n_T_918[16]), .Y(n2382) );
  AO22X1_LVT U3569 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[16]), .A3(n6901), 
        .A4(n_T_635[16]), .Y(n2383) );
  OR2X1_LVT U3570 ( .A1(n2382), .A2(n2383), .Y(n_T_702[16]) );
  AO22X1_LVT U3571 ( .A1(io_fpu_dmem_resp_data[7]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[7]), .A4(n9065), .Y(n2384) );
  AO22X1_LVT U3572 ( .A1(n_T_628[7]), .A2(n2493), .A3(n_T_918[7]), .A4(n9066), 
        .Y(n2385) );
  OR2X1_LVT U3573 ( .A1(n2384), .A2(n2385), .Y(io_fpu_fromint_data[7]) );
  INVX0_LVT U3574 ( .A(io_dmem_s2_nack), .Y(n2386) );
  AND3X1_LVT U3575 ( .A1(wb_reg_valid), .A2(wb_ctrl_fence_i), .A3(n2386), .Y(
        io_imem_flush_icache) );
  NAND2X0_LVT U3576 ( .A1(n_T_427[1630]), .A2(n3652), .Y(n2387) );
  AND3X1_LVT U3577 ( .A1(n2387), .A2(n7881), .A3(n7882), .Y(n2388) );
  AND4X1_LVT U3578 ( .A1(n7879), .A2(n2388), .A3(n7878), .A4(n7877), .Y(n2389)
         );
  NAND4X0_LVT U3579 ( .A1(n3054), .A2(n2389), .A3(n3055), .A4(n3056), .Y(N711)
         );
  AO222X1_LVT U3580 ( .A1(n9296), .A2(n2515), .A3(n_T_702[26]), .A4(n9301), 
        .A5(n4058), .A6(n_T_702[58]), .Y(N519) );
  NAND2X0_LVT U3581 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[3]), .Y(n2390) );
  NAND4X0_LVT U3582 ( .A1(n9157), .A2(n9155), .A3(n9156), .A4(n2390), .Y(
        n_T_702[3]) );
  AO222X1_LVT U3583 ( .A1(n6249), .A2(mem_br_target[17]), .A3(n_T_918[17]), 
        .A4(n6855), .A5(io_fpu_toint_data[17]), .A6(n6856), .Y(N615) );
  AOI22X1_LVT U3584 ( .A1(n_T_918[63]), .A2(n6855), .A3(io_fpu_toint_data[63]), 
        .A4(n6856), .Y(n2391) );
  NAND2X0_LVT U3585 ( .A1(n6857), .A2(n2391), .Y(N661) );
  OA221X1_LVT U3586 ( .A1(n5396), .A2(io_fpu_inst[26]), .A3(n5396), .A4(n1847), 
        .A5(n2873), .Y(n2392) );
  INVX0_LVT U3587 ( .A(n5063), .Y(n2393) );
  OA221X1_LVT U3588 ( .A1(n2392), .A2(id_reg_fence), .A3(n2393), .A4(n2392), 
        .A5(n4498), .Y(n1821) );
  INVX0_LVT U3589 ( .A(ibuf_io_pc[30]), .Y(n2394) );
  INVX0_LVT U3590 ( .A(n9492), .Y(n2395) );
  AO22X1_LVT U3591 ( .A1(ibuf_io_pc[30]), .A2(n9492), .A3(n2394), .A4(n2395), 
        .Y(n4587) );
  AOI22X1_LVT U3592 ( .A1(n3745), .A2(n_T_427[246]), .A3(n3771), .A4(
        n_T_427[757]), .Y(n3719) );
  AO22X1_LVT U3593 ( .A1(io_fpu_dmem_resp_data[13]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[13]), .A4(n9065), .Y(n2396) );
  AO22X1_LVT U3594 ( .A1(n_T_628[13]), .A2(n2493), .A3(n_T_918[13]), .A4(n9066), .Y(n2397) );
  OR2X1_LVT U3595 ( .A1(n2396), .A2(n2397), .Y(io_fpu_fromint_data[13]) );
  INVX0_LVT U3596 ( .A(csr_io_interrupt_cause[3]), .Y(n2398) );
  OA21X1_LVT U3597 ( .A1(n9448), .A2(n2398), .A3(n74), .Y(n2507) );
  OA22X1_LVT U3598 ( .A1(n5237), .A2(n5292), .A3(n5295), .A4(n5238), .Y(n2399)
         );
  AO22X1_LVT U3599 ( .A1(n3793), .A2(n_T_1298[11]), .A3(n5298), .A4(n5239), 
        .Y(n2400) );
  AND2X1_LVT U3600 ( .A1(n2399), .A2(n2400), .Y(N790) );
  NAND2X0_LVT U3601 ( .A1(n_T_427[1627]), .A2(n3651), .Y(n2401) );
  AND3X1_LVT U3602 ( .A1(n2401), .A2(n7793), .A3(n7794), .Y(n2402) );
  AND4X1_LVT U3603 ( .A1(n7791), .A2(n2402), .A3(n7790), .A4(n7789), .Y(n2403)
         );
  NAND4X0_LVT U3604 ( .A1(n3051), .A2(n2403), .A3(n3052), .A4(n3053), .Y(N708)
         );
  AO222X1_LVT U3605 ( .A1(n_T_702[4]), .A2(n2515), .A3(n_T_702[20]), .A4(n9301), .A5(n4058), .A6(n_T_702[52]), .Y(N513) );
  AO22X1_LVT U3606 ( .A1(n6813), .A2(n_T_427[842]), .A3(n2826), .A4(
        n_T_427[11]), .Y(n2404) );
  OAI22X1_LVT U3607 ( .A1(n3879), .A2(n5681), .A3(n3186), .A4(n3596), .Y(n2405) );
  NOR4X0_LVT U3608 ( .A1(n5676), .A2(n5675), .A3(n2404), .A4(n2405), .Y(n2406)
         );
  AOI22X1_LVT U3609 ( .A1(n3827), .A2(n_T_427[1674]), .A3(n3890), .A4(
        n_T_427[1546]), .Y(n2407) );
  AOI22X1_LVT U3610 ( .A1(n3922), .A2(n_T_427[1482]), .A3(n_T_427[1610]), .A4(
        n3889), .Y(n2408) );
  AOI22X2_LVT U3611 ( .A1(n3828), .A2(n_T_427[1801]), .A3(n_T_427[1738]), .A4(
        n2866), .Y(n2409) );
  AND4X1_LVT U3612 ( .A1(n2407), .A2(n2750), .A3(n2409), .A4(n2408), .Y(n2410)
         );
  AO22X1_LVT U3613 ( .A1(n3932), .A2(n_T_427[1418]), .A3(n_T_427[1354]), .A4(
        n3921), .Y(n2411) );
  AO22X1_LVT U3614 ( .A1(n3942), .A2(n_T_427[1162]), .A3(n_T_427[1290]), .A4(
        n3931), .Y(n2412) );
  AO22X1_LVT U3615 ( .A1(n3952), .A2(n_T_427[1098]), .A3(n_T_427[1226]), .A4(
        n3941), .Y(n2413) );
  AO22X1_LVT U3616 ( .A1(n3898), .A2(n_T_427[1034]), .A3(n_T_427[970]), .A4(
        n3951), .Y(n2414) );
  NOR4X0_LVT U3617 ( .A1(n2411), .A2(n2412), .A3(n2413), .A4(n2414), .Y(n2415)
         );
  NAND2X0_LVT U3618 ( .A1(n3819), .A2(n_T_427[523]), .Y(n2416) );
  NAND4X0_LVT U3619 ( .A1(n2406), .A2(n2410), .A3(n2415), .A4(n2416), .Y(
        id_rs_1[11]) );
  AO222X1_LVT U3620 ( .A1(n6249), .A2(mem_br_target[19]), .A3(n_T_918[19]), 
        .A4(n6855), .A5(io_fpu_toint_data[19]), .A6(n6856), .Y(N617) );
  AOI22X1_LVT U3621 ( .A1(n_T_918[58]), .A2(n6855), .A3(io_fpu_toint_data[58]), 
        .A4(n6856), .Y(n2417) );
  NAND2X0_LVT U3622 ( .A1(n6857), .A2(n2417), .Y(N656) );
  INVX0_LVT U3623 ( .A(n4507), .Y(n2418) );
  OA22X1_LVT U3624 ( .A1(io_fpu_inst[5]), .A2(n9109), .A3(io_fpu_inst[13]), 
        .A4(n2418), .Y(n2419) );
  AOI22X1_LVT U3625 ( .A1(io_fpu_inst[5]), .A2(n3077), .A3(n2552), .A4(n5067), 
        .Y(n2420) );
  NAND2X0_LVT U3626 ( .A1(n2639), .A2(n5074), .Y(n2421) );
  NAND4X0_LVT U3627 ( .A1(n5174), .A2(n2419), .A3(n2420), .A4(n2421), .Y(
        id_ctrl_wxd) );
  OR4X1_LVT U3628 ( .A1(ex_ctrl_div), .A2(ex_ctrl_csr[0]), .A3(ex_ctrl_csr[2]), 
        .A4(io_dmem_req_bits_tag[0]), .Y(n2422) );
  NOR4X0_LVT U3629 ( .A1(ex_ctrl_mem), .A2(ex_ctrl_jalr), .A3(ex_ctrl_csr[1]), 
        .A4(n2422), .Y(n5051) );
  INVX0_LVT U3630 ( .A(n5191), .Y(n2423) );
  NAND3X0_LVT U3631 ( .A1(n5185), .A2(io_fpu_dmem_resp_tag[0]), .A3(n2423), 
        .Y(n5270) );
  AND3X1_LVT U3632 ( .A1(n5481), .A2(ex_reg_rs_bypass_1), .A3(n5483), .Y(n6899) );
  AO222X1_LVT U3633 ( .A1(n3851), .A2(io_dmem_resp_bits_data[11]), .A3(
        div_io_resp_bits_data[11]), .A4(n3854), .A5(n3850), .A6(
        io_imem_sfence_bits_addr[11]), .Y(n2424) );
  AOI21X1_LVT U3634 ( .A1(csr_io_rw_rdata[11]), .A2(n3842), .A3(n2424), .Y(
        n3186) );
  AO22X1_LVT U3635 ( .A1(io_fpu_dmem_resp_data[15]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[15]), .A4(n9065), .Y(n2425) );
  AO22X1_LVT U3636 ( .A1(n_T_628[15]), .A2(n2493), .A3(n_T_918[15]), .A4(n9066), .Y(n2426) );
  OR2X1_LVT U3637 ( .A1(n2425), .A2(n2426), .Y(io_fpu_fromint_data[15]) );
  AND4X1_LVT U3638 ( .A1(n2927), .A2(n3677), .A3(n2926), .A4(n3676), .Y(n2427)
         );
  NAND3X0_LVT U3639 ( .A1(n3779), .A2(n2427), .A3(n3690), .Y(N715) );
  AO222X1_LVT U3640 ( .A1(n_T_702[2]), .A2(n2515), .A3(n_T_702[18]), .A4(n9301), .A5(n4058), .A6(n_T_702[50]), .Y(N511) );
  AND4X1_LVT U3641 ( .A1(n2841), .A2(n2840), .A3(n2839), .A4(n2838), .Y(n2428)
         );
  AO22X1_LVT U3642 ( .A1(n3928), .A2(n_T_427[1298]), .A3(n_T_427[1426]), .A4(
        n3934), .Y(n2430) );
  AO22X1_LVT U3643 ( .A1(n3938), .A2(n_T_427[1234]), .A3(n_T_427[1170]), .A4(
        n3944), .Y(n2431) );
  AO22X1_LVT U3644 ( .A1(n3948), .A2(n_T_427[978]), .A3(n_T_427[1106]), .A4(
        n3954), .Y(n2432) );
  AO22X1_LVT U3645 ( .A1(n2830), .A2(n_T_427[211]), .A3(n_T_427[1042]), .A4(
        n3900), .Y(n2433) );
  NOR4X0_LVT U3646 ( .A1(n2430), .A2(n2431), .A3(n2432), .A4(n2433), .Y(n2434)
         );
  NAND3X0_LVT U3647 ( .A1(n2428), .A2(n2429), .A3(n2434), .Y(id_rs_1[19]) );
  AO222X1_LVT U3648 ( .A1(n6249), .A2(mem_br_target[14]), .A3(n_T_918[14]), 
        .A4(n6855), .A5(io_fpu_toint_data[14]), .A6(n6856), .Y(N612) );
  AO222X1_LVT U3649 ( .A1(n6249), .A2(mem_br_target[25]), .A3(n_T_918[25]), 
        .A4(n6855), .A5(io_fpu_toint_data[25]), .A6(n6856), .Y(N623) );
  AOI22X1_LVT U3650 ( .A1(n_T_918[59]), .A2(n6855), .A3(io_fpu_toint_data[59]), 
        .A4(n6856), .Y(n2435) );
  NAND2X0_LVT U3651 ( .A1(n6857), .A2(n2435), .Y(N657) );
  AOI21X1_LVT U3652 ( .A1(io_dmem_req_bits_cmd[1]), .A2(n560), .A3(n5078), .Y(
        n2436) );
  OA221X1_LVT U3653 ( .A1(io_dmem_req_bits_cmd[3]), .A2(
        io_dmem_req_bits_cmd[2]), .A3(io_dmem_req_bits_cmd[3]), .A4(n2436), 
        .A5(n3245), .Y(n997) );
  INVX0_LVT U3654 ( .A(n5169), .Y(n2437) );
  AO22X1_LVT U3655 ( .A1(io_imem_req_bits_speculative), .A2(mem_reg_replay), 
        .A3(io_imem_bht_update_valid), .A4(n2437), .Y(N530) );
  INVX0_LVT U3656 ( .A(io_fpu_sboard_clra[3]), .Y(n2438) );
  AND2X1_LVT U3657 ( .A1(n2438), .A2(io_fpu_sboard_clra[4]), .Y(n5258) );
  INVX0_LVT U3658 ( .A(io_fpu_sboard_clra[4]), .Y(n2439) );
  NAND2X0_LVT U3659 ( .A1(io_fpu_sboard_clra[3]), .A2(n2439), .Y(n5245) );
  AO22X1_LVT U3660 ( .A1(io_fpu_dmem_resp_data[10]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[10]), .A4(n9065), .Y(n2440) );
  AO22X1_LVT U3661 ( .A1(n_T_628[10]), .A2(n2497), .A3(n_T_918[10]), .A4(n9066), .Y(n2441) );
  OR2X1_LVT U3662 ( .A1(n2440), .A2(n2441), .Y(io_fpu_fromint_data[10]) );
  NAND2X0_LVT U3663 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[4]), .Y(n2442) );
  NAND4X0_LVT U3664 ( .A1(n9161), .A2(n9159), .A3(n9160), .A4(n2442), .Y(
        n_T_702[4]) );
  AO222X1_LVT U3665 ( .A1(n_T_702[0]), .A2(n2515), .A3(n_T_702[16]), .A4(n9301), .A5(n4058), .A6(n_T_702[48]), .Y(N509) );
  NAND2X0_LVT U3666 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[2]), .Y(n2443) );
  NAND4X0_LVT U3667 ( .A1(n9150), .A2(n9148), .A3(n9149), .A4(n2443), .Y(
        n_T_702[2]) );
  AO22X1_LVT U3668 ( .A1(n3932), .A2(n_T_427[1432]), .A3(n_T_427[1368]), .A4(
        n3921), .Y(n2444) );
  AO22X1_LVT U3669 ( .A1(n3942), .A2(n_T_427[1176]), .A3(n_T_427[1304]), .A4(
        n3931), .Y(n2445) );
  AO22X1_LVT U3670 ( .A1(n3952), .A2(n_T_427[1112]), .A3(n_T_427[1240]), .A4(
        n3941), .Y(n2446) );
  AO22X1_LVT U3671 ( .A1(n3898), .A2(n_T_427[1048]), .A3(n_T_427[984]), .A4(
        n3951), .Y(n2447) );
  NOR4X0_LVT U3672 ( .A1(n2444), .A2(n2445), .A3(n2446), .A4(n2447), .Y(n2448)
         );
  AO22X1_LVT U3673 ( .A1(n3922), .A2(n_T_427[1496]), .A3(n_T_427[1624]), .A4(
        n3889), .Y(n2449) );
  NOR4X0_LVT U3674 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n2449), .Y(n2450)
         );
  NOR4X0_LVT U3675 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .Y(n2451)
         );
  NAND3X0_LVT U3676 ( .A1(n2448), .A2(n2450), .A3(n2451), .Y(id_rs_1[25]) );
  AO222X1_LVT U3677 ( .A1(mem_br_target[8]), .A2(n6249), .A3(n_T_918[8]), .A4(
        n6855), .A5(io_fpu_toint_data[8]), .A6(n6856), .Y(N606) );
  AO222X1_LVT U3678 ( .A1(n6249), .A2(mem_br_target[15]), .A3(n_T_918[15]), 
        .A4(n6855), .A5(io_fpu_toint_data[15]), .A6(n6856), .Y(N613) );
  AO222X1_LVT U3679 ( .A1(mem_br_target[21]), .A2(n6249), .A3(n_T_918[21]), 
        .A4(n6855), .A5(io_fpu_toint_data[21]), .A6(n6856), .Y(N619) );
  AO222X1_LVT U3680 ( .A1(n6249), .A2(mem_br_target[27]), .A3(n_T_918[27]), 
        .A4(n6855), .A5(io_fpu_toint_data[27]), .A6(n6856), .Y(N625) );
  AOI22X1_LVT U3681 ( .A1(n_T_918[60]), .A2(n6855), .A3(io_fpu_toint_data[60]), 
        .A4(n6856), .Y(n2452) );
  NAND2X0_LVT U3682 ( .A1(n6857), .A2(n2452), .Y(N658) );
  OA221X1_LVT U3683 ( .A1(n1853), .A2(n3597), .A3(io_fpu_inst[3]), .A4(n9445), 
        .A5(n9109), .Y(n2453) );
  NOR2X0_LVT U3684 ( .A1(n1431), .A2(n2453), .Y(N275) );
  INVX0_LVT U3685 ( .A(io_imem_req_bits_speculative), .Y(n2454) );
  AOI221X1_LVT U3686 ( .A1(mem_reg_valid), .A2(mem_reg_sfence), .A3(
        mem_reg_valid), .A4(io_imem_bht_update_bits_mispredict), .A5(n2454), 
        .Y(n9418) );
  NAND2X0_LVT U3687 ( .A1(n118), .A2(n9361), .Y(n2455) );
  OA221X1_LVT U3688 ( .A1(n9501), .A2(n_T_698[22]), .A3(n118), .A4(n9361), 
        .A5(n2455), .Y(n4603) );
  INVX0_LVT U3689 ( .A(n5191), .Y(n2456) );
  NAND3X0_LVT U3690 ( .A1(io_fpu_dmem_resp_tag[1]), .A2(n5184), .A3(n2456), 
        .Y(n5261) );
  AO22X1_LVT U3691 ( .A1(io_fpu_dmem_resp_data[14]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[14]), .A4(n9065), .Y(n2457) );
  AO22X1_LVT U3692 ( .A1(n_T_628[14]), .A2(n2497), .A3(n_T_918[14]), .A4(n9066), .Y(n2458) );
  OR2X1_LVT U3693 ( .A1(n2457), .A2(n2458), .Y(io_fpu_fromint_data[14]) );
  AND2X1_LVT U3694 ( .A1(n_T_1187[29]), .A2(n2572), .Y(n2459) );
  NAND2X0_LVT U3695 ( .A1(n5385), .A2(n5314), .Y(n2460) );
  AO22X1_LVT U3696 ( .A1(n5383), .A2(n5317), .A3(n2459), .A4(n2460), .Y(N775)
         );
  OR4X1_LVT U3697 ( .A1(n8059), .A2(n8077), .A3(n8079), .A4(n8060), .Y(n2461)
         );
  AO222X1_LVT U3698 ( .A1(n_T_702[17]), .A2(n9301), .A3(n_T_702[1]), .A4(n2515), .A5(n4058), .A6(n_T_702[49]), .Y(N510) );
  AO222X1_LVT U3699 ( .A1(n6249), .A2(mem_br_target[9]), .A3(n_T_918[9]), .A4(
        n6855), .A5(io_fpu_toint_data[9]), .A6(n6856), .Y(N607) );
  AO222X1_LVT U3700 ( .A1(n6249), .A2(mem_br_target[16]), .A3(n_T_918[16]), 
        .A4(n6855), .A5(io_fpu_toint_data[16]), .A6(n6856), .Y(N614) );
  AO222X1_LVT U3701 ( .A1(n6249), .A2(mem_br_target[23]), .A3(n_T_918[23]), 
        .A4(n6855), .A5(io_fpu_toint_data[23]), .A6(n6856), .Y(N621) );
  AO222X1_LVT U3702 ( .A1(n6249), .A2(mem_br_target[29]), .A3(n_T_918[29]), 
        .A4(n6855), .A5(io_fpu_toint_data[29]), .A6(n6856), .Y(N627) );
  AO222X1_LVT U3703 ( .A1(n6249), .A2(mem_br_target[34]), .A3(n_T_918[34]), 
        .A4(n6855), .A5(io_fpu_toint_data[34]), .A6(n6856), .Y(N632) );
  AOI22X1_LVT U3704 ( .A1(n_T_918[61]), .A2(n6855), .A3(io_fpu_toint_data[61]), 
        .A4(n6856), .Y(n2462) );
  NAND2X0_LVT U3705 ( .A1(n6857), .A2(n2462), .Y(N659) );
  AOI22X1_LVT U3706 ( .A1(n5123), .A2(n5087), .A3(csr_io_decode_0_write_flush), 
        .A4(n5088), .Y(n2463) );
  INVX0_LVT U3707 ( .A(n1828), .Y(n2464) );
  NAND3X0_LVT U3708 ( .A1(n2463), .A2(n5122), .A3(n2464), .Y(n_T_731) );
  INVX0_LVT U3709 ( .A(div_io_req_ready), .Y(n2465) );
  NAND2X0_LVT U3710 ( .A1(n9422), .A2(n2465), .Y(n2466) );
  NAND3X0_LVT U3711 ( .A1(ex_reg_valid), .A2(n5175), .A3(ex_reg_load_use), .Y(
        n2467) );
  AND4X1_LVT U3712 ( .A1(n3233), .A2(n5095), .A3(n2466), .A4(n2467), .Y(n9421)
         );
  OA22X2_LVT U3713 ( .A1(n3803), .A2(n3170), .A3(n3488), .A4(n3800), .Y(n2468)
         );
  OA22X1_LVT U3714 ( .A1(n3082), .A2(n3489), .A3(n3081), .A4(n3171), .Y(n2469)
         );
  AOI22X1_LVT U3715 ( .A1(n3894), .A2(n_T_427[1598]), .A3(n_T_427[1662]), .A4(
        n3889), .Y(n2470) );
  AND4X1_LVT U3716 ( .A1(n2468), .A2(n6881), .A3(n2470), .A4(n2469), .Y(n2471)
         );
  AO22X1_LVT U3717 ( .A1(n3909), .A2(n_T_427[191]), .A3(n3911), .A4(
        n_T_427[511]), .Y(n2472) );
  AO22X1_LVT U3718 ( .A1(n3916), .A2(n_T_427[639]), .A3(n_T_427[63]), .A4(
        n3913), .Y(n2473) );
  AO22X1_LVT U3719 ( .A1(n3899), .A2(n_T_427[1086]), .A3(n_T_427[958]), .A4(
        n2831), .Y(n2474) );
  AO22X1_LVT U3720 ( .A1(n3905), .A2(n_T_427[766]), .A3(n_T_427[830]), .A4(
        n2861), .Y(n2475) );
  NOR4X0_LVT U3721 ( .A1(n2472), .A2(n2473), .A3(n2474), .A4(n2475), .Y(n2476)
         );
  AO22X1_LVT U3722 ( .A1(n3922), .A2(n_T_427[1534]), .A3(n_T_427[1406]), .A4(
        n3917), .Y(n2477) );
  AO22X1_LVT U3723 ( .A1(n3933), .A2(n_T_427[1470]), .A3(n_T_427[1342]), .A4(
        n3927), .Y(n2478) );
  AO22X1_LVT U3724 ( .A1(n3942), .A2(n_T_427[1214]), .A3(n_T_427[1278]), .A4(
        n3937), .Y(n2479) );
  AO22X1_LVT U3725 ( .A1(n3952), .A2(n_T_427[1150]), .A3(n_T_427[1022]), .A4(
        n3947), .Y(n2480) );
  NOR4X0_LVT U3726 ( .A1(n2477), .A2(n2478), .A3(n2479), .A4(n2480), .Y(n2481)
         );
  NAND2X0_LVT U3727 ( .A1(n4496), .A2(n3959), .Y(n2482) );
  NAND4X0_LVT U3728 ( .A1(n2471), .A2(n2476), .A3(n2481), .A4(n2482), .Y(
        id_rs_1[63]) );
  INVX0_LVT U3729 ( .A(io_fpu_sboard_clra[1]), .Y(n2483) );
  AND2X1_LVT U3730 ( .A1(n2483), .A2(io_fpu_sboard_clr), .Y(n5183) );
  NAND2X0_LVT U3731 ( .A1(n_T_427[59]), .A2(n8944), .Y(n2484) );
  NAND3X0_LVT U3732 ( .A1(n2484), .A2(n8887), .A3(n8886), .Y(n2582) );
  OAI21X1_LVT U3733 ( .A1(n2968), .A2(n1262), .A3(n9412), .Y(n9383) );
  INVX0_LVT U3734 ( .A(n5191), .Y(n2485) );
  NAND3X0_LVT U3735 ( .A1(io_fpu_dmem_resp_tag[0]), .A2(
        io_fpu_dmem_resp_tag[1]), .A3(n2485), .Y(n5292) );
  AO22X1_LVT U3736 ( .A1(io_fpu_dmem_resp_data[11]), .A2(n9064), .A3(
        io_imem_sfence_bits_addr[11]), .A4(n9065), .Y(n2486) );
  AO22X1_LVT U3737 ( .A1(n_T_628[11]), .A2(n2493), .A3(n_T_918[11]), .A4(n9066), .Y(n2487) );
  OR2X1_LVT U3738 ( .A1(n2486), .A2(n2487), .Y(io_fpu_fromint_data[11]) );
  AND3X1_LVT U3739 ( .A1(n9179), .A2(n9173), .A3(n9200), .Y(n9199) );
  AO222X1_LVT U3740 ( .A1(n_T_702[21]), .A2(n9301), .A3(n_T_702[5]), .A4(n2515), .A5(n4058), .A6(n_T_702[53]), .Y(N514) );
  INVX0_LVT U3741 ( .A(n5483), .Y(n2488) );
  NAND2X0_LVT U3742 ( .A1(io_fpu_dmem_resp_data[1]), .A2(n2488), .Y(n2489) );
  NAND4X0_LVT U3743 ( .A1(n9135), .A2(n9136), .A3(n9137), .A4(n2489), .Y(
        n_T_702[1]) );
  AO222X1_LVT U3744 ( .A1(n6249), .A2(mem_br_target[10]), .A3(n_T_918[10]), 
        .A4(n6855), .A5(io_fpu_toint_data[10]), .A6(n6856), .Y(N608) );
  AO222X1_LVT U3745 ( .A1(n6249), .A2(mem_br_target[18]), .A3(n_T_918[18]), 
        .A4(n6855), .A5(io_fpu_toint_data[18]), .A6(n6856), .Y(N616) );
  AO222X1_LVT U3746 ( .A1(n6249), .A2(mem_br_target[20]), .A3(n_T_918[20]), 
        .A4(n6855), .A5(io_fpu_toint_data[20]), .A6(n6856), .Y(N618) );
  AO222X1_LVT U3747 ( .A1(mem_br_target[22]), .A2(n6249), .A3(n_T_918[22]), 
        .A4(n6855), .A5(io_fpu_toint_data[22]), .A6(n6856), .Y(N620) );
  AO222X1_LVT U3748 ( .A1(n6249), .A2(mem_br_target[24]), .A3(n_T_918[24]), 
        .A4(n6855), .A5(io_fpu_toint_data[24]), .A6(n6856), .Y(N622) );
  AO222X1_LVT U3749 ( .A1(n6249), .A2(mem_br_target[26]), .A3(n_T_918[26]), 
        .A4(n6855), .A5(io_fpu_toint_data[26]), .A6(n6856), .Y(N624) );
  AO222X1_LVT U3750 ( .A1(n6249), .A2(mem_br_target[28]), .A3(n_T_918[28]), 
        .A4(n6855), .A5(io_fpu_toint_data[28]), .A6(n6856), .Y(N626) );
  AO222X1_LVT U3751 ( .A1(n6249), .A2(mem_br_target[30]), .A3(n_T_918[30]), 
        .A4(n6855), .A5(io_fpu_toint_data[30]), .A6(n6856), .Y(N628) );
  AO222X1_LVT U3752 ( .A1(n6249), .A2(mem_br_target[36]), .A3(n_T_918[36]), 
        .A4(n6855), .A5(io_fpu_toint_data[36]), .A6(n6856), .Y(N634) );
  AO222X1_LVT U3753 ( .A1(n6249), .A2(mem_br_target[37]), .A3(n_T_918[37]), 
        .A4(n6855), .A5(io_fpu_toint_data[37]), .A6(n6856), .Y(N635) );
  AOI22X1_LVT U3754 ( .A1(n_T_918[62]), .A2(n6855), .A3(io_fpu_toint_data[62]), 
        .A4(n6856), .Y(n2490) );
  NAND2X0_LVT U3755 ( .A1(n6857), .A2(n2490), .Y(N660) );
  AO221X1_LVT U3756 ( .A1(n1853), .A2(io_fpu_inst[31]), .A3(n1853), .A4(n5099), 
        .A5(io_fpu_inst[6]), .Y(id_ctrl_mem_cmd_2_) );
  IBUFFX2_LVT U3757 ( .A(n3081), .Y(n2765) );
  IBUFFX2_LVT U3758 ( .A(n3081), .Y(n3830) );
  IBUFFX2_LVT U3759 ( .A(n3081), .Y(n3828) );
  IBUFFX2_LVT U3760 ( .A(n3081), .Y(n3829) );
  IBUFFX2_LVT U3761 ( .A(n6765), .Y(n3805) );
  AND2X4_LVT U3762 ( .A1(n5453), .A2(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(
        n6765) );
  IBUFFX2_LVT U3763 ( .A(n3805), .Y(n3804) );
  IBUFFX2_LVT U3764 ( .A(n3012), .Y(n9008) );
  DELLN1X2_LVT U3765 ( .A(n3803), .Y(n2875) );
  IBUFFX2_LVT U3766 ( .A(n3186), .Y(n4351) );
  AOI21X2_LVT U3767 ( .A1(n3841), .A2(csr_io_rw_rdata[4]), .A3(n5529), .Y(
        n3190) );
  IBUFFX2_LVT U3768 ( .A(n3190), .Y(n4330) );
  IBUFFX2_LVT U3769 ( .A(n3692), .Y(n3989) );
  IBUFFX2_LVT U3770 ( .A(n3692), .Y(n2969) );
  IBUFFX2_LVT U3771 ( .A(n3692), .Y(n3988) );
  IBUFFX2_LVT U3772 ( .A(n6871), .Y(n3876) );
  AND2X4_LVT U3773 ( .A1(n5449), .A2(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(
        n6871) );
  IBUFFX2_LVT U3774 ( .A(n3876), .Y(n3875) );
  IBUFFX2_LVT U3775 ( .A(n3876), .Y(n3874) );
  IBUFFX2_LVT U3776 ( .A(n3783), .Y(n2552) );
  IBUFFX2_LVT U3777 ( .A(n9524), .Y(n9446) );
  NBUFFX2_LVT U3778 ( .A(n9036), .Y(n3060) );
  NBUFFX2_LVT U3779 ( .A(n9036), .Y(n2982) );
  IBUFFX2_LVT U3780 ( .A(n3184), .Y(n4023) );
  IBUFFX2_LVT U3781 ( .A(n3184), .Y(n4025) );
  IBUFFX2_LVT U3782 ( .A(n3184), .Y(n4024) );
  IBUFFX2_LVT U3783 ( .A(n6422), .Y(n6866) );
  DELLN1X2_LVT U3784 ( .A(n6866), .Y(n3864) );
  IBUFFX2_LVT U3785 ( .A(n6767), .Y(n6867) );
  DELLN1X2_LVT U3786 ( .A(n6867), .Y(n3865) );
  IBUFFX2_LVT U3787 ( .A(io_fpu_inst[12]), .Y(n3583) );
  IBUFFX2_LVT U3788 ( .A(clock), .Y(n3784) );
  DELLN1X2_LVT U3789 ( .A(n4499), .Y(n3594) );
  DELLN1X2_LVT U3790 ( .A(n4499), .Y(n3595) );
  INVX1_LVT U3791 ( .A(n3101), .Y(n2497) );
  INVX1_LVT U3792 ( .A(n3246), .Y(n2498) );
  AOI21X2_LVT U3793 ( .A1(io_fpu_inst[25]), .A2(n1847), .A3(n1828), .Y(n4855)
         );
  NAND3X2_LVT U3794 ( .A1(n9075), .A2(n9522), .A3(n9435), .Y(n4856) );
  NAND3X2_LVT U3795 ( .A1(io_fpu_inst[24]), .A2(n9522), .A3(io_fpu_inst[21]), 
        .Y(n5151) );
  AND2X1_LVT U3806 ( .A1(n1699), .A2(n3039), .Y(n2512) );
  AND2X1_LVT U3813 ( .A1(div_io_req_ready), .A2(n9422), .Y(n2524) );
  NBUFFX2_LVT U3814 ( .A(n2527), .Y(n2526) );
  NAND2X0_LVT U3815 ( .A1(n2527), .A2(n_T_427[424]), .Y(n8219) );
  NAND2X0_LVT U3816 ( .A1(n2527), .A2(n_T_427[436]), .Y(n2598) );
  NAND2X0_LVT U3817 ( .A1(n2527), .A2(n_T_427[429]), .Y(n8395) );
  NAND2X0_LVT U3818 ( .A1(n2527), .A2(n_T_427[446]), .Y(n8998) );
  NAND2X0_LVT U3819 ( .A1(n2527), .A2(n_T_427[441]), .Y(n8811) );
  NAND2X0_LVT U3820 ( .A1(n2527), .A2(n_T_427[423]), .Y(n8157) );
  NAND2X0_LVT U3821 ( .A1(n2527), .A2(n_T_427[417]), .Y(n7963) );
  NAND2X0_LVT U3822 ( .A1(n2527), .A2(n_T_427[437]), .Y(n8641) );
  NAND2X0_LVT U3823 ( .A1(n2526), .A2(n_T_427[432]), .Y(n8486) );
  NAND2X0_LVT U3824 ( .A1(n2526), .A2(n_T_427[419]), .Y(n8025) );
  NAND2X0_LVT U3825 ( .A1(n2526), .A2(n_T_427[421]), .Y(n8106) );
  NAND2X0_LVT U3826 ( .A1(n2526), .A2(n_T_427[438]), .Y(n8679) );
  AND2X4_LVT U3827 ( .A1(n8105), .A2(n3968), .Y(n2527) );
  NAND3X0_LVT U3828 ( .A1(n5142), .A2(n9437), .A3(n9443), .Y(n2528) );
  NAND2X0_LVT U3829 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[24]), .Y(n7683)
         );
  NAND2X0_LVT U3830 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[16]), .Y(n7442)
         );
  NAND2X0_LVT U3831 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[21]), .Y(n7591)
         );
  NAND2X0_LVT U3832 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[18]), .Y(n7499)
         );
  NAND2X0_LVT U3833 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[19]), .Y(n7532)
         );
  NAND2X0_LVT U3834 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[20]), .Y(n7559)
         );
  NAND2X0_LVT U3835 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[22]), .Y(n7622)
         );
  NAND2X0_LVT U3836 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[23]), .Y(n7655)
         );
  NAND2X0_LVT U3837 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[25]), .Y(n7718)
         );
  NAND2X0_LVT U3838 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[26]), .Y(n7751)
         );
  NAND2X0_LVT U3839 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[27]), .Y(n7783)
         );
  NAND2X0_LVT U3840 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[28]), .Y(n7815)
         );
  NAND2X0_LVT U3841 ( .A1(n2529), .A2(ibuf_io_inst_0_bits_raw[29]), .Y(n7848)
         );
  NAND2X0_LVT U3842 ( .A1(n2529), .A2(n1859), .Y(n7875) );
  NAND2X0_LVT U3843 ( .A1(n2529), .A2(n2494), .Y(n7903) );
  AND3X1_LVT U3844 ( .A1(n8943), .A2(n8945), .A3(n2531), .Y(n2530) );
  NAND2X0_LVT U3845 ( .A1(n3707), .A2(n_T_427[125]), .Y(n2531) );
  NAND4X0_LVT U3846 ( .A1(n2630), .A2(n2670), .A3(n9446), .A4(n9104), .Y(n2629) );
  AND2X4_LVT U3847 ( .A1(n3590), .A2(io_fpu_inst[6]), .Y(n5163) );
  AND3X1_LVT U3848 ( .A1(n6908), .A2(n6909), .A3(n6907), .Y(n2532) );
  OA21X1_LVT U3849 ( .A1(n9395), .A2(n9386), .A3(n9397), .Y(n9388) );
  AND3X1_LVT U3850 ( .A1(n3073), .A2(n6913), .A3(n6935), .Y(n6914) );
  NOR2X0_LVT U3851 ( .A1(n6910), .A2(n6911), .Y(n2533) );
  AND3X1_LVT U3852 ( .A1(n2534), .A2(n2535), .A3(n2536), .Y(n3737) );
  AND3X1_LVT U3853 ( .A1(n8627), .A2(n8626), .A3(n8625), .Y(n2534) );
  AND2X1_LVT U3854 ( .A1(n8632), .A2(n2617), .Y(n2535) );
  AND2X1_LVT U3855 ( .A1(n8629), .A2(n8628), .Y(n2536) );
  NAND2X0_LVT U3856 ( .A1(n4844), .A2(n4845), .Y(n2538) );
  NAND4X1_LVT U3857 ( .A1(n5162), .A2(n5161), .A3(n2624), .A4(n2623), .Y(n2539) );
  OR2X2_LVT U3858 ( .A1(n9524), .A2(n3078), .Y(n9079) );
  NAND3X1_LVT U3859 ( .A1(n5067), .A2(n9524), .A3(n9528), .Y(n1531) );
  OR2X2_LVT U3860 ( .A1(io_fpu_inst[12]), .A2(n9524), .Y(n5075) );
  NBUFFX2_LVT U3861 ( .A(n9521), .Y(io_fpu_inst[27]) );
  OR2X4_LVT U3862 ( .A1(n9520), .A2(n9521), .Y(n5099) );
  OA22X2_LVT U3863 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .Y(n5160)
         );
  NAND3X0_LVT U3864 ( .A1(n2541), .A2(n2542), .A3(n2543), .Y(N724) );
  AND4X1_LVT U3865 ( .A1(n2956), .A2(n2957), .A3(n8350), .A4(n2590), .Y(n2541)
         );
  AND3X1_LVT U3866 ( .A1(n8357), .A2(n8356), .A3(n8355), .Y(n2542) );
  AND3X2_LVT U3867 ( .A1(n6991), .A2(n9288), .A3(n6992), .Y(n2544) );
  OR2X2_LVT U3868 ( .A1(n9111), .A2(n5073), .Y(n5077) );
  AND2X4_LVT U3869 ( .A1(n6238), .A2(n5437), .Y(n5446) );
  AND2X4_LVT U3870 ( .A1(n6238), .A2(n5448), .Y(n5457) );
  NAND4X1_LVT U3871 ( .A1(n5433), .A2(n5430), .A3(n5432), .A4(n5431), .Y(n6238) );
  NAND3X0_LVT U3872 ( .A1(n6991), .A2(n9288), .A3(n6992), .Y(n1262) );
  NBUFFX2_LVT U3873 ( .A(n9527), .Y(io_fpu_inst[4]) );
  NAND2X0_LVT U3874 ( .A1(n_T_427[1899]), .A2(n3992), .Y(n7483) );
  AOI21X2_LVT U3875 ( .A1(n3039), .A2(n5069), .A3(n5068), .Y(n5123) );
  OR2X2_LVT U3876 ( .A1(n5099), .A2(n2568), .Y(n2669) );
  OA21X2_LVT U3877 ( .A1(n3276), .A2(n3993), .A3(n7934), .Y(n7937) );
  OR2X4_LVT U3878 ( .A1(n3531), .A2(n3993), .Y(n7077) );
  OR2X4_LVT U3879 ( .A1(n2496), .A2(n3993), .Y(n8352) );
  OR2X4_LVT U3880 ( .A1(n3277), .A2(n3993), .Y(n2593) );
  NAND2X0_LVT U3881 ( .A1(n3782), .A2(n3588), .Y(n9288) );
  NOR3X4_LVT U3882 ( .A1(io_fpu_inst[29]), .A2(n5130), .A3(io_fpu_inst[7]), 
        .Y(n5131) );
  AND4X2_LVT U3883 ( .A1(n9230), .A2(io_fpu_inst[6]), .A3(io_fpu_inst[29]), 
        .A4(n5136), .Y(n5137) );
  AND2X1_LVT U3884 ( .A1(n2544), .A2(n6906), .Y(n2548) );
  IBUFFX2_LVT U3885 ( .A(n9519), .Y(n9436) );
  NAND3X2_LVT U3886 ( .A1(n5138), .A2(n9445), .A3(io_fpu_inst[29]), .Y(n2641)
         );
  NAND3X2_LVT U3887 ( .A1(io_fpu_inst[29]), .A2(n3078), .A3(n9445), .Y(n5152)
         );
  NAND3X0_LVT U3888 ( .A1(n2549), .A2(n2550), .A3(n2551), .Y(N734) );
  AND3X1_LVT U3889 ( .A1(n8681), .A2(n8680), .A3(n8679), .Y(n2549) );
  AND3X1_LVT U3890 ( .A1(n3718), .A2(n3719), .A3(n3720), .Y(n2550) );
  NOR2X0_LVT U3891 ( .A1(n8705), .A2(n8706), .Y(n2551) );
  DELLN2X2_LVT U3892 ( .A(n9529), .Y(io_fpu_inst[2]) );
  AND2X4_LVT U3893 ( .A1(n9105), .A2(n9529), .Y(n9097) );
  AO21X2_LVT U3894 ( .A1(io_fpu_inst[13]), .A2(n9105), .A3(n9529), .Y(n5100)
         );
  NAND3X2_LVT U3895 ( .A1(io_dmem_resp_bits_replay), .A2(n2029), .A3(n2626), 
        .Y(n5403) );
  NAND2X0_LVT U3896 ( .A1(n4351), .A2(n3060), .Y(n2595) );
  DELLN3X2_LVT U3897 ( .A(n9036), .Y(n3665) );
  AND2X1_LVT U3898 ( .A1(n3765), .A2(n6923), .Y(n3773) );
  IBUFFX2_LVT U3899 ( .A(n5134), .Y(n5132) );
  NAND4X1_LVT U3900 ( .A1(n5166), .A2(n3049), .A3(n2130), .A4(io_fpu_inst[26]), 
        .Y(n6964) );
  NOR3X4_LVT U3901 ( .A1(n9438), .A2(n9110), .A3(n5129), .Y(n5070) );
  OR3X2_LVT U3902 ( .A1(io_fpu_inst[31]), .A2(io_fpu_inst[14]), .A3(n5129), 
        .Y(n5134) );
  AND2X1_LVT U3903 ( .A1(n6923), .A2(n6922), .Y(n6975) );
  IBUFFX2_LVT U3904 ( .A(n9518), .Y(n9435) );
  NBUFFX2_LVT U3905 ( .A(n9520), .Y(io_fpu_inst[28]) );
  OR2X2_LVT U3906 ( .A1(n8424), .A2(n3632), .Y(n8425) );
  NAND3X0_LVT U3907 ( .A1(n2555), .A2(n2556), .A3(n2557), .Y(N717) );
  AND3X1_LVT U3908 ( .A1(n2952), .A2(n2951), .A3(n2950), .Y(n2555) );
  AND3X1_LVT U3909 ( .A1(n8108), .A2(n8107), .A3(n8106), .Y(n2556) );
  NAND3X0_LVT U3910 ( .A1(n2558), .A2(n2559), .A3(n2560), .Y(N712) );
  AND3X1_LVT U3911 ( .A1(n7909), .A2(n7908), .A3(n7907), .Y(n2558) );
  AND3X1_LVT U3912 ( .A1(n7924), .A2(n7923), .A3(n7922), .Y(n2559) );
  AND3X1_LVT U3913 ( .A1(n2919), .A2(n2918), .A3(n2585), .Y(n2560) );
  AND2X1_LVT U3914 ( .A1(n6964), .A2(n2548), .Y(n6923) );
  NAND3X0_LVT U3915 ( .A1(n2562), .A2(n2563), .A3(n2564), .Y(N731) );
  AND3X1_LVT U3916 ( .A1(n8575), .A2(n8574), .A3(n8573), .Y(n2562) );
  AND3X1_LVT U3917 ( .A1(n3725), .A2(n3726), .A3(n3727), .Y(n2563) );
  NOR2X0_LVT U3918 ( .A1(n8600), .A2(n8599), .Y(n2564) );
  AND4X2_LVT U3919 ( .A1(n9442), .A2(n9438), .A3(n9441), .A4(n5148), .Y(n2565)
         );
  AO21X1_LVT U3920 ( .A1(n2629), .A2(n5108), .A3(n2669), .Y(n5165) );
  NAND3X1_LVT U3921 ( .A1(n9445), .A2(n3078), .A3(n2618), .Y(n3580) );
  NAND3X2_LVT U3922 ( .A1(n6995), .A2(n9288), .A3(n6992), .Y(n6944) );
  NAND3X1_LVT U3923 ( .A1(n6993), .A2(n572), .A3(n6992), .Y(n6994) );
  OR2X4_LVT U3924 ( .A1(n5051), .A2(n6992), .Y(n9281) );
  NAND4X1_LVT U3925 ( .A1(n4758), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .A3(
        n4757), .A4(n6963), .Y(n4759) );
  OA21X2_LVT U3926 ( .A1(n4996), .A2(n4995), .A3(n2825), .Y(n4997) );
  OR3X2_LVT U3927 ( .A1(n2878), .A2(ibuf_io_inst_0_bits_inst_rs2[4]), .A3(
        n5435), .Y(n5421) );
  AND2X1_LVT U3928 ( .A1(ibuf_io_inst_0_bits_inst_rs2[3]), .A2(
        ibuf_io_inst_0_bits_inst_rs2[4]), .Y(n5437) );
  XOR2X1_LVT U3929 ( .A1(n3782), .A2(n2566), .Y(n3581) );
  AND3X2_LVT U3930 ( .A1(n2068), .A2(n6957), .A3(n6975), .Y(n3769) );
  AND3X2_LVT U3931 ( .A1(n6975), .A2(n6954), .A3(n6973), .Y(n9015) );
  IBUFFX2_LVT U3932 ( .A(n9527), .Y(n3577) );
  AND4X1_LVT U3933 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n2625), .Y(n2567)
         );
  NAND4X1_LVT U3934 ( .A1(n9442), .A2(n9438), .A3(n9441), .A4(n5148), .Y(n5143) );
  AND3X2_LVT U3935 ( .A1(n9107), .A2(io_fpu_inst[5]), .A3(n9108), .Y(n1823) );
  AND3X2_LVT U3936 ( .A1(n2671), .A2(n2561), .A3(n6922), .Y(n3715) );
  NAND3X2_LVT U3937 ( .A1(n4857), .A2(io_fpu_inst[5]), .A3(n9104), .Y(n1532)
         );
  OR2X2_LVT U3938 ( .A1(io_fpu_inst[5]), .A2(io_fpu_inst[12]), .Y(n5133) );
  NAND3X2_LVT U3939 ( .A1(n9440), .A2(io_fpu_inst[4]), .A3(n9443), .Y(n5130)
         );
  NOR3X2_LVT U3940 ( .A1(n1262), .A2(n6935), .A3(n2968), .Y(n6937) );
  IBUFFX2_LVT U3941 ( .A(io_fpu_inst[26]), .Y(n9439) );
  AND2X4_LVT U3942 ( .A1(n2981), .A2(n6796), .Y(n6886) );
  AND2X4_LVT U3943 ( .A1(n6877), .A2(n3836), .Y(n6887) );
  AND2X4_LVT U3944 ( .A1(n6877), .A2(n3812), .Y(n6885) );
  AND2X4_LVT U3945 ( .A1(n2981), .A2(n3863), .Y(n6812) );
  AND2X4_LVT U3946 ( .A1(n2981), .A2(n3871), .Y(n6774) );
  AND2X4_LVT U3947 ( .A1(n6877), .A2(n3865), .Y(n6830) );
  AND2X4_LVT U3948 ( .A1(n6877), .A2(n3811), .Y(n6882) );
  AND2X4_LVT U3949 ( .A1(n6877), .A2(n6765), .Y(n6884) );
  AND2X4_LVT U3950 ( .A1(n2981), .A2(n3840), .Y(n6888) );
  AND2X4_LVT U3951 ( .A1(n2981), .A2(n3859), .Y(n6773) );
  AND2X4_LVT U3952 ( .A1(n6877), .A2(n6868), .Y(n6810) );
  AND2X4_LVT U3953 ( .A1(n6877), .A2(n6871), .Y(n6813) );
  NAND3X2_LVT U3954 ( .A1(n3773), .A2(n6973), .A3(n6972), .Y(n3663) );
  AND3X2_LVT U3955 ( .A1(n6973), .A2(n6948), .A3(n3709), .Y(n3666) );
  AND3X2_LVT U3956 ( .A1(n6975), .A2(n6948), .A3(n6973), .Y(n9030) );
  AND3X2_LVT U3957 ( .A1(n6973), .A2(n6972), .A3(n2983), .Y(n3768) );
  NAND4X1_LVT U3958 ( .A1(n5148), .A2(io_fpu_inst[28]), .A3(n9445), .A4(n9440), 
        .Y(n5150) );
  OR2X2_LVT U3959 ( .A1(n3079), .A2(n9520), .Y(n5129) );
  NAND3X2_LVT U3960 ( .A1(n2650), .A2(n6923), .A3(n6922), .Y(n3012) );
  AND3X2_LVT U3961 ( .A1(n6941), .A2(n6974), .A3(n6940), .Y(n9021) );
  AND3X2_LVT U3962 ( .A1(n6940), .A2(n6972), .A3(n3772), .Y(n9012) );
  AND2X4_LVT U3963 ( .A1(n2143), .A2(n6917), .Y(n6940) );
  INVX1_LVT U3964 ( .A(n9418), .Y(io_imem_req_valid) );
  IBUFFX2_LVT U3965 ( .A(n3683), .Y(n2645) );
  INVX1_LVT U3966 ( .A(n9383), .Y(n6995) );
  NOR4X1_LVT U3967 ( .A1(n1917), .A2(n9284), .A3(n9283), .A4(n9285), .Y(n1822)
         );
  AND2X1_LVT U3968 ( .A1(n6962), .A2(n6965), .Y(n6922) );
  INVX1_LVT U3969 ( .A(io_dmem_req_bits_addr[38]), .Y(n9328) );
  INVX1_LVT U3970 ( .A(n9280), .Y(n2834) );
  INVX1_LVT U3971 ( .A(n5021), .Y(n4934) );
  INVX1_LVT U3972 ( .A(n9099), .Y(n2675) );
  INVX1_LVT U3973 ( .A(n4040), .Y(n4038) );
  NOR2X1_LVT U3974 ( .A1(n9243), .A2(bpu_io_xcpt_if), .Y(n9099) );
  INVX1_LVT U3975 ( .A(n9413), .Y(n4931) );
  INVX1_LVT U3976 ( .A(n4040), .Y(n4039) );
  NOR2X0_LVT U3977 ( .A1(n6991), .A2(n2569), .Y(n2673) );
  INVX1_LVT U3978 ( .A(n6954), .Y(n4772) );
  INVX1_LVT U3979 ( .A(n6957), .Y(n4771) );
  INVX1_LVT U3980 ( .A(n4040), .Y(n9040) );
  INVX1_LVT U3981 ( .A(bpu_io_xcpt_if), .Y(n9244) );
  INVX1_LVT U3982 ( .A(n4729), .Y(n4707) );
  INVX1_LVT U3983 ( .A(n6948), .Y(n4773) );
  INVX1_LVT U3984 ( .A(n4364), .Y(n3710) );
  INVX1_LVT U3985 ( .A(n6972), .Y(n4774) );
  INVX1_LVT U3986 ( .A(n4318), .Y(n3686) );
  AND3X1_LVT U3987 ( .A1(n2570), .A2(n3077), .A3(n9446), .Y(n5396) );
  INVX1_LVT U3988 ( .A(n9288), .Y(n2569) );
  INVX1_LVT U3989 ( .A(n9109), .Y(n9073) );
  INVX1_LVT U3990 ( .A(n4691), .Y(n4692) );
  INVX1_LVT U3991 ( .A(n4401), .Y(n3645) );
  INVX1_LVT U3992 ( .A(n4445), .Y(n3660) );
  AND2X1_LVT U3993 ( .A1(n4642), .A2(ibuf_io_inst_0_bits_inst_rd[1]), .Y(n4729) );
  INVX1_LVT U3994 ( .A(n3097), .Y(n4388) );
  NOR2X0_LVT U3995 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(
        ibuf_io_inst_0_bits_inst_rd[1]), .Y(n4731) );
  INVX1_LVT U3996 ( .A(n4321), .Y(n3679) );
  AND2X1_LVT U3997 ( .A1(n4971), .A2(n2038), .Y(n6946) );
  INVX1_LVT U3998 ( .A(n5144), .Y(n5139) );
  INVX1_LVT U3999 ( .A(ibuf_io_inst_0_bits_inst_rd[0]), .Y(n4642) );
  INVX1_LVT U4000 ( .A(n9089), .Y(n9091) );
  INVX1_LVT U4001 ( .A(n5086), .Y(n9108) );
  INVX1_LVT U4002 ( .A(n3099), .Y(n4403) );
  INVX1_LVT U4003 ( .A(ibuf_io_inst_0_bits_inst_rd[4]), .Y(n4719) );
  INVX1_LVT U4004 ( .A(ibuf_io_inst_0_bits_inst_rd[1]), .Y(n4641) );
  INVX1_LVT U4005 ( .A(n3090), .Y(n4395) );
  INVX1_LVT U4006 ( .A(n4398), .Y(n3711) );
  INVX1_LVT U4007 ( .A(n4436), .Y(n3688) );
  INVX1_LVT U4008 ( .A(n9511), .Y(n9346) );
  INVX1_LVT U4009 ( .A(n3091), .Y(n4408) );
  INVX1_LVT U4010 ( .A(n9507), .Y(n9348) );
  INVX1_LVT U4011 ( .A(io_fpu_inst[20]), .Y(n9444) );
  INVX1_LVT U4012 ( .A(n3183), .Y(n4413) );
  INVX1_LVT U4013 ( .A(io_fpu_inst[9]), .Y(n3587) );
  INVX1_LVT U4014 ( .A(n4475), .Y(n3644) );
  INVX1_LVT U4015 ( .A(n2981), .Y(n3586) );
  NOR2X1_LVT U4016 ( .A1(io_fpu_inst[23]), .A2(io_fpu_inst[7]), .Y(n2616) );
  INVX1_LVT U4017 ( .A(n3092), .Y(n4356) );
  INVX1_LVT U4018 ( .A(ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4662) );
  INVX1_LVT U4019 ( .A(n4858), .Y(n4634) );
  INVX1_LVT U4020 ( .A(n3094), .Y(n4380) );
  INVX1_LVT U4021 ( .A(n3093), .Y(n4361) );
  INVX1_LVT U4022 ( .A(n9485), .Y(n9342) );
  INVX1_LVT U4023 ( .A(ibuf_io_inst_0_bits_inst_rs1[0]), .Y(n4747) );
  INVX1_LVT U4024 ( .A(n3096), .Y(n4390) );
  INVX0_LVT U4025 ( .A(ibuf_io_inst_0_bits_inst_rs1[1]), .Y(n2790) );
  INVX1_LVT U4026 ( .A(n4442), .Y(n3659) );
  INVX1_LVT U4027 ( .A(n9499), .Y(n9344) );
  INVX1_LVT U4028 ( .A(n9484), .Y(n9340) );
  INVX1_LVT U4029 ( .A(n9495), .Y(n9338) );
  INVX1_LVT U4030 ( .A(ibuf_io_inst_0_bits_replay), .Y(n9433) );
  INVX1_LVT U4031 ( .A(n4416), .Y(n3687) );
  INVX1_LVT U4032 ( .A(n5456), .Y(n4905) );
  INVX1_LVT U4033 ( .A(n5451), .Y(n4894) );
  INVX1_LVT U4034 ( .A(n3083), .Y(n3861) );
  NOR2X0_LVT U4035 ( .A1(n5436), .A2(n5435), .Y(n6837) );
  INVX1_LVT U4036 ( .A(n3083), .Y(n3862) );
  INVX1_LVT U4037 ( .A(n3095), .Y(n4378) );
  INVX1_LVT U4038 ( .A(n9425), .Y(n1281) );
  INVX1_LVT U4039 ( .A(n3098), .Y(n4421) );
  INVX1_LVT U4040 ( .A(n9503), .Y(n9336) );
  INVX1_LVT U4041 ( .A(n5454), .Y(n4873) );
  INVX1_LVT U4042 ( .A(n5449), .Y(n4874) );
  INVX1_LVT U4043 ( .A(n5450), .Y(n5438) );
  AND2X1_LVT U4044 ( .A1(n4890), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5451) );
  OR2X1_LVT U4045 ( .A1(n5434), .A2(n2878), .Y(n5447) );
  INVX1_LVT U4046 ( .A(n5452), .Y(n4906) );
  INVX1_LVT U4047 ( .A(n4890), .Y(n4898) );
  AND2X1_LVT U4048 ( .A1(n4889), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5450) );
  AND2X1_LVT U4049 ( .A1(n4900), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5449) );
  INVX1_LVT U4050 ( .A(n4889), .Y(n4899) );
  INVX1_LVT U4051 ( .A(n4860), .Y(n4633) );
  INVX0_LVT U4052 ( .A(ibuf_io_inst_0_bits_rvc), .Y(n4497) );
  INVX0_LVT U4053 ( .A(n9332), .Y(n9378) );
  INVX1_LVT U4054 ( .A(n3185), .Y(n2572) );
  INVX1_LVT U4055 ( .A(ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n4815) );
  OR2X1_LVT U4056 ( .A1(n9399), .A2(n9398), .Y(n9402) );
  INVX1_LVT U4057 ( .A(n5358), .Y(n5304) );
  AND2X1_LVT U4058 ( .A1(n5358), .A2(n5302), .Y(n3185) );
  AOI21X1_LVT U4059 ( .A1(n9256), .A2(n9255), .A3(n9254), .Y(n9276) );
  INVX1_LVT U4060 ( .A(n5254), .Y(n5256) );
  INVX1_LVT U4061 ( .A(io_fpu_fromint_data[62]), .Y(n9307) );
  INVX1_LVT U4062 ( .A(io_fpu_fromint_data[63]), .Y(n9308) );
  INVX1_LVT U4063 ( .A(io_fpu_fromint_data[61]), .Y(n9309) );
  INVX1_LVT U4064 ( .A(io_fpu_fromint_data[59]), .Y(n9310) );
  INVX1_LVT U4065 ( .A(io_fpu_fromint_data[60]), .Y(n9303) );
  INVX1_LVT U4066 ( .A(io_fpu_fromint_data[58]), .Y(n9304) );
  INVX1_LVT U4067 ( .A(io_fpu_fromint_data[56]), .Y(n9305) );
  INVX1_LVT U4068 ( .A(io_fpu_fromint_data[57]), .Y(n9306) );
  AND3X1_LVT U4069 ( .A1(n9392), .A2(n2574), .A3(n2061), .Y(n9405) );
  INVX1_LVT U4070 ( .A(n9397), .Y(n9399) );
  INVX1_LVT U4071 ( .A(n9386), .Y(n9387) );
  INVX1_LVT U4072 ( .A(n9403), .Y(n9400) );
  AND3X1_LVT U4073 ( .A1(n5314), .A2(n3046), .A3(n2575), .Y(n5307) );
  AND3X1_LVT U4074 ( .A1(n3046), .A2(n5351), .A3(n2575), .Y(n5357) );
  AND2X1_LVT U4075 ( .A1(n9120), .A2(ex_reg_rs_bypass_1), .Y(n9165) );
  AND2X1_LVT U4076 ( .A1(n9201), .A2(ex_ctrl_sel_alu2[1]), .Y(n9227) );
  NOR2X1_LVT U4077 ( .A1(n9201), .A2(n9200), .Y(n9222) );
  INVX1_LVT U4078 ( .A(wb_cause[0]), .Y(n9256) );
  INVX1_LVT U4079 ( .A(n5408), .Y(n5406) );
  INVX1_LVT U4080 ( .A(n5051), .Y(n5052) );
  INVX1_LVT U4081 ( .A(n5084), .Y(n5082) );
  INVX1_LVT U4082 ( .A(n5009), .Y(n4866) );
  INVX1_LVT U4083 ( .A(ibuf_io_inst_0_bits_raw[27]), .Y(n4781) );
  INVX1_LVT U4084 ( .A(n5301), .Y(n4944) );
  INVX0_LVT U4085 ( .A(n9179), .Y(n9201) );
  INVX1_LVT U4086 ( .A(n9172), .Y(n9174) );
  INVX1_LVT U4087 ( .A(n9178), .Y(n9180) );
  AND2X1_LVT U4088 ( .A1(n7017), .A2(n7019), .Y(n9064) );
  INVX1_LVT U4089 ( .A(n5326), .Y(n5327) );
  INVX1_LVT U4090 ( .A(n5412), .Y(n5414) );
  INVX1_LVT U4091 ( .A(n5303), .Y(n5392) );
  INVX1_LVT U4092 ( .A(n5306), .Y(n5427) );
  INVX1_LVT U4093 ( .A(n5313), .Y(n2575) );
  INVX1_LVT U4094 ( .A(n4948), .Y(n4859) );
  INVX1_LVT U4095 ( .A(csr_io_status_isa[2]), .Y(n6912) );
  INVX1_LVT U4096 ( .A(div_io_req_ready), .Y(n4917) );
  INVX1_LVT U4097 ( .A(n9330), .Y(n9331) );
  INVX1_LVT U4098 ( .A(n5413), .Y(n6860) );
  INVX0_LVT U4099 ( .A(reset), .Y(n4498) );
  INVX1_LVT U4100 ( .A(io_fpu_dec_ren2), .Y(n4837) );
  INVX1_LVT U4101 ( .A(io_fpu_sboard_clra[0]), .Y(n5182) );
  INVX0_LVT U4102 ( .A(io_dmem_s2_xcpt_pf_ld), .Y(n9246) );
  INVX1_LVT U4103 ( .A(io_fpu_dmem_resp_tag[0]), .Y(n5184) );
  INVX0_LVT U4104 ( .A(io_dmem_s2_xcpt_ma_ld), .Y(n9247) );
  INVX1_LVT U4105 ( .A(io_fpu_dec_ren3), .Y(n4838) );
  INVX0_LVT U4106 ( .A(n2030), .Y(n4943) );
  INVX1_LVT U4107 ( .A(io_fpu_sboard_clra[2]), .Y(n5257) );
  INVX1_LVT U4108 ( .A(io_fpu_dec_ren1), .Y(n4945) );
  INVX1_LVT U4109 ( .A(io_fpu_sboard_clr), .Y(n5177) );
  INVX1_LVT U4110 ( .A(io_fpu_dmem_resp_tag[2]), .Y(n5259) );
  NAND4X0_LVT U4111 ( .A1(n3023), .A2(n2655), .A3(n3705), .A4(n3022), .Y(N701)
         );
  NOR2X1_LVT U4112 ( .A1(n8835), .A2(n8836), .Y(n3732) );
  NOR2X1_LVT U4113 ( .A1(n8872), .A2(n8871), .Y(n3729) );
  NAND4X0_LVT U4114 ( .A1(n3021), .A2(n2651), .A3(n3020), .A4(n3696), .Y(N697)
         );
  NOR2X1_LVT U4115 ( .A1(n9033), .A2(n9034), .Y(n3749) );
  OA21X1_LVT U4116 ( .A1(n3476), .A2(n3994), .A3(n8553), .Y(n8556) );
  AND3X1_LVT U4117 ( .A1(n7545), .A2(n2664), .A3(n2663), .Y(n2662) );
  AO21X1_LVT U4118 ( .A1(n7350), .A2(n7351), .A3(n2645), .Y(n7352) );
  OR2X1_LVT U4119 ( .A1(n8842), .A2(n2645), .Y(n8843) );
  OR2X1_LVT U4120 ( .A1(n3371), .A2(n3988), .Y(n2661) );
  OR2X1_LVT U4121 ( .A1(n3309), .A2(n4012), .Y(n2607) );
  AOI22X1_LVT U4122 ( .A1(n_T_427[1162]), .A2(n2611), .A3(n3639), .A4(
        n_T_427[1226]), .Y(n7301) );
  AOI21X1_LVT U4123 ( .A1(n3717), .A2(n_T_427[1078]), .A3(n3776), .Y(n8740) );
  AOI21X1_LVT U4124 ( .A1(n3717), .A2(n_T_427[1064]), .A3(n3777), .Y(n8256) );
  OA21X1_LVT U4125 ( .A1(n2081), .A2(n3306), .A3(n8975), .Y(n8978) );
  OA21X1_LVT U4126 ( .A1(n4008), .A2(n3336), .A3(n8113), .Y(n8116) );
  OR2X1_LVT U4127 ( .A1(n3341), .A2(n4011), .Y(n2608) );
  OR2X1_LVT U4128 ( .A1(n8319), .A2(n2154), .Y(n8320) );
  OA21X1_LVT U4129 ( .A1(n3664), .A2(n3298), .A3(n7970), .Y(n7973) );
  OA21X1_LVT U4130 ( .A1(n2081), .A2(n3342), .A3(n8362), .Y(n8365) );
  OA21X1_LVT U4131 ( .A1(n4009), .A2(n3354), .A3(n8595), .Y(n8598) );
  OR2X1_LVT U4132 ( .A1(n9088), .A2(n1431), .Y(n9233) );
  NAND4X0_LVT U4133 ( .A1(n2677), .A2(n9231), .A3(io_fpu_inst[30]), .A4(n9230), 
        .Y(n9232) );
  OR2X1_LVT U4134 ( .A1(n9077), .A2(n1431), .Y(n9228) );
  INVX0_LVT U4135 ( .A(n2984), .Y(n4011) );
  NBUFFX2_LVT U4136 ( .A(n3658), .Y(n2897) );
  XOR2X1_LVT U4137 ( .A1(n9377), .A2(ibuf_io_pc[39]), .Y(n4574) );
  AO21X1_LVT U4138 ( .A1(n9439), .A2(n2539), .A3(n3075), .Y(n6936) );
  XOR2X1_LVT U4139 ( .A1(n9508), .A2(ibuf_io_pc[36]), .Y(n4565) );
  XOR2X1_LVT U4140 ( .A1(n9498), .A2(ibuf_io_pc[38]), .Y(n4521) );
  XOR2X1_LVT U4141 ( .A1(n9505), .A2(ibuf_io_pc[32]), .Y(n4593) );
  NOR2X1_LVT U4142 ( .A1(n5845), .A2(n5844), .Y(n5855) );
  NOR2X1_LVT U4143 ( .A1(n5566), .A2(n5565), .Y(n5576) );
  NOR2X1_LVT U4144 ( .A1(n5935), .A2(n5934), .Y(n5945) );
  XOR2X1_LVT U4145 ( .A1(n9493), .A2(ibuf_io_pc[33]), .Y(n4583) );
  NOR2X1_LVT U4146 ( .A1(n5658), .A2(n5657), .Y(n5668) );
  XOR2X1_LVT U4147 ( .A1(n9374), .A2(ibuf_io_pc[35]), .Y(n4576) );
  XOR2X1_LVT U4148 ( .A1(n9502), .A2(ibuf_io_pc[31]), .Y(n4563) );
  XOR2X1_LVT U4149 ( .A1(n9373), .A2(n4557), .Y(n4558) );
  NOR2X1_LVT U4150 ( .A1(n6330), .A2(n6329), .Y(n6340) );
  NOR2X1_LVT U4151 ( .A1(n6495), .A2(n6494), .Y(n6505) );
  NOR2X1_LVT U4152 ( .A1(n6172), .A2(n6171), .Y(n6182) );
  NOR2X1_LVT U4153 ( .A1(n5979), .A2(n5978), .Y(n5989) );
  NOR2X1_LVT U4154 ( .A1(n5515), .A2(n5514), .Y(n5525) );
  OA22X1_LVT U4155 ( .A1(n3559), .A2(n3882), .A3(n3877), .A4(n6549), .Y(n6552)
         );
  OA22X1_LVT U4156 ( .A1(n3539), .A2(n3880), .A3(n3879), .A4(n5751), .Y(n5753)
         );
  OA22X1_LVT U4157 ( .A1(n3542), .A2(n3881), .A3(n3879), .A4(n5813), .Y(n5814)
         );
  AOI22X1_LVT U4158 ( .A1(n3834), .A2(n_T_427[405]), .A3(n_T_427[469]), .A4(
        n2824), .Y(n2845) );
  OA22X1_LVT U4159 ( .A1(n3564), .A2(n3882), .A3(n1993), .A4(n6674), .Y(n6677)
         );
  OA22X1_LVT U4160 ( .A1(n3533), .A2(n3880), .A3(n3879), .A4(n5595), .Y(n5598)
         );
  OA22X1_LVT U4161 ( .A1(n3560), .A2(n3882), .A3(n1993), .A4(n6577), .Y(n6580)
         );
  AOI22X1_LVT U4162 ( .A1(n5776), .A2(n1992), .A3(n_T_427[1897]), .A4(n3884), 
        .Y(n2756) );
  OA22X1_LVT U4163 ( .A1(n3540), .A2(n3880), .A3(n3879), .A4(n5784), .Y(n5788)
         );
  OA22X1_LVT U4164 ( .A1(n3558), .A2(n3882), .A3(n1993), .A4(n6500), .Y(n6502)
         );
  AOI22X1_LVT U4165 ( .A1(n2856), .A2(n_T_427[342]), .A3(n_T_427[86]), .A4(
        n2872), .Y(n2683) );
  AOI22X1_LVT U4166 ( .A1(n2872), .A2(n_T_427[71]), .A3(n_T_427[902]), .A4(
        n3897), .Y(n2729) );
  OA22X1_LVT U4167 ( .A1(n3562), .A2(n3882), .A3(n3877), .A4(n6622), .Y(n6625)
         );
  OA22X1_LVT U4168 ( .A1(n3277), .A2(n3882), .A3(n1993), .A4(n6525), .Y(n6527)
         );
  AOI22X1_LVT U4169 ( .A1(n5495), .A2(n6877), .A3(n_T_427[1884]), .A4(n3884), 
        .Y(n2789) );
  OA22X1_LVT U4170 ( .A1(n3536), .A2(n3880), .A3(n3879), .A4(n5663), .Y(n5666)
         );
  AOI22X1_LVT U4171 ( .A1(n5545), .A2(n6877), .A3(n_T_427[1886]), .A4(n3884), 
        .Y(n2785) );
  AND4X1_LVT U4172 ( .A1(n9096), .A2(n9095), .A3(n9109), .A4(n9094), .Y(n2676)
         );
  NOR2X1_LVT U4173 ( .A1(n6280), .A2(n6279), .Y(n6290) );
  OA22X1_LVT U4174 ( .A1(n3538), .A2(n3880), .A3(n3879), .A4(n5712), .Y(n5714)
         );
  OA22X1_LVT U4175 ( .A1(n3531), .A2(n3880), .A3(n3879), .A4(n5520), .Y(n5523)
         );
  AOI22X1_LVT U4176 ( .A1(n6258), .A2(n6877), .A3(n_T_427[1919]), .A4(n3884), 
        .Y(n2760) );
  AOI22X1_LVT U4177 ( .A1(n3798), .A2(n_T_427[1762]), .A3(n_T_427[1823]), .A4(
        n3830), .Y(n2746) );
  AOI22X1_LVT U4178 ( .A1(n6772), .A2(n1992), .A3(n_T_427[1939]), .A4(n3884), 
        .Y(n2823) );
  AOI22X1_LVT U4179 ( .A1(n3901), .A2(n_T_427[1070]), .A3(n_T_427[239]), .A4(
        n6773), .Y(n2736) );
  AOI22X1_LVT U4180 ( .A1(n3835), .A2(n_T_427[431]), .A3(n_T_427[750]), .A4(
        n3905), .Y(n2737) );
  AOI22X1_LVT U4181 ( .A1(n3902), .A2(n_T_427[1081]), .A3(n_T_427[250]), .A4(
        n3807), .Y(n2732) );
  OR3X1_LVT U4182 ( .A1(n5133), .A2(n9109), .A3(n9096), .Y(n1612) );
  AOI22X1_LVT U4183 ( .A1(n2864), .A2(n_T_427[429]), .A3(n_T_427[109]), .A4(
        n3833), .Y(n2709) );
  OA22X1_LVT U4184 ( .A1(n3555), .A2(n3882), .A3(n3877), .A4(n6402), .Y(n6405)
         );
  OA22X1_LVT U4185 ( .A1(n3532), .A2(n3880), .A3(n3879), .A4(n5571), .Y(n5574)
         );
  OA22X1_LVT U4186 ( .A1(n3537), .A2(n3880), .A3(n3879), .A4(n5694), .Y(n5697)
         );
  AOI22X1_LVT U4187 ( .A1(n6376), .A2(n1992), .A3(n_T_427[1924]), .A4(n3884), 
        .Y(n2764) );
  NOR2X1_LVT U4188 ( .A1(n5689), .A2(n5688), .Y(n5699) );
  AOI22X1_LVT U4189 ( .A1(n2867), .A2(n_T_427[1756]), .A3(n_T_427[1818]), .A4(
        n3829), .Y(n2766) );
  XOR2X1_LVT U4190 ( .A1(n9486), .A2(ibuf_io_pc[20]), .Y(n4585) );
  XOR2X1_LVT U4191 ( .A1(n9501), .A2(ibuf_io_pc[22]), .Y(n4584) );
  OA22X1_LVT U4192 ( .A1(n3535), .A2(n3880), .A3(n3879), .A4(n5639), .Y(n5642)
         );
  XOR2X1_LVT U4193 ( .A1(n9364), .A2(ibuf_io_pc[24]), .Y(n4590) );
  XOR2X1_LVT U4194 ( .A1(n9368), .A2(ibuf_io_pc[28]), .Y(n4589) );
  XOR2X1_LVT U4195 ( .A1(n9488), .A2(ibuf_io_pc[23]), .Y(n4560) );
  XOR2X1_LVT U4196 ( .A1(n9483), .A2(ibuf_io_pc[26]), .Y(n4520) );
  XOR2X1_LVT U4197 ( .A1(n9489), .A2(ibuf_io_pc[27]), .Y(n4561) );
  OA22X1_LVT U4198 ( .A1(n3534), .A2(n3880), .A3(n3879), .A4(n5615), .Y(n5618)
         );
  AOI22X1_LVT U4199 ( .A1(n3893), .A2(n_T_427[1579]), .A3(n_T_427[1643]), .A4(
        n3887), .Y(n2763) );
  AOI22X1_LVT U4200 ( .A1(n3945), .A2(n_T_427[1194]), .A3(n_T_427[1258]), .A4(
        n3940), .Y(n2694) );
  XOR2X1_LVT U4201 ( .A1(n9506), .A2(ibuf_io_pc[14]), .Y(n4555) );
  AOI22X1_LVT U4202 ( .A1(n3945), .A2(n_T_427[1198]), .A3(n_T_427[1262]), .A4(
        n3939), .Y(n2734) );
  XOR2X1_LVT U4203 ( .A1(n9491), .A2(ibuf_io_pc[12]), .Y(n4554) );
  AOI22X1_LVT U4204 ( .A1(n3955), .A2(n_T_427[1130]), .A3(n_T_427[1002]), .A4(
        n3950), .Y(n2695) );
  AOI22X1_LVT U4205 ( .A1(n3955), .A2(n_T_427[1134]), .A3(n_T_427[1006]), .A4(
        n3949), .Y(n2735) );
  OR2X1_LVT U4206 ( .A1(n2644), .A2(n5143), .Y(n2643) );
  NOR2X1_LVT U4207 ( .A1(csr_io_interrupt), .A2(bpu_io_debug_if), .Y(n5167) );
  XOR2X1_LVT U4208 ( .A1(n9496), .A2(ibuf_io_pc[18]), .Y(n4556) );
  AOI22X1_LVT U4209 ( .A1(n3955), .A2(n_T_427[1132]), .A3(n_T_427[1004]), .A4(
        n3949), .Y(n2707) );
  AOI22X1_LVT U4210 ( .A1(n3945), .A2(n_T_427[1196]), .A3(n_T_427[1260]), .A4(
        n3939), .Y(n2706) );
  AOI22X1_LVT U4211 ( .A1(n3901), .A2(n_T_427[1059]), .A3(n_T_427[931]), .A4(
        n3895), .Y(n2740) );
  AOI22X1_LVT U4212 ( .A1(n2824), .A2(n_T_427[484]), .A3(n_T_427[739]), .A4(
        n3904), .Y(n2741) );
  AOI22X1_LVT U4213 ( .A1(n3955), .A2(n_T_427[1135]), .A3(n_T_427[1007]), .A4(
        n3950), .Y(n2723) );
  INVX1_LVT U4214 ( .A(n4040), .Y(n4037) );
  AOI22X1_LVT U4215 ( .A1(n3945), .A2(n_T_427[1191]), .A3(n_T_427[1255]), .A4(
        n3939), .Y(n2718) );
  AOI22X1_LVT U4216 ( .A1(n3955), .A2(n_T_427[1127]), .A3(n_T_427[999]), .A4(
        n3949), .Y(n2719) );
  NAND3X0_LVT U4217 ( .A1(n2565), .A2(n3078), .A3(n9436), .Y(n5146) );
  AOI22X1_LVT U4218 ( .A1(n2861), .A2(n_T_427[810]), .A3(n_T_427[746]), .A4(
        n3904), .Y(n2697) );
  XOR2X1_LVT U4219 ( .A1(n9497), .A2(ibuf_io_pc[25]), .Y(n4582) );
  AOI22X1_LVT U4220 ( .A1(n2866), .A2(n_T_427[1760]), .A3(n_T_427[1821]), .A4(
        n3829), .Y(n2751) );
  XOR2X1_LVT U4221 ( .A1(n9356), .A2(n4518), .Y(n4519) );
  AOI22X1_LVT U4222 ( .A1(n3945), .A2(n_T_427[1200]), .A3(n_T_427[1264]), .A4(
        n3939), .Y(n2698) );
  AOI22X1_LVT U4223 ( .A1(n3955), .A2(n_T_427[1136]), .A3(n_T_427[1008]), .A4(
        n3949), .Y(n2699) );
  AOI22X1_LVT U4224 ( .A1(n3890), .A2(n_T_427[1537]), .A3(n_T_427[1601]), .A4(
        n3885), .Y(n2788) );
  AOI22X1_LVT U4225 ( .A1(n3893), .A2(n_T_427[1581]), .A3(n_T_427[1645]), .A4(
        n3888), .Y(n2780) );
  AOI22X1_LVT U4226 ( .A1(n6428), .A2(n1992), .A3(n_T_427[1926]), .A4(n3884), 
        .Y(n2781) );
  AOI22X1_LVT U4227 ( .A1(n3924), .A2(n_T_427[1498]), .A3(n_T_427[1370]), .A4(
        n3918), .Y(n2773) );
  AOI22X1_LVT U4228 ( .A1(n3901), .A2(n_T_427[1068]), .A3(n_T_427[940]), .A4(
        n2831), .Y(n2708) );
  AOI22X1_LVT U4229 ( .A1(n3945), .A2(n_T_427[1199]), .A3(n_T_427[1263]), .A4(
        n3940), .Y(n2722) );
  AOI22X1_LVT U4230 ( .A1(n2861), .A2(n_T_427[788]), .A3(n_T_427[341]), .A4(
        n2857), .Y(n2843) );
  INVX1_LVT U4231 ( .A(n6949), .Y(n8982) );
  AOI22X1_LVT U4232 ( .A1(n2824), .A2(n_T_427[470]), .A3(n_T_427[917]), .A4(
        n2831), .Y(n2682) );
  NOR2X1_LVT U4233 ( .A1(n6956), .A2(n6947), .Y(n9038) );
  AOI22X1_LVT U4234 ( .A1(n3923), .A2(n_T_427[1491]), .A3(n_T_427[1363]), .A4(
        n3918), .Y(n2802) );
  AOI22X1_LVT U4235 ( .A1(n3956), .A2(n_T_427[1144]), .A3(n_T_427[1016]), .A4(
        n3951), .Y(n2743) );
  AOI22X1_LVT U4236 ( .A1(n3946), .A2(n_T_427[1208]), .A3(n_T_427[1272]), .A4(
        n3941), .Y(n2742) );
  AOI22X1_LVT U4237 ( .A1(n3927), .A2(n_T_427[1280]), .A3(n_T_427[1216]), .A4(
        n3937), .Y(n2855) );
  AOI22X1_LVT U4238 ( .A1(n2860), .A2(n_T_427[825]), .A3(n_T_427[761]), .A4(
        n3905), .Y(n2733) );
  AOI22X1_LVT U4239 ( .A1(n3956), .A2(n_T_427[1145]), .A3(n_T_427[1017]), .A4(
        n3951), .Y(n2731) );
  AOI22X1_LVT U4240 ( .A1(n3946), .A2(n_T_427[1209]), .A3(n_T_427[1273]), .A4(
        n3941), .Y(n2730) );
  INVX0_LVT U4241 ( .A(n6991), .Y(n6993) );
  AOI22X1_LVT U4242 ( .A1(n3923), .A2(n_T_427[1481]), .A3(n_T_427[1353]), .A4(
        n3917), .Y(n2794) );
  NOR2X1_LVT U4243 ( .A1(n1531), .A2(io_fpu_inst[14]), .Y(n5116) );
  AOI22X1_LVT U4244 ( .A1(n3924), .A2(n_T_427[1489]), .A3(n_T_427[1361]), .A4(
        n3918), .Y(n2818) );
  NAND2X0_LVT U4245 ( .A1(n5067), .A2(n3578), .Y(n2635) );
  AOI22X1_LVT U4246 ( .A1(n1919), .A2(n_T_427[337]), .A3(n_T_427[529]), .A4(
        n3819), .Y(n2679) );
  AOI22X1_LVT U4247 ( .A1(n3823), .A2(n_T_427[848]), .A3(n_T_427[657]), .A4(
        n3821), .Y(n2681) );
  AOI22X1_LVT U4248 ( .A1(n3894), .A2(n_T_427[1595]), .A3(n_T_427[1659]), .A4(
        n3888), .Y(n2822) );
  AOI22X1_LVT U4249 ( .A1(n3829), .A2(n_T_427[1846]), .A3(n_T_427[1723]), .A4(
        n3824), .Y(n2821) );
  AOI22X1_LVT U4250 ( .A1(n3907), .A2(n_T_427[786]), .A3(n_T_427[467]), .A4(
        n3910), .Y(n2839) );
  AOI22X1_LVT U4251 ( .A1(n3924), .A2(n_T_427[1480]), .A3(n_T_427[1352]), .A4(
        n3917), .Y(n2814) );
  AOI22X1_LVT U4252 ( .A1(n3955), .A2(n_T_427[1138]), .A3(n_T_427[1010]), .A4(
        n3950), .Y(n2711) );
  AOI22X1_LVT U4253 ( .A1(n3945), .A2(n_T_427[1202]), .A3(n_T_427[1266]), .A4(
        n3940), .Y(n2710) );
  AOI22X1_LVT U4254 ( .A1(n3956), .A2(n_T_427[1141]), .A3(n_T_427[1013]), .A4(
        n3951), .Y(n2691) );
  AOI22X1_LVT U4255 ( .A1(n3946), .A2(n_T_427[1205]), .A3(n_T_427[1269]), .A4(
        n3941), .Y(n2690) );
  AOI22X1_LVT U4256 ( .A1(n3818), .A2(n_T_427[512]), .A3(n_T_427[576]), .A4(
        n3916), .Y(n2880) );
  AOI22X1_LVT U4257 ( .A1(n3956), .A2(n_T_427[1143]), .A3(n_T_427[1015]), .A4(
        n3950), .Y(n2703) );
  AOI22X1_LVT U4258 ( .A1(n3946), .A2(n_T_427[1207]), .A3(n_T_427[1271]), .A4(
        n3940), .Y(n2702) );
  NAND3X0_LVT U4259 ( .A1(n3566), .A2(n5136), .A3(n3567), .Y(n2644) );
  INVX1_LVT U4260 ( .A(n3097), .Y(n4387) );
  NAND3X0_LVT U4261 ( .A1(n9076), .A2(n9075), .A3(io_fpu_inst[30]), .Y(n9077)
         );
  AND2X1_LVT U4262 ( .A1(n4749), .A2(n2038), .Y(n6954) );
  OR2X1_LVT U4263 ( .A1(n2825), .A2(n6955), .Y(n6949) );
  NOR2X1_LVT U4264 ( .A1(n6956), .A2(n6955), .Y(n3182) );
  INVX1_LVT U4265 ( .A(n6955), .Y(n6926) );
  INVX1_LVT U4266 ( .A(n4730), .Y(n4708) );
  INVX0_LVT U4267 ( .A(n4847), .Y(n4618) );
  NAND4X0_LVT U4268 ( .A1(n4690), .A2(n3046), .A3(n4689), .A4(n4688), .Y(n4695) );
  XOR2X1_LVT U4269 ( .A1(n9487), .A2(ibuf_io_pc[17]), .Y(n4551) );
  NAND4X0_LVT U4270 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n2625), .Y(n5036) );
  XOR2X1_LVT U4271 ( .A1(n9507), .A2(ibuf_io_pc[9]), .Y(n4547) );
  XOR2X1_LVT U4272 ( .A1(n9511), .A2(ibuf_io_pc[8]), .Y(n4549) );
  AND2X1_LVT U4273 ( .A1(n4641), .A2(ibuf_io_inst_0_bits_inst_rd[0]), .Y(n4732) );
  INVX1_LVT U4274 ( .A(n3195), .Y(n4358) );
  OR2X1_LVT U4275 ( .A1(io_fpu_inst[6]), .A2(io_fpu_inst[2]), .Y(n9109) );
  AOI21X1_LVT U4276 ( .A1(n3843), .A2(csr_io_rw_rdata[25]), .A3(n5953), .Y(
        n3097) );
  NAND4X0_LVT U4277 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n3046), .Y(n5003) );
  INVX1_LVT U4278 ( .A(n3195), .Y(n4357) );
  XOR2X1_LVT U4279 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n3202), .Y(n4946) );
  NAND4X0_LVT U4280 ( .A1(n9445), .A2(n1867), .A3(io_fpu_inst[6]), .A4(n3577), 
        .Y(n9081) );
  AO21X1_LVT U4281 ( .A1(io_fpu_inst[5]), .A2(io_fpu_inst[14]), .A3(
        io_fpu_inst[2]), .Y(n9094) );
  AND3X1_LVT U4282 ( .A1(n3044), .A2(io_fpu_inst[14]), .A3(n9435), .Y(n5107)
         );
  NAND2X0_LVT U4283 ( .A1(n5100), .A2(n2552), .Y(n2636) );
  NAND2X0_LVT U4284 ( .A1(n5446), .A2(n5452), .Y(n3082) );
  INVX1_LVT U4285 ( .A(n3189), .Y(n4345) );
  AO21X1_LVT U4286 ( .A1(io_fpu_inst[14]), .A2(n9105), .A3(n9435), .Y(n5097)
         );
  INVX1_LVT U4287 ( .A(n3192), .Y(n4342) );
  OR2X1_LVT U4288 ( .A1(io_fpu_inst[21]), .A2(io_fpu_inst[20]), .Y(n5394) );
  INVX1_LVT U4289 ( .A(n3193), .Y(n4354) );
  XOR2X1_LVT U4290 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n588), .Y(n5031)
         );
  XOR2X1_LVT U4291 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n590), .Y(n5033)
         );
  NOR4X0_LVT U4292 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n2877), .A3(
        ibuf_io_inst_0_bits_inst_rs1[0]), .A4(ibuf_io_inst_0_bits_inst_rs1[2]), 
        .Y(n3588) );
  NOR2X1_LVT U4293 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(
        ibuf_io_inst_0_bits_inst_rd[4]), .Y(n4700) );
  INVX1_LVT U4294 ( .A(n3192), .Y(n4340) );
  INVX1_LVT U4295 ( .A(ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4733) );
  INVX1_LVT U4296 ( .A(n3190), .Y(n4329) );
  INVX1_LVT U4297 ( .A(n3092), .Y(n4355) );
  INVX1_LVT U4298 ( .A(n3193), .Y(n4352) );
  AND2X1_LVT U4299 ( .A1(n5434), .A2(n6238), .Y(n6877) );
  INVX1_LVT U4300 ( .A(n3189), .Y(n4343) );
  INVX1_LVT U4301 ( .A(n3099), .Y(n4402) );
  INVX1_LVT U4302 ( .A(n3091), .Y(n4407) );
  IBUFFX2_LVT U4303 ( .A(n6238), .Y(n6898) );
  INVX1_LVT U4304 ( .A(n3090), .Y(n4394) );
  INVX1_LVT U4305 ( .A(n3193), .Y(n4353) );
  INVX1_LVT U4306 ( .A(n3183), .Y(n4412) );
  XOR2X1_LVT U4307 ( .A1(n9485), .A2(ibuf_io_pc[6]), .Y(n4546) );
  INVX1_LVT U4308 ( .A(n3192), .Y(n4341) );
  INVX1_LVT U4309 ( .A(n3190), .Y(n4328) );
  INVX1_LVT U4310 ( .A(n3189), .Y(n4344) );
  INVX1_LVT U4311 ( .A(n3186), .Y(n4350) );
  INVX1_LVT U4312 ( .A(n3196), .Y(n4323) );
  AOI21X1_LVT U4313 ( .A1(n3842), .A2(csr_io_rw_rdata[13]), .A3(n5707), .Y(
        n3092) );
  INVX1_LVT U4314 ( .A(n3187), .Y(n4326) );
  INVX1_LVT U4315 ( .A(n3197), .Y(n4332) );
  INVX1_LVT U4316 ( .A(n3194), .Y(n4335) );
  INVX1_LVT U4317 ( .A(n3191), .Y(n4338) );
  NOR2X1_LVT U4318 ( .A1(csr_io_interrupt), .A2(ibuf_io_inst_0_bits_replay), 
        .Y(n9385) );
  AOI21X1_LVT U4319 ( .A1(n3842), .A2(csr_io_rw_rdata[12]), .A3(n5683), .Y(
        n3193) );
  AOI21X1_LVT U4320 ( .A1(n3843), .A2(csr_io_rw_rdata[28]), .A3(n6014), .Y(
        n3090) );
  INVX1_LVT U4321 ( .A(n3187), .Y(n4327) );
  INVX1_LVT U4322 ( .A(n3196), .Y(n4322) );
  INVX1_LVT U4323 ( .A(ibuf_io_inst_0_bits_inst_rs1[4]), .Y(n6963) );
  INVX1_LVT U4324 ( .A(n3197), .Y(n4331) );
  INVX1_LVT U4325 ( .A(n3094), .Y(n4379) );
  INVX1_LVT U4326 ( .A(n3191), .Y(n4339) );
  INVX1_LVT U4327 ( .A(n3096), .Y(n4389) );
  AOI21X1_LVT U4328 ( .A1(n3843), .A2(csr_io_rw_rdata[31]), .A3(n6083), .Y(
        n3099) );
  AOI21X1_LVT U4329 ( .A1(n3842), .A2(csr_io_rw_rdata[9]), .A3(n5628), .Y(
        n3189) );
  INVX1_LVT U4330 ( .A(n3196), .Y(n4324) );
  AOI21X1_LVT U4331 ( .A1(n3842), .A2(csr_io_rw_rdata[8]), .A3(n5604), .Y(
        n3192) );
  INVX1_LVT U4332 ( .A(n3197), .Y(n4333) );
  INVX1_LVT U4333 ( .A(n3187), .Y(n4325) );
  INVX1_LVT U4334 ( .A(n3194), .Y(n4334) );
  INVX1_LVT U4335 ( .A(csr_io_interrupt), .Y(n9448) );
  INVX1_LVT U4336 ( .A(n3191), .Y(n4337) );
  INVX1_LVT U4337 ( .A(n3194), .Y(n4336) );
  INVX1_LVT U4338 ( .A(n3093), .Y(n4360) );
  INVX1_LVT U4339 ( .A(n3186), .Y(n4349) );
  OR2X1_LVT U4340 ( .A1(csr_io_status_isa[3]), .A2(n3583), .Y(n3570) );
  AOI21X1_LVT U4341 ( .A1(n3841), .A2(csr_io_rw_rdata[7]), .A3(n5584), .Y(
        n3191) );
  AOI21X1_LVT U4342 ( .A1(n3841), .A2(csr_io_rw_rdata[3]), .A3(n5505), .Y(
        n3187) );
  INVX1_LVT U4343 ( .A(n3188), .Y(n4348) );
  INVX0_LVT U4344 ( .A(n9525), .Y(n5067) );
  AOI21X1_LVT U4345 ( .A1(n3841), .A2(csr_io_rw_rdata[6]), .A3(n5560), .Y(
        n3194) );
  IBUFFX2_LVT U4346 ( .A(n5075), .Y(n2571) );
  INVX1_LVT U4347 ( .A(n3083), .Y(n3863) );
  NBUFFX2_LVT U4348 ( .A(n6794), .Y(n3811) );
  AOI21X1_LVT U4349 ( .A1(n3843), .A2(csr_io_rw_rdata[15]), .A3(n5746), .Y(
        n3093) );
  AOI21X1_LVT U4350 ( .A1(n3843), .A2(csr_io_rw_rdata[26]), .A3(n5973), .Y(
        n3096) );
  INVX1_LVT U4351 ( .A(n3188), .Y(n4346) );
  INVX1_LVT U4352 ( .A(n3188), .Y(n4347) );
  AOI21X1_LVT U4353 ( .A1(n3841), .A2(csr_io_rw_rdata[2]), .A3(n5486), .Y(
        n3196) );
  AOI21X1_LVT U4354 ( .A1(n3841), .A2(csr_io_rw_rdata[5]), .A3(n5536), .Y(
        n3197) );
  INVX1_LVT U4355 ( .A(n3095), .Y(n4377) );
  INVX1_LVT U4356 ( .A(n3098), .Y(n4420) );
  AND2X1_LVT U4357 ( .A1(n4890), .A2(n4816), .Y(n5456) );
  INVX1_LVT U4358 ( .A(n5435), .Y(n5455) );
  AOI21X1_LVT U4359 ( .A1(n3844), .A2(csr_io_rw_rdata[21]), .A3(n5863), .Y(
        n3095) );
  AOI21X1_LVT U4360 ( .A1(n3842), .A2(csr_io_rw_rdata[10]), .A3(n5652), .Y(
        n3188) );
  NBUFFX2_LVT U4361 ( .A(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(n3781) );
  OR2X1_LVT U4362 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n4814), .Y(n5435) );
  AOI21X1_LVT U4363 ( .A1(n3842), .A2(csr_io_rw_rdata[38]), .A3(n6232), .Y(
        n3098) );
  AND2X1_LVT U4364 ( .A1(n4889), .A2(n4816), .Y(n5452) );
  AND2X1_LVT U4365 ( .A1(n4900), .A2(n4816), .Y(n5454) );
  NOR2X0_LVT U4366 ( .A1(wb_reg_flush_pipe), .A2(n9332), .Y(
        io_imem_req_bits_speculative) );
  NOR2X1_LVT U4367 ( .A1(n_T_726[1]), .A2(n_T_726[0]), .Y(n9430) );
  NAND4X0_LVT U4368 ( .A1(n4870), .A2(n4869), .A3(n3046), .A4(n4868), .Y(n4888) );
  AND2X1_LVT U4369 ( .A1(n9387), .A2(n9388), .Y(n9394) );
  NOR2X1_LVT U4370 ( .A1(n9400), .A2(n9402), .Y(n9401) );
  NOR2X1_LVT U4371 ( .A1(n9331), .A2(n4065), .Y(n9414) );
  NOR2X0_LVT U4372 ( .A1(n9403), .A2(n9402), .Y(n9410) );
  OR2X1_LVT U4373 ( .A1(n5359), .A2(n5358), .Y(n5393) );
  NOR2X1_LVT U4374 ( .A1(n5362), .A2(n5358), .Y(n5378) );
  OR2X1_LVT U4375 ( .A1(n5327), .A2(n5358), .Y(n5334) );
  NOR2X1_LVT U4376 ( .A1(n5381), .A2(n5358), .Y(n5366) );
  NOR2X1_LVT U4377 ( .A1(n5365), .A2(n5358), .Y(n5383) );
  NAND2X0_LVT U4378 ( .A1(n9380), .A2(n4498), .Y(n5358) );
  AO21X1_LVT U4379 ( .A1(n9103), .A2(io_fpu_fromint_data[43]), .A3(n9102), .Y(
        alu_io_in1[43]) );
  AO21X1_LVT U4380 ( .A1(n9103), .A2(io_fpu_fromint_data[41]), .A3(n9102), .Y(
        alu_io_in1[41]) );
  NOR2X1_LVT U4381 ( .A1(n5365), .A2(n5254), .Y(n5275) );
  AO22X1_LVT U4382 ( .A1(n_T_698[27]), .A2(n9101), .A3(io_fpu_fromint_data[27]), .A4(n9103), .Y(alu_io_in1[27]) );
  AO22X1_LVT U4383 ( .A1(n_T_698[28]), .A2(n9101), .A3(io_fpu_fromint_data[28]), .A4(n9103), .Y(alu_io_in1[28]) );
  AO21X1_LVT U4384 ( .A1(n9103), .A2(io_fpu_fromint_data[55]), .A3(n9102), .Y(
        alu_io_in1[55]) );
  NOR2X1_LVT U4385 ( .A1(n5381), .A2(n5254), .Y(n5265) );
  AO22X1_LVT U4386 ( .A1(n_T_698[25]), .A2(n9101), .A3(io_fpu_fromint_data[25]), .A4(n9103), .Y(alu_io_in1[25]) );
  AO21X1_LVT U4387 ( .A1(n9103), .A2(io_fpu_fromint_data[51]), .A3(n9102), .Y(
        alu_io_in1[51]) );
  AO22X1_LVT U4388 ( .A1(n4054), .A2(n_T_698[26]), .A3(io_fpu_fromint_data[26]), .A4(n9103), .Y(alu_io_in1[26]) );
  AO21X1_LVT U4389 ( .A1(n9103), .A2(io_fpu_fromint_data[49]), .A3(n9102), .Y(
        alu_io_in1[49]) );
  AO22X1_LVT U4390 ( .A1(n9101), .A2(n_T_698[11]), .A3(io_fpu_fromint_data[11]), .A4(n9103), .Y(alu_io_in1[11]) );
  AO21X1_LVT U4391 ( .A1(n9103), .A2(io_fpu_fromint_data[39]), .A3(n9102), .Y(
        alu_io_in1[39]) );
  AO22X1_LVT U4392 ( .A1(n_T_698[8]), .A2(n4054), .A3(io_fpu_fromint_data[8]), 
        .A4(n9103), .Y(alu_io_in1[8]) );
  AO22X1_LVT U4393 ( .A1(n_T_698[9]), .A2(n4054), .A3(io_fpu_fromint_data[9]), 
        .A4(n9103), .Y(alu_io_in1[9]) );
  AO22X1_LVT U4394 ( .A1(n9101), .A2(n_T_698[5]), .A3(io_fpu_fromint_data[5]), 
        .A4(n9103), .Y(alu_io_in1[5]) );
  NOR2X1_LVT U4395 ( .A1(n5362), .A2(n5254), .Y(n5285) );
  AO21X1_LVT U4396 ( .A1(n9103), .A2(io_fpu_fromint_data[63]), .A3(n9102), .Y(
        alu_io_in1[63]) );
  AND3X1_LVT U4397 ( .A1(n9400), .A2(n9398), .A3(n9397), .Y(n9396) );
  AO22X1_LVT U4398 ( .A1(n_T_698[31]), .A2(n9101), .A3(io_fpu_fromint_data[31]), .A4(n9103), .Y(alu_io_in1[31]) );
  NOR2X1_LVT U4399 ( .A1(n5392), .A2(n5254), .Y(n5248) );
  OR2X1_LVT U4400 ( .A1(n7905), .A2(n7904), .Y(io_fpu_fromint_data[31]) );
  NAND2X0_LVT U4401 ( .A1(csr_io_retire), .A2(n5176), .Y(n5254) );
  INVX0_LVT U4402 ( .A(ibuf_io_inst_0_bits_raw[1]), .Y(n3646) );
  IBUFFX2_LVT U4403 ( .A(n3042), .Y(n2573) );
  NOR3X1_LVT U4404 ( .A1(n3203), .A2(n9330), .A3(csr_io_exception), .Y(
        csr_io_retire) );
  IBUFFX2_LVT U4405 ( .A(n3040), .Y(n2574) );
  MUX21X1_LVT U4406 ( .A1(wb_reg_cause[1]), .A2(n9251), .S0(n576), .Y(
        wb_cause[1]) );
  NOR2X1_LVT U4407 ( .A1(n_T_728[1]), .A2(n_T_728[0]), .Y(n9118) );
  OR2X1_LVT U4408 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(
        ibuf_io_inst_0_bits_raw[28]), .Y(n4804) );
  NOR2X0_LVT U4409 ( .A1(n6860), .A2(n5415), .Y(n6861) );
  NOR2X1_LVT U4410 ( .A1(mem_ctrl_jalr), .A2(mem_reg_sfence), .Y(n4591) );
  NOR2X1_LVT U4411 ( .A1(n5426), .A2(n5428), .Y(n5314) );
  INVX0_LVT U4412 ( .A(ibuf_io_inst_0_bits_raw[28]), .Y(n4782) );
  AND3X1_LVT U4413 ( .A1(n7019), .A2(n3101), .A3(n3255), .Y(n9066) );
  OR2X1_LVT U4414 ( .A1(io_dmem_s2_nack), .A2(wb_reg_replay), .Y(n9330) );
  NBUFFX2_LVT U4415 ( .A(net34480), .Y(n4285) );
  INVX1_LVT U4416 ( .A(n3784), .Y(n3785) );
  INVX1_LVT U4417 ( .A(io_fpu_dmem_resp_tag[4]), .Y(n5228) );
  AND2X1_LVT U4418 ( .A1(io_dmem_resp_valid), .A2(io_dmem_resp_bits_has_data), 
        .Y(n2626) );
  INVX1_LVT U4419 ( .A(io_fpu_dmem_resp_tag[1]), .Y(n5185) );
  INVX0_LVT U4420 ( .A(io_dmem_perf_grant), .Y(n5065) );
  INVX1_LVT U4421 ( .A(io_fpu_dmem_resp_tag[3]), .Y(n5249) );
  INVX0_LVT U4422 ( .A(io_fpu_fcsr_rdy), .Y(n4918) );
  INVX0_LVT U4423 ( .A(io_dmem_req_ready), .Y(n5064) );
  OR2X1_LVT U4424 ( .A1(io_fpu_dmem_resp_tag[3]), .A2(io_fpu_dmem_resp_tag[4]), 
        .Y(n5192) );
  NAND3X0_LVT U4425 ( .A1(n8870), .A2(n8868), .A3(n2577), .Y(n8871) );
  OA21X1_LVT U4426 ( .A1(n4011), .A2(n3368), .A3(n8869), .Y(n2577) );
  OA21X1_LVT U4427 ( .A1(n4012), .A2(n3356), .A3(n8618), .Y(n2578) );
  OA21X1_LVT U4428 ( .A1(n4012), .A2(n3347), .A3(n8451), .Y(n2579) );
  OA21X1_LVT U4429 ( .A1(n4013), .A2(n3350), .A3(n8515), .Y(n2580) );
  NAND2X0_LVT U4430 ( .A1(n_T_427[490]), .A2(n3614), .Y(n8264) );
  IBUFFX2_LVT U4431 ( .A(n3663), .Y(n2611) );
  NAND4X0_LVT U4432 ( .A1(n3662), .A2(n3780), .A3(n2910), .A4(n2581), .Y(N735)
         );
  NOR3X0_LVT U4433 ( .A1(n2582), .A2(n8888), .A3(n8889), .Y(n3730) );
  AND3X1_LVT U4434 ( .A1(n7355), .A2(n7356), .A3(n2583), .Y(n2958) );
  OA21X1_LVT U4435 ( .A1(n3439), .A2(n4008), .A3(n7357), .Y(n2583) );
  AND3X1_LVT U4436 ( .A1(n2935), .A2(n7271), .A3(n7272), .Y(n2584) );
  AND3X1_LVT U4437 ( .A1(n7937), .A2(n7936), .A3(n7938), .Y(n2585) );
  NAND2X0_LVT U4438 ( .A1(n_T_427[486]), .A2(n3614), .Y(n8125) );
  IBUFFX2_LVT U4439 ( .A(n2984), .Y(n4012) );
  OR2X1_LVT U4440 ( .A1(n3427), .A2(n3653), .Y(n2586) );
  NAND2X0_LVT U4441 ( .A1(n2611), .A2(n_T_427[1155]), .Y(n2587) );
  NAND2X0_LVT U4442 ( .A1(n_T_427[1219]), .A2(n3638), .Y(n2588) );
  OR3X2_LVT U4443 ( .A1(io_fpu_inst[4]), .A2(n3593), .A3(n9528), .Y(n9113) );
  NAND2X0_LVT U4444 ( .A1(n_T_427[303]), .A2(n3790), .Y(n2589) );
  AND2X1_LVT U4445 ( .A1(n8218), .A2(n8219), .Y(n2602) );
  NAND2X0_LVT U4446 ( .A1(n_T_427[498]), .A2(n3614), .Y(n8550) );
  AND4X1_LVT U4447 ( .A1(n8099), .A2(n8100), .A3(n8098), .A4(n8097), .Y(n2950)
         );
  NAND2X0_LVT U4448 ( .A1(n_T_427[480]), .A2(n3614), .Y(n7923) );
  AND2X1_LVT U4449 ( .A1(n8349), .A2(n8348), .Y(n2590) );
  AND4X1_LVT U4450 ( .A1(n7958), .A2(n7957), .A3(n7956), .A4(n7955), .Y(n2963)
         );
  NAND2X0_LVT U4451 ( .A1(n_T_427[312]), .A2(n3790), .Y(n2591) );
  NAND2X0_LVT U4452 ( .A1(n_T_427[1431]), .A2(n3629), .Y(n2592) );
  AND3X1_LVT U4453 ( .A1(n2594), .A2(n8961), .A3(n3050), .Y(n2987) );
  AND2X1_LVT U4454 ( .A1(n8962), .A2(n8960), .Y(n2594) );
  AOI21X1_LVT U4455 ( .A1(n9429), .A2(n9107), .A3(n9445), .Y(n2657) );
  NAND2X0_LVT U4456 ( .A1(n2596), .A2(n2646), .Y(n4513) );
  NOR4X1_LVT U4457 ( .A1(n4501), .A2(n9437), .A3(n2606), .A4(n4500), .Y(n2596)
         );
  OR2X1_LVT U4458 ( .A1(n3191), .A2(n2089), .Y(n2597) );
  AND2X1_LVT U4459 ( .A1(n3960), .A2(n8105), .Y(n9052) );
  AND2X1_LVT U4460 ( .A1(n8631), .A2(n2598), .Y(n2617) );
  DELLN1X2_LVT U4461 ( .A(n9052), .Y(n3614) );
  AND2X1_LVT U4462 ( .A1(n3678), .A2(n2599), .Y(n2910) );
  AND3X1_LVT U4463 ( .A1(n8739), .A2(n8738), .A3(n8740), .Y(n2599) );
  NOR3X0_LVT U4464 ( .A1(n2601), .A2(n8222), .A3(n8221), .Y(n3746) );
  OA21X1_LVT U4465 ( .A1(n4011), .A2(n3344), .A3(n8383), .Y(n2604) );
  OA21X1_LVT U4466 ( .A1(n4012), .A2(n3300), .A3(n8418), .Y(n2605) );
  OR2X1_LVT U4467 ( .A1(io_fpu_inst[7]), .A2(io_fpu_inst[26]), .Y(n2606) );
  NAND4X0_LVT U4468 ( .A1(n9032), .A2(n9027), .A3(n9031), .A4(n2607), .Y(n9033) );
  NAND4X0_LVT U4469 ( .A1(n8204), .A2(n8202), .A3(n8203), .A4(n2609), .Y(n8205) );
  OR2X1_LVT U4470 ( .A1(n3338), .A2(n4013), .Y(n2609) );
  NAND2X0_LVT U4471 ( .A1(n_T_427[1457]), .A2(n3627), .Y(n8562) );
  OA21X1_LVT U4472 ( .A1(n3752), .A2(n3282), .A3(n7426), .Y(n2610) );
  IBUFFX2_LVT U4473 ( .A(n3768), .Y(n3664) );
  IBUFFX2_LVT U4474 ( .A(n3768), .Y(n4008) );
  IBUFFX2_LVT U4475 ( .A(n3768), .Y(n4009) );
  AOI22X1_LVT U4476 ( .A1(n4330), .A2(n2982), .A3(n2966), .A4(n_T_427[1411]), 
        .Y(n7105) );
  OR2X1_LVT U4477 ( .A1(n3459), .A2(n3658), .Y(n2612) );
  NAND4X0_LVT U4478 ( .A1(n8074), .A2(n8076), .A3(n8075), .A4(n2613), .Y(n8077) );
  OR2X1_LVT U4479 ( .A1(n3455), .A2(n3658), .Y(n2613) );
  OR2X1_LVT U4480 ( .A1(n3403), .A2(n3658), .Y(n2614) );
  AND2X1_LVT U4481 ( .A1(n9446), .A2(n2616), .Y(n2615) );
  NBUFFX2_LVT U4482 ( .A(io_fpu_inst[12]), .Y(n2618) );
  IBUFFX2_LVT U4483 ( .A(n3683), .Y(n3631) );
  IBUFFX2_LVT U4484 ( .A(n9527), .Y(n3783) );
  NAND2X0_LVT U4485 ( .A1(n9438), .A2(n5144), .Y(n2620) );
  AND2X1_LVT U4486 ( .A1(n2544), .A2(n6906), .Y(n2621) );
  OA21X1_LVT U4487 ( .A1(n4010), .A2(n3428), .A3(n7190), .Y(n2622) );
  OA21X1_LVT U4488 ( .A1(n2643), .A2(n2639), .A3(n2640), .Y(n2624) );
  XNOR2X1_LVT U4489 ( .A1(n3782), .A2(n589), .Y(n2625) );
  OR2X2_LVT U4490 ( .A1(n5036), .A2(n5013), .Y(n6992) );
  INVX1_LVT U4491 ( .A(n6931), .Y(n6947) );
  NAND2X0_LVT U4492 ( .A1(n6956), .A2(n6931), .Y(n4040) );
  AND2X1_LVT U4493 ( .A1(n2038), .A2(n4970), .Y(n6931) );
  MUX21X1_LVT U4494 ( .A1(n3043), .A2(n5313), .S0(n9381), .Y(n3042) );
  MUX21X1_LVT U4495 ( .A1(io_fpu_dmem_resp_tag[2]), .A2(
        div_io_resp_bits_tag[2]), .S0(n5403), .Y(n5313) );
  NAND2X0_LVT U4496 ( .A1(n2153), .A2(n4685), .Y(n5413) );
  AND3X1_LVT U4497 ( .A1(n5124), .A2(n2628), .A3(n2627), .Y(n6939) );
  NAND2X0_LVT U4498 ( .A1(n5122), .A2(n3049), .Y(n6916) );
  OA21X1_LVT U4499 ( .A1(n3072), .A2(n5123), .A3(
        csr_io_decode_0_system_illegal), .Y(n6915) );
  OR2X1_LVT U4500 ( .A1(csr_io_status_isa[2]), .A2(n4497), .Y(n2628) );
  AND2X1_LVT U4501 ( .A1(n5106), .A2(n5105), .Y(n2630) );
  AND2X1_LVT U4502 ( .A1(n2631), .A2(n2658), .Y(n2633) );
  OA22X1_LVT U4503 ( .A1(n2635), .A2(n2636), .A3(n5098), .A4(n2634), .Y(n2631)
         );
  AND4X1_LVT U4504 ( .A1(n5104), .A2(n5103), .A3(n9445), .A4(n2632), .Y(n2637)
         );
  NAND2X0_LVT U4505 ( .A1(n3635), .A2(n_T_427[1271]), .Y(n2638) );
  OA21X1_LVT U4506 ( .A1(n5135), .A2(n5134), .A3(n5140), .Y(n2640) );
  OR2X1_LVT U4507 ( .A1(n3656), .A2(n8521), .Y(n8522) );
  AO21X1_LVT U4508 ( .A1(n7321), .A2(n7322), .A3(n2154), .Y(n7323) );
  AO21X1_LVT U4509 ( .A1(n7377), .A2(n7378), .A3(n3632), .Y(n7379) );
  AO21X1_LVT U4510 ( .A1(n7779), .A2(n7780), .A3(n2645), .Y(n7781) );
  AO21X1_LVT U4511 ( .A1(n7811), .A2(n7812), .A3(n2154), .Y(n7813) );
  AO21X1_LVT U4512 ( .A1(n7747), .A2(n7748), .A3(n2155), .Y(n7749) );
  AO21X1_LVT U4513 ( .A1(n7871), .A2(n7872), .A3(n3656), .Y(n7873) );
  AND2X1_LVT U4514 ( .A1(n4503), .A2(n4502), .Y(n2646) );
  AND2X1_LVT U4515 ( .A1(n3577), .A2(n9439), .Y(n2647) );
  AND2X1_LVT U4516 ( .A1(n3077), .A2(n3577), .Y(n2648) );
  AND2X1_LVT U4517 ( .A1(io_fpu_inst[3]), .A2(n5163), .Y(n9428) );
  NAND2X0_LVT U4518 ( .A1(n3577), .A2(n5067), .Y(n9095) );
  AND3X1_LVT U4519 ( .A1(n6966), .A2(n6917), .A3(n6946), .Y(n2650) );
  AND4X1_LVT U4520 ( .A1(n2652), .A2(n7455), .A3(n2653), .A4(n3697), .Y(n2651)
         );
  AND2X1_LVT U4521 ( .A1(n7456), .A2(n7457), .Y(n2652) );
  OR2X1_LVT U4522 ( .A1(n3139), .A2(n3987), .Y(n2653) );
  AND4X1_LVT U4523 ( .A1(n3706), .A2(n2656), .A3(n7576), .A4(n2654), .Y(n2655)
         );
  AND2X1_LVT U4524 ( .A1(n7577), .A2(n7578), .Y(n2654) );
  AND2X1_LVT U4525 ( .A1(n5102), .A2(n9104), .Y(n9429) );
  NAND2X0_LVT U4526 ( .A1(n3991), .A2(n_T_427[1903]), .Y(n2660) );
  AND3X1_LVT U4527 ( .A1(n3701), .A2(n3702), .A3(n2659), .Y(n3028) );
  AND4X1_LVT U4528 ( .A1(n7609), .A2(n7608), .A3(n2661), .A4(n2660), .Y(n2659)
         );
  NAND2X0_LVT U4529 ( .A1(n2882), .A2(n_T_427[1901]), .Y(n2663) );
  AND4X1_LVT U4530 ( .A1(n3703), .A2(n3704), .A3(n7546), .A4(n2662), .Y(n3017)
         );
  NAND3X0_LVT U4531 ( .A1(n3006), .A2(n2666), .A3(n2665), .Y(N710) );
  AND4X1_LVT U4532 ( .A1(n3005), .A2(n3065), .A3(n3064), .A4(n2668), .Y(n2665)
         );
  AND2X1_LVT U4533 ( .A1(n2667), .A2(n7860), .Y(n2666) );
  AND2X1_LVT U4534 ( .A1(n7861), .A2(n7862), .Y(n2667) );
  AND2X1_LVT U4535 ( .A1(n3180), .A2(n3580), .Y(n2670) );
  AND2X1_LVT U4536 ( .A1(n3765), .A2(n2561), .Y(n6941) );
  AND2X1_LVT U4537 ( .A1(n2143), .A2(n2672), .Y(n2671) );
  AND2X1_LVT U4538 ( .A1(n6917), .A2(n6954), .Y(n2672) );
  XOR2X1_LVT U4539 ( .A1(n2876), .A2(n591), .Y(n5037) );
  NAND2X0_LVT U4540 ( .A1(n2673), .A2(n2538), .Y(n5094) );
  AOI21X1_LVT U4541 ( .A1(n2676), .A2(n9116), .A3(n2675), .Y(N279) );
  INVX1_LVT U4542 ( .A(n4732), .Y(n4675) );
  AND2X1_LVT U4543 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(
        ibuf_io_inst_0_bits_inst_rd[0]), .Y(n4730) );
  AOI21X1_LVT U4544 ( .A1(n9281), .A2(n3048), .A3(n9280), .Y(n9283) );
  AOI22X1_LVT U4545 ( .A1(n3903), .A2(n_T_427[721]), .A3(n_T_427[17]), .A4(
        n3914), .Y(n2680) );
  AOI22X1_LVT U4546 ( .A1(n3908), .A2(n_T_427[149]), .A3(n_T_427[277]), .A4(
        n2828), .Y(n2844) );
  AOI22X1_LVT U4547 ( .A1(n2864), .A2(n_T_427[401]), .A3(n_T_427[1040]), .A4(
        n3898), .Y(n2678) );
  AND4X1_LVT U4548 ( .A1(n2678), .A2(n2679), .A3(n2680), .A4(n2681), .Y(n5794)
         );
  AND2X1_LVT U4549 ( .A1(n2682), .A2(n2683), .Y(n5895) );
  AOI22X1_LVT U4550 ( .A1(n3902), .A2(n_T_427[1080]), .A3(n_T_427[249]), .A4(
        n3808), .Y(n2744) );
  OA22X1_LVT U4551 ( .A1(n3371), .A2(n3080), .A3(n3881), .A4(n2684), .Y(n2775)
         );
  AND2X1_LVT U4552 ( .A1(n2685), .A2(n2686), .Y(n6132) );
  AOI22X1_LVT U4553 ( .A1(n3833), .A2(n_T_427[97]), .A3(n_T_427[225]), .A4(
        n3806), .Y(n2685) );
  AOI22X1_LVT U4554 ( .A1(n2831), .A2(n_T_427[928]), .A3(n_T_427[161]), .A4(
        n2862), .Y(n2686) );
  AOI22X1_LVT U4555 ( .A1(n3900), .A2(n_T_427[1055]), .A3(n_T_427[224]), .A4(
        n3808), .Y(n2687) );
  AOI22X1_LVT U4556 ( .A1(n2870), .A2(n_T_427[608]), .A3(n_T_427[32]), .A4(
        n2879), .Y(n2688) );
  AOI22X1_LVT U4557 ( .A1(n3819), .A2(n_T_427[544]), .A3(n_T_427[863]), .A4(
        n3823), .Y(n2689) );
  AND4X1_LVT U4558 ( .A1(n2690), .A2(n2691), .A3(n2692), .A4(n2693), .Y(n6628)
         );
  AOI22X1_LVT U4559 ( .A1(n3902), .A2(n_T_427[1077]), .A3(n_T_427[949]), .A4(
        n3895), .Y(n2692) );
  AOI22X1_LVT U4560 ( .A1(n3906), .A2(n_T_427[821]), .A3(n_T_427[438]), .A4(
        n2865), .Y(n2693) );
  AND4X1_LVT U4561 ( .A1(n2694), .A2(n2695), .A3(n2696), .A4(n2697), .Y(n6362)
         );
  AOI22X1_LVT U4562 ( .A1(n3901), .A2(n_T_427[1066]), .A3(n_T_427[938]), .A4(
        n3896), .Y(n2696) );
  AND4X1_LVT U4563 ( .A1(n2698), .A2(n2699), .A3(n2700), .A4(n2701), .Y(n6506)
         );
  AOI22X1_LVT U4564 ( .A1(n3901), .A2(n_T_427[1072]), .A3(n_T_427[113]), .A4(
        n3833), .Y(n2700) );
  AOI22X1_LVT U4565 ( .A1(n3910), .A2(n_T_427[497]), .A3(n_T_427[752]), .A4(
        n2827), .Y(n2701) );
  AND4X1_LVT U4566 ( .A1(n2702), .A2(n2703), .A3(n2704), .A4(n2705), .Y(n6680)
         );
  AOI22X1_LVT U4567 ( .A1(n3902), .A2(n_T_427[1079]), .A3(n_T_427[951]), .A4(
        n3897), .Y(n2704) );
  AOI22X1_LVT U4568 ( .A1(n3835), .A2(n_T_427[440]), .A3(n_T_427[184]), .A4(
        n2863), .Y(n2705) );
  AOI22X1_LVT U4569 ( .A1(n2856), .A2(n_T_427[351]), .A3(n_T_427[95]), .A4(
        n3831), .Y(n2847) );
  AND4X1_LVT U4570 ( .A1(n2706), .A2(n2707), .A3(n2708), .A4(n2709), .Y(n6408)
         );
  AND4X1_LVT U4571 ( .A1(n2710), .A2(n2711), .A3(n2712), .A4(n2713), .Y(n6555)
         );
  AOI22X1_LVT U4572 ( .A1(n3902), .A2(n_T_427[1074]), .A3(n_T_427[243]), .A4(
        n2830), .Y(n2712) );
  AOI22X1_LVT U4573 ( .A1(n2832), .A2(n_T_427[946]), .A3(n_T_427[754]), .A4(
        n2827), .Y(n2713) );
  AND4X1_LVT U4574 ( .A1(n2714), .A2(n2715), .A3(n2716), .A4(n2717), .Y(n6224)
         );
  AOI22X1_LVT U4575 ( .A1(n3944), .A2(n_T_427[1188]), .A3(n_T_427[1252]), .A4(
        n3939), .Y(n2714) );
  AOI22X1_LVT U4576 ( .A1(n3954), .A2(n_T_427[1124]), .A3(n_T_427[996]), .A4(
        n3949), .Y(n2715) );
  AOI22X1_LVT U4577 ( .A1(n3901), .A2(n_T_427[1060]), .A3(n_T_427[229]), .A4(
        n3807), .Y(n2716) );
  AOI22X1_LVT U4578 ( .A1(n3832), .A2(n_T_427[101]), .A3(n_T_427[740]), .A4(
        n6884), .Y(n2717) );
  AND4X1_LVT U4579 ( .A1(n2718), .A2(n2719), .A3(n2720), .A4(n2721), .Y(n6291)
         );
  AOI22X1_LVT U4580 ( .A1(n3901), .A2(n_T_427[1063]), .A3(n_T_427[232]), .A4(
        n3808), .Y(n2720) );
  AOI22X1_LVT U4581 ( .A1(n3833), .A2(n_T_427[104]), .A3(n_T_427[935]), .A4(
        n3896), .Y(n2721) );
  AND4X1_LVT U4582 ( .A1(n2722), .A2(n2723), .A3(n2724), .A4(n2725), .Y(n6482)
         );
  AOI22X1_LVT U4583 ( .A1(n3901), .A2(n_T_427[1071]), .A3(n_T_427[240]), .A4(
        n3807), .Y(n2724) );
  AOI22X1_LVT U4584 ( .A1(n3834), .A2(n_T_427[432]), .A3(n_T_427[943]), .A4(
        n2832), .Y(n2725) );
  AND4X1_LVT U4585 ( .A1(n2726), .A2(n2727), .A3(n2728), .A4(n2729), .Y(n5601)
         );
  AOI22X1_LVT U4586 ( .A1(n3943), .A2(n_T_427[1158]), .A3(n_T_427[1222]), .A4(
        n3937), .Y(n2726) );
  AOI22X1_LVT U4587 ( .A1(n3953), .A2(n_T_427[1094]), .A3(n_T_427[966]), .A4(
        n3947), .Y(n2727) );
  AOI22X1_LVT U4588 ( .A1(n3899), .A2(n_T_427[1030]), .A3(n_T_427[199]), .A4(
        n3808), .Y(n2728) );
  AND4X1_LVT U4589 ( .A1(n2730), .A2(n2731), .A3(n2732), .A4(n2733), .Y(n6726)
         );
  AND4X1_LVT U4590 ( .A1(n2734), .A2(n2735), .A3(n2736), .A4(n2737), .Y(n6457)
         );
  AND4X1_LVT U4591 ( .A1(n2738), .A2(n2739), .A3(n2740), .A4(n2741), .Y(n6203)
         );
  AOI22X1_LVT U4592 ( .A1(n3944), .A2(n_T_427[1187]), .A3(n_T_427[1251]), .A4(
        n3939), .Y(n2738) );
  AOI22X1_LVT U4593 ( .A1(n3954), .A2(n_T_427[1123]), .A3(n_T_427[995]), .A4(
        n3949), .Y(n2739) );
  AND4X1_LVT U4594 ( .A1(n2742), .A2(n2743), .A3(n2744), .A4(n2745), .Y(n6701)
         );
  AOI22X1_LVT U4595 ( .A1(n3831), .A2(n_T_427[121]), .A3(n_T_427[760]), .A4(
        n3905), .Y(n2745) );
  IBUFFX2_LVT U4596 ( .A(n6878), .Y(n3884) );
  AND4X1_LVT U4597 ( .A1(n2746), .A2(n2747), .A3(n2748), .A4(n2749), .Y(n6184)
         );
  AOI22X1_LVT U4598 ( .A1(n2028), .A2(n_T_427[1876]), .A3(n3884), .A4(
        n_T_427[1915]), .Y(n2747) );
  AOI22X1_LVT U4599 ( .A1(n3827), .A2(n_T_427[1698]), .A3(n_T_427[1570]), .A4(
        n3890), .Y(n2748) );
  AOI22X1_LVT U4600 ( .A1(n3889), .A2(n_T_427[1634]), .A3(n_T_427[1506]), .A4(
        n3922), .Y(n2749) );
  AOI22X1_LVT U4601 ( .A1(n2028), .A2(n_T_427[1857]), .A3(n3884), .A4(
        n_T_427[1892]), .Y(n2750) );
  AND4X1_LVT U4602 ( .A1(n2751), .A2(n2752), .A3(n2753), .A4(n2754), .Y(n6134)
         );
  AOI22X1_LVT U4603 ( .A1(n3801), .A2(n_T_427[1874]), .A3(n3884), .A4(
        n_T_427[1913]), .Y(n2752) );
  AOI22X1_LVT U4604 ( .A1(n3827), .A2(n_T_427[1696]), .A3(n_T_427[1568]), .A4(
        n3890), .Y(n2753) );
  AOI22X1_LVT U4605 ( .A1(n3889), .A2(n_T_427[1632]), .A3(n_T_427[1504]), .A4(
        n3922), .Y(n2754) );
  AOI22X1_LVT U4606 ( .A1(n6764), .A2(n_T_427[1862]), .A3(n_T_427[1743]), .A4(
        n3798), .Y(n2755) );
  AND4X1_LVT U4607 ( .A1(n2757), .A2(n2758), .A3(n2759), .A4(n2760), .Y(n6270)
         );
  AOI22X1_LVT U4608 ( .A1(n3801), .A2(n_T_427[1878]), .A3(n_T_427[1766]), .A4(
        n2867), .Y(n2757) );
  AOI22X1_LVT U4609 ( .A1(n2765), .A2(n_T_427[1827]), .A3(n_T_427[1702]), .A4(
        n3825), .Y(n2758) );
  AOI22X1_LVT U4610 ( .A1(n3892), .A2(n_T_427[1574]), .A3(n_T_427[1638]), .A4(
        n3887), .Y(n2759) );
  AND4X1_LVT U4611 ( .A1(n2761), .A2(n2762), .A3(n2763), .A4(n2764), .Y(n6388)
         );
  AOI22X1_LVT U4612 ( .A1(n6764), .A2(n_T_427[1879]), .A3(n_T_427[1771]), .A4(
        n2866), .Y(n2761) );
  AOI22X1_LVT U4613 ( .A1(n3828), .A2(n_T_427[1832]), .A3(n_T_427[1707]), .A4(
        n3825), .Y(n2762) );
  AND4X1_LVT U4614 ( .A1(n2766), .A2(n2767), .A3(n2768), .A4(n2769), .Y(n6047)
         );
  AOI22X1_LVT U4615 ( .A1(n3801), .A2(n_T_427[1872]), .A3(n3884), .A4(
        n_T_427[1910]), .Y(n2767) );
  AOI22X1_LVT U4616 ( .A1(n3826), .A2(n_T_427[1692]), .A3(n_T_427[1564]), .A4(
        n3890), .Y(n2768) );
  AOI22X1_LVT U4617 ( .A1(n3889), .A2(n_T_427[1628]), .A3(n_T_427[1500]), .A4(
        n3922), .Y(n2769) );
  AND4X1_LVT U4618 ( .A1(n2770), .A2(n2771), .A3(n2772), .A4(n2773), .Y(n6011)
         );
  AOI22X1_LVT U4619 ( .A1(n6764), .A2(n_T_427[1870]), .A3(n_T_427[1754]), .A4(
        n2867), .Y(n2770) );
  AOI22X1_LVT U4620 ( .A1(n3830), .A2(n_T_427[1816]), .A3(n_T_427[1690]), .A4(
        n3826), .Y(n2771) );
  AOI22X1_LVT U4621 ( .A1(n3892), .A2(n_T_427[1562]), .A3(n_T_427[1626]), .A4(
        n3886), .Y(n2772) );
  AND4X1_LVT U4622 ( .A1(n2774), .A2(n2775), .A3(n2776), .A4(n2777), .Y(n5897)
         );
  AOI22X1_LVT U4623 ( .A1(n3798), .A2(n_T_427[1749]), .A3(n_T_427[1811]), .A4(
        n2765), .Y(n2774) );
  AOI22X1_LVT U4624 ( .A1(n3827), .A2(n_T_427[1685]), .A3(n_T_427[1557]), .A4(
        n3890), .Y(n2776) );
  AOI22X1_LVT U4625 ( .A1(n3889), .A2(n_T_427[1621]), .A3(n_T_427[1493]), .A4(
        n3922), .Y(n2777) );
  AND4X1_LVT U4626 ( .A1(n2778), .A2(n2779), .A3(n2780), .A4(n2781), .Y(n6435)
         );
  AOI22X1_LVT U4627 ( .A1(n3802), .A2(n_T_427[1880]), .A3(n_T_427[1773]), .A4(
        n2867), .Y(n2778) );
  AOI22X1_LVT U4628 ( .A1(n3828), .A2(n_T_427[1834]), .A3(n_T_427[1709]), .A4(
        n3825), .Y(n2779) );
  AND4X1_LVT U4629 ( .A1(n2782), .A2(n2783), .A3(n2784), .A4(n2785), .Y(n5552)
         );
  AOI22X1_LVT U4630 ( .A1(n6764), .A2(n_T_427[1851]), .A3(n_T_427[1732]), .A4(
        n2866), .Y(n2782) );
  AOI22X1_LVT U4631 ( .A1(n3828), .A2(n_T_427[1795]), .A3(n_T_427[1668]), .A4(
        n3826), .Y(n2783) );
  AOI22X1_LVT U4632 ( .A1(n3892), .A2(n_T_427[1540]), .A3(n_T_427[1604]), .A4(
        n3885), .Y(n2784) );
  AND4X1_LVT U4633 ( .A1(n2786), .A2(n2787), .A3(n2788), .A4(n2789), .Y(n5501)
         );
  AOI22X1_LVT U4634 ( .A1(n3802), .A2(n_T_427[1848]), .A3(n_T_427[1729]), .A4(
        n2867), .Y(n2786) );
  AOI22X1_LVT U4635 ( .A1(n3829), .A2(n_T_427[1792]), .A3(n_T_427[1665]), .A4(
        n3826), .Y(n2787) );
  AND4X1_LVT U4636 ( .A1(n2791), .A2(n2792), .A3(n2793), .A4(n2794), .Y(n5670)
         );
  AOI22X1_LVT U4637 ( .A1(n3801), .A2(n_T_427[1856]), .A3(n_T_427[1737]), .A4(
        n2868), .Y(n2791) );
  AOI22X1_LVT U4638 ( .A1(n3830), .A2(n_T_427[1800]), .A3(n_T_427[1673]), .A4(
        n3826), .Y(n2792) );
  AOI22X1_LVT U4639 ( .A1(n3891), .A2(n_T_427[1545]), .A3(n_T_427[1609]), .A4(
        n3885), .Y(n2793) );
  AND4X1_LVT U4640 ( .A1(n2795), .A2(n2796), .A3(n2797), .A4(n2798), .Y(n5622)
         );
  AOI22X1_LVT U4641 ( .A1(n3802), .A2(n_T_427[1854]), .A3(n_T_427[1735]), .A4(
        n2867), .Y(n2795) );
  AOI22X1_LVT U4642 ( .A1(n2765), .A2(n_T_427[1798]), .A3(n_T_427[1671]), .A4(
        n3826), .Y(n2796) );
  AOI22X1_LVT U4643 ( .A1(n3891), .A2(n_T_427[1543]), .A3(n_T_427[1607]), .A4(
        n3885), .Y(n2797) );
  AOI22X1_LVT U4644 ( .A1(n3923), .A2(n_T_427[1479]), .A3(n_T_427[1351]), .A4(
        n3917), .Y(n2798) );
  AND4X1_LVT U4645 ( .A1(n2799), .A2(n2800), .A3(n2801), .A4(n2802), .Y(n5857)
         );
  AOI22X1_LVT U4646 ( .A1(n3802), .A2(n_T_427[1865]), .A3(n_T_427[1747]), .A4(
        n2866), .Y(n2799) );
  AOI22X1_LVT U4647 ( .A1(n3892), .A2(n_T_427[1555]), .A3(n_T_427[1619]), .A4(
        n3886), .Y(n2801) );
  AND4X1_LVT U4648 ( .A1(n2803), .A2(n2804), .A3(n2805), .A4(n2806), .Y(n5701)
         );
  AOI22X1_LVT U4649 ( .A1(n3801), .A2(n_T_427[1858]), .A3(n_T_427[1739]), .A4(
        n2868), .Y(n2803) );
  AOI22X1_LVT U4650 ( .A1(n3828), .A2(n_T_427[1802]), .A3(n_T_427[1675]), .A4(
        n3826), .Y(n2804) );
  AOI22X1_LVT U4651 ( .A1(n3891), .A2(n_T_427[1547]), .A3(n_T_427[1611]), .A4(
        n3885), .Y(n2805) );
  AOI22X1_LVT U4652 ( .A1(n3923), .A2(n_T_427[1483]), .A3(n_T_427[1355]), .A4(
        n3917), .Y(n2806) );
  AND4X1_LVT U4653 ( .A1(n2807), .A2(n2808), .A3(n2809), .A4(n2810), .Y(n5578)
         );
  AOI22X1_LVT U4654 ( .A1(n3802), .A2(n_T_427[1852]), .A3(n_T_427[1733]), .A4(
        n2868), .Y(n2807) );
  AOI22X1_LVT U4655 ( .A1(n3829), .A2(n_T_427[1796]), .A3(n_T_427[1669]), .A4(
        n3826), .Y(n2808) );
  AOI22X1_LVT U4656 ( .A1(n3891), .A2(n_T_427[1541]), .A3(n_T_427[1605]), .A4(
        n3885), .Y(n2809) );
  AOI22X1_LVT U4657 ( .A1(n3923), .A2(n_T_427[1477]), .A3(n_T_427[1349]), .A4(
        n3917), .Y(n2810) );
  AND4X1_LVT U4658 ( .A1(n2811), .A2(n2812), .A3(n2813), .A4(n2814), .Y(n5646)
         );
  AOI22X1_LVT U4659 ( .A1(n3801), .A2(n_T_427[1855]), .A3(n_T_427[1736]), .A4(
        n2866), .Y(n2811) );
  AOI22X1_LVT U4660 ( .A1(n3830), .A2(n_T_427[1799]), .A3(n_T_427[1672]), .A4(
        n3826), .Y(n2812) );
  AOI22X1_LVT U4661 ( .A1(n3891), .A2(n_T_427[1544]), .A3(n_T_427[1608]), .A4(
        n3885), .Y(n2813) );
  AND4X1_LVT U4662 ( .A1(n2815), .A2(n2816), .A3(n2817), .A4(n2818), .Y(n5820)
         );
  AOI22X1_LVT U4663 ( .A1(n6764), .A2(n_T_427[1863]), .A3(n_T_427[1745]), .A4(
        n2867), .Y(n2815) );
  AOI22X1_LVT U4664 ( .A1(n3830), .A2(n_T_427[1807]), .A3(n_T_427[1681]), .A4(
        n3825), .Y(n2816) );
  AOI22X1_LVT U4665 ( .A1(n3892), .A2(n_T_427[1553]), .A3(n_T_427[1617]), .A4(
        n3886), .Y(n2817) );
  AOI22X1_LVT U4666 ( .A1(n2028), .A2(n_T_427[1860]), .A3(n_T_427[1741]), .A4(
        n3798), .Y(n2819) );
  AND4X1_LVT U4667 ( .A1(n2820), .A2(n2821), .A3(n2822), .A4(n2823), .Y(n6786)
         );
  AOI22X1_LVT U4668 ( .A1(n6764), .A2(n_T_427[1881]), .A3(n_T_427[1787]), .A4(
        n3798), .Y(n2820) );
  NBUFFX2_LVT U4669 ( .A(n6887), .Y(n2824) );
  NBUFFX2_LVT U4670 ( .A(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(n2825) );
  NBUFFX2_LVT U4671 ( .A(n6888), .Y(n2826) );
  NBUFFX2_LVT U4672 ( .A(n6884), .Y(n2827) );
  NBUFFX2_LVT U4673 ( .A(n6774), .Y(n2828) );
  NBUFFX2_LVT U4674 ( .A(n6812), .Y(n2829) );
  NBUFFX2_LVT U4675 ( .A(n6773), .Y(n2830) );
  IBUFFX2_LVT U4676 ( .A(n3781), .Y(n5436) );
  INVX1_LVT U4677 ( .A(n5906), .Y(n6796) );
  NBUFFX2_LVT U4678 ( .A(n6882), .Y(n2831) );
  NBUFFX2_LVT U4679 ( .A(n6882), .Y(n2832) );
  AOI22X1_LVT U4680 ( .A1(n3895), .A2(n_T_427[926]), .A3(n_T_427[735]), .A4(
        n3904), .Y(n2846) );
  AOI22X1_LVT U4681 ( .A1(n3834), .A2(n_T_427[385]), .A3(n_T_427[65]), .A4(
        n3832), .Y(n2852) );
  NBUFFX2_LVT U4682 ( .A(n6813), .Y(n2833) );
  NAND2X0_LVT U4683 ( .A1(n2834), .A2(n2835), .Y(n5060) );
  AND3X1_LVT U4684 ( .A1(n5008), .A2(n5007), .A3(n5006), .Y(n2835) );
  NBUFFX2_LVT U4685 ( .A(n9041), .Y(n2836) );
  NBUFFX2_LVT U4686 ( .A(n9041), .Y(n2837) );
  XOR2X1_LVT U4687 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n3202), .Y(
        n4846) );
  AOI22X1_LVT U4688 ( .A1(n3835), .A2(n_T_427[403]), .A3(n_T_427[83]), .A4(
        n2871), .Y(n2838) );
  AOI22X1_LVT U4689 ( .A1(n3817), .A2(n_T_427[339]), .A3(n6774), .A4(
        n_T_427[275]), .Y(n2840) );
  AND2X1_LVT U4690 ( .A1(n5833), .A2(n5832), .Y(n2841) );
  AND4X1_LVT U4691 ( .A1(n2842), .A2(n2843), .A3(n2844), .A4(n2845), .Y(n5877)
         );
  AND2X1_LVT U4692 ( .A1(n5870), .A2(n5869), .Y(n2842) );
  AND4X1_LVT U4693 ( .A1(n2846), .A2(n2847), .A3(n2848), .A4(n2849), .Y(n6097)
         );
  AOI22X1_LVT U4694 ( .A1(n3823), .A2(n_T_427[862]), .A3(n_T_427[159]), .A4(
        n2863), .Y(n2848) );
  AND2X1_LVT U4695 ( .A1(n6089), .A2(n6090), .Y(n2849) );
  NBUFFX2_LVT U4696 ( .A(n6811), .Y(n2850) );
  NBUFFX2_LVT U4697 ( .A(n6811), .Y(n2851) );
  INVX1_LVT U4698 ( .A(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(n4816) );
  AOI22X1_LVT U4699 ( .A1(n3943), .A2(n_T_427[1152]), .A3(n_T_427[1024]), .A4(
        n3898), .Y(n2853) );
  AOI22X1_LVT U4700 ( .A1(n3953), .A2(n_T_427[1088]), .A3(n_T_427[960]), .A4(
        n3947), .Y(n2854) );
  IBUFFX2_LVT U4701 ( .A(n6423), .Y(n6865) );
  NBUFFX2_LVT U4702 ( .A(n6810), .Y(n2856) );
  NBUFFX2_LVT U4703 ( .A(n6810), .Y(n2857) );
  NBUFFX2_LVT U4704 ( .A(n8932), .Y(n2858) );
  NBUFFX2_LVT U4705 ( .A(n6885), .Y(n2860) );
  NBUFFX2_LVT U4706 ( .A(n6885), .Y(n2861) );
  NBUFFX2_LVT U4707 ( .A(n6886), .Y(n2862) );
  NBUFFX2_LVT U4708 ( .A(n6886), .Y(n2863) );
  NBUFFX2_LVT U4709 ( .A(n6830), .Y(n2864) );
  NBUFFX2_LVT U4710 ( .A(n6830), .Y(n2865) );
  NBUFFX2_LVT U4711 ( .A(n6763), .Y(n2866) );
  IBUFFX2_LVT U4712 ( .A(n3799), .Y(n2867) );
  IBUFFX2_LVT U4713 ( .A(n3799), .Y(n2868) );
  AND2X1_LVT U4714 ( .A1(n5446), .A2(n2034), .Y(n6763) );
  IBUFFX2_LVT U4715 ( .A(n6763), .Y(n3800) );
  NBUFFX2_LVT U4716 ( .A(n6889), .Y(n2869) );
  NBUFFX2_LVT U4717 ( .A(n6889), .Y(n2870) );
  NBUFFX2_LVT U4718 ( .A(n6829), .Y(n2871) );
  NBUFFX2_LVT U4719 ( .A(n6829), .Y(n2872) );
  AND2X1_LVT U4720 ( .A1(n9417), .A2(n5062), .Y(n2873) );
  AND3X1_LVT U4721 ( .A1(n5395), .A2(n5396), .A3(n406), .Y(n5401) );
  NAND2X0_LVT U4722 ( .A1(n9417), .A2(n5062), .Y(n2874) );
  AND2X1_LVT U4723 ( .A1(n406), .A2(n9383), .Y(N744) );
  AND2X1_LVT U4724 ( .A1(n2873), .A2(n9382), .Y(N745) );
  AND2X1_LVT U4725 ( .A1(n9286), .A2(n2873), .Y(io_fpu_valid) );
  AND2X1_LVT U4726 ( .A1(n9417), .A2(n5062), .Y(n406) );
  NBUFFX2_LVT U4727 ( .A(ibuf_io_inst_0_bits_inst_rs1[1]), .Y(n2876) );
  NBUFFX2_LVT U4728 ( .A(ibuf_io_inst_0_bits_inst_rs1[1]), .Y(n2877) );
  NBUFFX2_LVT U4729 ( .A(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(n2878) );
  NBUFFX2_LVT U4730 ( .A(n6888), .Y(n2879) );
  AND2X1_LVT U4731 ( .A1(n5444), .A2(n5445), .Y(n2881) );
  IBUFFX2_LVT U4732 ( .A(n3012), .Y(n2882) );
  AND3X1_LVT U4733 ( .A1(n6986), .A2(n6985), .A3(n6984), .Y(n2883) );
  AND3X1_LVT U4734 ( .A1(n6982), .A2(n6981), .A3(n6980), .Y(n2884) );
  INVX1_LVT U4735 ( .A(n6766), .Y(n6868) );
  AND3X1_LVT U4736 ( .A1(n7118), .A2(n7117), .A3(n7116), .Y(n2885) );
  AND3X1_LVT U4737 ( .A1(n7114), .A2(n7113), .A3(n7112), .Y(n2886) );
  AND3X1_LVT U4738 ( .A1(n7397), .A2(n7396), .A3(n7395), .Y(n2887) );
  AND3X1_LVT U4739 ( .A1(n7393), .A2(n7392), .A3(n7391), .Y(n2888) );
  AND3X1_LVT U4740 ( .A1(n7312), .A2(n7311), .A3(n7310), .Y(n2889) );
  AND3X1_LVT U4741 ( .A1(n7308), .A2(n7307), .A3(n7306), .Y(n2890) );
  AND3X1_LVT U4742 ( .A1(n7256), .A2(n7255), .A3(n7254), .Y(n2891) );
  AND3X1_LVT U4743 ( .A1(n7252), .A2(n7251), .A3(n7250), .Y(n2892) );
  AND3X1_LVT U4744 ( .A1(n7230), .A2(n7229), .A3(n7228), .Y(n2893) );
  AND3X1_LVT U4745 ( .A1(n7226), .A2(n7225), .A3(n7224), .Y(n2894) );
  AND3X1_LVT U4746 ( .A1(n7058), .A2(n7057), .A3(n7056), .Y(n2895) );
  AND3X1_LVT U4747 ( .A1(n7054), .A2(n7053), .A3(n7052), .Y(n2896) );
  AND3X1_LVT U4748 ( .A1(n6988), .A2(n6989), .A3(n6990), .Y(n2898) );
  AND3X1_LVT U4749 ( .A1(n7014), .A2(n7013), .A3(n7012), .Y(n2899) );
  AND3X1_LVT U4750 ( .A1(n6998), .A2(n6997), .A3(n6996), .Y(n2900) );
  NAND3X0_LVT U4751 ( .A1(n2901), .A2(n2902), .A3(n2903), .Y(N673) );
  AND3X1_LVT U4752 ( .A1(n2953), .A2(n2954), .A3(n2955), .Y(n2901) );
  AND3X1_LVT U4753 ( .A1(n6929), .A2(n6928), .A3(n6927), .Y(n2902) );
  AND3X1_LVT U4754 ( .A1(n6921), .A2(n6920), .A3(n6919), .Y(n2903) );
  AND3X1_LVT U4755 ( .A1(n7368), .A2(n7367), .A3(n7366), .Y(n2904) );
  AND3X1_LVT U4756 ( .A1(n7364), .A2(n7363), .A3(n7362), .Y(n2905) );
  AND3X1_LVT U4757 ( .A1(n7146), .A2(n7145), .A3(n7144), .Y(n2906) );
  AND3X1_LVT U4758 ( .A1(n7142), .A2(n7141), .A3(n7140), .Y(n2907) );
  AND3X1_LVT U4759 ( .A1(n7030), .A2(n7029), .A3(n7028), .Y(n2908) );
  AND3X1_LVT U4760 ( .A1(n7026), .A2(n7025), .A3(n7024), .Y(n2909) );
  AND3X1_LVT U4761 ( .A1(n8733), .A2(n8732), .A3(n8731), .Y(n2911) );
  AND4X1_LVT U4762 ( .A1(n2912), .A2(n2913), .A3(n2914), .A4(n2915), .Y(n5463)
         );
  OA22X1_LVT U4763 ( .A1(n1994), .A2(n3633), .A3(n3256), .A4(n3799), .Y(n2912)
         );
  AOI22X1_LVT U4764 ( .A1(n3828), .A2(n_T_427[1791]), .A3(n_T_427[1663]), .A4(
        n3824), .Y(n2913) );
  AOI22X1_LVT U4765 ( .A1(n3892), .A2(n_T_427[1535]), .A3(n_T_427[1599]), .A4(
        n3886), .Y(n2914) );
  AOI22X1_LVT U4766 ( .A1(n3924), .A2(n_T_427[1471]), .A3(n_T_427[1343]), .A4(
        n3919), .Y(n2915) );
  AND3X1_LVT U4767 ( .A1(n7341), .A2(n7340), .A3(n7339), .Y(n2916) );
  AND3X1_LVT U4768 ( .A1(n7337), .A2(n7336), .A3(n7335), .Y(n2917) );
  AND3X1_LVT U4769 ( .A1(n7932), .A2(n7931), .A3(n7930), .Y(n2918) );
  AND3X1_LVT U4770 ( .A1(n7928), .A2(n7927), .A3(n7926), .Y(n2919) );
  AND2X1_LVT U4771 ( .A1(n2920), .A2(n2921), .Y(n3741) );
  AND3X1_LVT U4772 ( .A1(n8441), .A2(n8440), .A3(n8439), .Y(n2920) );
  AND3X1_LVT U4773 ( .A1(n8445), .A2(n8444), .A3(n8443), .Y(n2921) );
  NBUFFX2_LVT U4774 ( .A(n9012), .Y(n2922) );
  AND3X1_LVT U4775 ( .A1(n7997), .A2(n7996), .A3(n7995), .Y(n2923) );
  AND3X1_LVT U4776 ( .A1(n8001), .A2(n8000), .A3(n7999), .Y(n2924) );
  AND2X1_LVT U4777 ( .A1(n3623), .A2(n3622), .Y(n2925) );
  AND3X1_LVT U4778 ( .A1(n8030), .A2(n8029), .A3(n8028), .Y(n2926) );
  AND3X1_LVT U4779 ( .A1(n8034), .A2(n8033), .A3(n8032), .Y(n2927) );
  OA22X1_LVT U4780 ( .A1(n2875), .A2(n3654), .A3(n3257), .A4(n3799), .Y(n2928)
         );
  AOI22X1_LVT U4781 ( .A1(n3827), .A2(n_T_427[1664]), .A3(n_T_427[1600]), .A4(
        n3885), .Y(n2929) );
  AOI22X1_LVT U4782 ( .A1(n3891), .A2(n_T_427[1536]), .A3(n_T_427[1408]), .A4(
        n3932), .Y(n2930) );
  AOI22X1_LVT U4783 ( .A1(n3923), .A2(n_T_427[1472]), .A3(n_T_427[1344]), .A4(
        n3917), .Y(n2931) );
  AND3X1_LVT U4784 ( .A1(n8293), .A2(n8292), .A3(n8291), .Y(n2932) );
  AND3X1_LVT U4785 ( .A1(n8289), .A2(n8288), .A3(n8287), .Y(n2933) );
  AND2X1_LVT U4786 ( .A1(n8278), .A2(n8277), .Y(n2934) );
  AND3X1_LVT U4787 ( .A1(n7277), .A2(n7276), .A3(n7275), .Y(n2935) );
  AND3X1_LVT U4788 ( .A1(n7269), .A2(n7268), .A3(n7267), .Y(n2936) );
  AND3X1_LVT U4789 ( .A1(n7243), .A2(n7242), .A3(n7241), .Y(n2937) );
  AND3X1_LVT U4790 ( .A1(n7410), .A2(n7409), .A3(n7408), .Y(n2938) );
  AND3X1_LVT U4791 ( .A1(n7329), .A2(n7328), .A3(n7327), .Y(n2939) );
  AND3X1_LVT U4792 ( .A1(n7333), .A2(n7332), .A3(n7331), .Y(n2940) );
  AND3X1_LVT U4793 ( .A1(n7325), .A2(n7324), .A3(n7323), .Y(n2941) );
  AND3X1_LVT U4794 ( .A1(n7075), .A2(n7074), .A3(n7073), .Y(n2942) );
  AND3X1_LVT U4795 ( .A1(n7079), .A2(n7078), .A3(n7077), .Y(n2943) );
  AND3X1_LVT U4796 ( .A1(n7071), .A2(n7070), .A3(n7069), .Y(n2944) );
  NAND3X0_LVT U4797 ( .A1(n2945), .A2(n2946), .A3(n2947), .Y(N728) );
  AND3X1_LVT U4798 ( .A1(n8487), .A2(n8486), .A3(n8485), .Y(n2946) );
  NOR2X0_LVT U4799 ( .A1(n8497), .A2(n8496), .Y(n2947) );
  AND3X1_LVT U4800 ( .A1(n8249), .A2(n8248), .A3(n8247), .Y(n2948) );
  AND3X1_LVT U4801 ( .A1(n8245), .A2(n8244), .A3(n8243), .Y(n2949) );
  AND2X1_LVT U4802 ( .A1(n8096), .A2(n8095), .Y(n2951) );
  AND3X1_LVT U4803 ( .A1(n8094), .A2(n8092), .A3(n8093), .Y(n2952) );
  AND3X1_LVT U4804 ( .A1(n6944), .A2(n6943), .A3(n6942), .Y(n2953) );
  AND3X1_LVT U4805 ( .A1(n6934), .A2(n6933), .A3(n6932), .Y(n2954) );
  AND3X1_LVT U4806 ( .A1(n6978), .A2(n6977), .A3(n6976), .Y(n2955) );
  AND2X1_LVT U4807 ( .A1(n8345), .A2(n8344), .Y(n2956) );
  AND3X1_LVT U4808 ( .A1(n8343), .A2(n8341), .A3(n8342), .Y(n2957) );
  AND3X1_LVT U4809 ( .A1(n7358), .A2(n7359), .A3(n7360), .Y(n2959) );
  AND3X1_LVT U4810 ( .A1(n7354), .A2(n7353), .A3(n7352), .Y(n2960) );
  AND2X1_LVT U4811 ( .A1(n8478), .A2(n8477), .Y(n2961) );
  AND3X1_LVT U4812 ( .A1(n8476), .A2(n8474), .A3(n8475), .Y(n2962) );
  AND2X1_LVT U4813 ( .A1(n7954), .A2(n7953), .Y(n2964) );
  AND3X1_LVT U4814 ( .A1(n7952), .A2(n7951), .A3(n7950), .Y(n2965) );
  AND3X2_LVT U4815 ( .A1(n3773), .A2(n6946), .A3(n6973), .Y(n2966) );
  NBUFFX2_LVT U4816 ( .A(n9007), .Y(n2967) );
  AND2X1_LVT U4817 ( .A1(n4027), .A2(n8105), .Y(n8991) );
  AND2X1_LVT U4818 ( .A1(n4051), .A2(n8105), .Y(n8944) );
  AND2X1_LVT U4819 ( .A1(n4041), .A2(n8105), .Y(n8994) );
  AND2X1_LVT U4820 ( .A1(n3973), .A2(n8105), .Y(n9059) );
  AND2X4_LVT U4821 ( .A1(n8105), .A2(n3979), .Y(n9056) );
  AND2X1_LVT U4822 ( .A1(n4845), .A2(n4844), .Y(n2968) );
  AND2X1_LVT U4823 ( .A1(n5067), .A2(io_fpu_inst[4]), .Y(n5106) );
  AND3X2_LVT U4824 ( .A1(n6973), .A2(n6926), .A3(n2983), .Y(n9029) );
  NAND2X0_LVT U4825 ( .A1(n7910), .A2(n7911), .Y(n9047) );
  AND3X1_LVT U4826 ( .A1(n7389), .A2(n7388), .A3(n7387), .Y(n2970) );
  AND3X1_LVT U4827 ( .A1(n7383), .A2(n7384), .A3(n7385), .Y(n2971) );
  AND3X1_LVT U4828 ( .A1(n7381), .A2(n7380), .A3(n7379), .Y(n2972) );
  AND3X1_LVT U4829 ( .A1(n7222), .A2(n7221), .A3(n7220), .Y(n2973) );
  AND3X1_LVT U4830 ( .A1(n7214), .A2(n7213), .A3(n7212), .Y(n2974) );
  AND3X1_LVT U4831 ( .A1(n7167), .A2(n7166), .A3(n7165), .Y(n2975) );
  AND3X1_LVT U4832 ( .A1(n7161), .A2(n7162), .A3(n7163), .Y(n2976) );
  AND3X1_LVT U4833 ( .A1(n7159), .A2(n7158), .A3(n7157), .Y(n2977) );
  AND3X1_LVT U4834 ( .A1(n7050), .A2(n7049), .A3(n7048), .Y(n2978) );
  AND3X1_LVT U4835 ( .A1(n7043), .A2(n7042), .A3(n7041), .Y(n2979) );
  OR2X1_LVT U4836 ( .A1(n2069), .A2(n2980), .Y(n8246) );
  AND3X1_LVT U4837 ( .A1(n6964), .A2(n6963), .A3(n2627), .Y(n7910) );
  IBUFFX2_LVT U4838 ( .A(n3012), .Y(n2985) );
  IBUFFX2_LVT U4839 ( .A(n3012), .Y(n2986) );
  AND3X1_LVT U4840 ( .A1(n8954), .A2(n8953), .A3(n8952), .Y(n2988) );
  AND3X1_LVT U4841 ( .A1(n8950), .A2(n8949), .A3(n8948), .Y(n2989) );
  AND2X1_LVT U4842 ( .A1(n2990), .A2(n2991), .Y(n3738) );
  AND3X1_LVT U4843 ( .A1(n8509), .A2(n8508), .A3(n8507), .Y(n2990) );
  AND3X1_LVT U4844 ( .A1(n8505), .A2(n8504), .A3(n8503), .Y(n2991) );
  AND2X1_LVT U4845 ( .A1(n2992), .A2(n2993), .Y(n3034) );
  AND3X1_LVT U4846 ( .A1(n8303), .A2(n8304), .A3(n8305), .Y(n2992) );
  AND3X1_LVT U4847 ( .A1(n8301), .A2(n8300), .A3(n8299), .Y(n2993) );
  AND2X1_LVT U4848 ( .A1(n2994), .A2(n2995), .Y(n3731) );
  AND3X1_LVT U4849 ( .A1(n8827), .A2(n8826), .A3(n8825), .Y(n2994) );
  AND3X1_LVT U4850 ( .A1(n8823), .A2(n8822), .A3(n8821), .Y(n2995) );
  AND2X1_LVT U4851 ( .A1(n2996), .A2(n2997), .Y(n3735) );
  AND3X1_LVT U4852 ( .A1(n8612), .A2(n8611), .A3(n8610), .Y(n2996) );
  AND3X1_LVT U4853 ( .A1(n8608), .A2(n8607), .A3(n8606), .Y(n2997) );
  NBUFFX2_LVT U4854 ( .A(n9008), .Y(n2998) );
  NAND3X0_LVT U4855 ( .A1(n3001), .A2(n3000), .A3(n2999), .Y(N699) );
  AND3X1_LVT U4856 ( .A1(n3680), .A2(n3681), .A3(n3682), .Y(n2999) );
  AND3X1_LVT U4857 ( .A1(n7511), .A2(n7510), .A3(n7509), .Y(n3000) );
  AND3X1_LVT U4858 ( .A1(n7507), .A2(n7506), .A3(n7505), .Y(n3001) );
  NAND3X0_LVT U4859 ( .A1(n3002), .A2(n3003), .A3(n3004), .Y(N709) );
  AND3X1_LVT U4860 ( .A1(n3057), .A2(n3058), .A3(n3059), .Y(n3002) );
  AND3X1_LVT U4861 ( .A1(n7827), .A2(n7826), .A3(n7825), .Y(n3003) );
  AND3X1_LVT U4862 ( .A1(n7823), .A2(n7822), .A3(n7821), .Y(n3004) );
  AND3X1_LVT U4863 ( .A1(n7856), .A2(n7855), .A3(n7854), .Y(n3005) );
  AND3X1_LVT U4864 ( .A1(n7852), .A2(n7851), .A3(n7850), .Y(n3006) );
  AND3X1_LVT U4865 ( .A1(n7478), .A2(n7477), .A3(n7476), .Y(n3007) );
  AND3X1_LVT U4866 ( .A1(n7474), .A2(n7473), .A3(n7472), .Y(n3008) );
  NAND3X0_LVT U4867 ( .A1(n3011), .A2(n3010), .A3(n3009), .Y(N703) );
  AND3X1_LVT U4868 ( .A1(n3066), .A2(n3067), .A3(n3068), .Y(n3009) );
  AND3X1_LVT U4869 ( .A1(n7634), .A2(n7633), .A3(n7632), .Y(n3010) );
  AND3X1_LVT U4870 ( .A1(n7630), .A2(n7629), .A3(n7628), .Y(n3011) );
  OA22X1_LVT U4871 ( .A1(n3993), .A2(n3524), .A3(n3178), .A4(n3988), .Y(n3568)
         );
  AND3X1_LVT U4872 ( .A1(n7697), .A2(n7696), .A3(n7695), .Y(n3013) );
  AND3X1_LVT U4873 ( .A1(n7693), .A2(n7692), .A3(n7691), .Y(n3014) );
  AND3X1_LVT U4874 ( .A1(n7730), .A2(n7729), .A3(n7728), .Y(n3015) );
  AND3X1_LVT U4875 ( .A1(n7726), .A2(n7725), .A3(n7724), .Y(n3016) );
  NAND3X0_LVT U4876 ( .A1(n3017), .A2(n3018), .A3(n3019), .Y(N700) );
  AND3X1_LVT U4877 ( .A1(n7540), .A2(n7539), .A3(n7538), .Y(n3018) );
  AND3X1_LVT U4878 ( .A1(n7536), .A2(n7535), .A3(n7534), .Y(n3019) );
  AND3X1_LVT U4879 ( .A1(n7450), .A2(n7449), .A3(n7448), .Y(n3020) );
  AND3X1_LVT U4880 ( .A1(n7446), .A2(n7445), .A3(n7444), .Y(n3021) );
  AND3X1_LVT U4881 ( .A1(n7571), .A2(n7570), .A3(n7569), .Y(n3022) );
  AND3X1_LVT U4882 ( .A1(n7567), .A2(n7566), .A3(n7565), .Y(n3023) );
  AND2X1_LVT U4883 ( .A1(n3024), .A2(n3025), .Y(n3728) );
  AND3X1_LVT U4884 ( .A1(n8859), .A2(n8858), .A3(n8857), .Y(n3024) );
  AND3X1_LVT U4885 ( .A1(n8861), .A2(n8862), .A3(n8863), .Y(n3025) );
  AND2X1_LVT U4886 ( .A1(n3026), .A2(n3027), .Y(n3748) );
  AND3X1_LVT U4887 ( .A1(n9011), .A2(n9010), .A3(n9009), .Y(n3026) );
  AND3X1_LVT U4888 ( .A1(n9017), .A2(n9018), .A3(n9019), .Y(n3027) );
  NAND3X0_LVT U4889 ( .A1(n3028), .A2(n3029), .A3(n3030), .Y(N702) );
  AND3X1_LVT U4890 ( .A1(n7603), .A2(n7602), .A3(n7601), .Y(n3029) );
  AND3X1_LVT U4891 ( .A1(n7599), .A2(n7598), .A3(n7597), .Y(n3030) );
  NAND2X0_LVT U4892 ( .A1(n9231), .A2(n3031), .Y(n3574) );
  AND2X1_LVT U4893 ( .A1(n3575), .A2(csr_io_status_isa[12]), .Y(n3031) );
  NAND2X0_LVT U4894 ( .A1(n3032), .A2(n3033), .Y(n8774) );
  AND3X1_LVT U4895 ( .A1(n8768), .A2(n8769), .A3(n8767), .Y(n3032) );
  AND3X1_LVT U4896 ( .A1(n8773), .A2(n8772), .A3(n8771), .Y(n3033) );
  NAND3X0_LVT U4897 ( .A1(n3034), .A2(n3036), .A3(n3035), .Y(N723) );
  NOR3X0_LVT U4898 ( .A1(n8329), .A2(n8328), .A3(n8327), .Y(n3036) );
  NAND2X0_LVT U4899 ( .A1(n3037), .A2(n3038), .Y(n8923) );
  AND3X1_LVT U4900 ( .A1(n8918), .A2(n8917), .A3(n8916), .Y(n3037) );
  AND3X1_LVT U4901 ( .A1(n8922), .A2(n8921), .A3(n8920), .Y(n3038) );
  IBUFFX2_LVT U4902 ( .A(n6877), .Y(n3879) );
  IBUFFX2_LVT U4903 ( .A(n3082), .Y(n3826) );
  IBUFFX2_LVT U4904 ( .A(n3082), .Y(n3825) );
  MUX21X1_LVT U4905 ( .A1(n3041), .A2(n5306), .S0(n9381), .Y(n3040) );
  IBUFFX2_LVT U4906 ( .A(n9529), .Y(n3044) );
  AND2X1_LVT U4907 ( .A1(n3044), .A2(n5074), .Y(n9076) );
  NAND3X0_LVT U4908 ( .A1(n4843), .A2(n3044), .A3(n4842), .Y(n4845) );
  NAND3X0_LVT U4909 ( .A1(n9091), .A2(n1867), .A3(n9090), .Y(n9092) );
  IBUFFX2_LVT U4910 ( .A(n5075), .Y(n9075) );
  OR3X1_LVT U4911 ( .A1(reset), .A2(n3046), .A3(n9380), .Y(N746) );
  INVX1_LVT U4912 ( .A(n5905), .Y(n6838) );
  XOR2X1_LVT U4913 ( .A1(n2037), .A2(ibuf_io_inst_0_bits_inst_rs2[2]), .Y(
        n5425) );
  NAND3X0_LVT U4914 ( .A1(n9439), .A2(n2553), .A3(n5097), .Y(n5098) );
  AND3X2_LVT U4915 ( .A1(n6973), .A2(n6931), .A3(n3709), .Y(n9004) );
  AND3X2_LVT U4916 ( .A1(n6973), .A2(n6931), .A3(n3709), .Y(n3613) );
  XOR2X1_LVT U4917 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n2574), .Y(
        n5431) );
  MUX21X1_LVT U4918 ( .A1(n3199), .A2(n5426), .S0(n9381), .Y(n9403) );
  MUX21X1_LVT U4919 ( .A1(n3198), .A2(n5428), .S0(n9381), .Y(n9398) );
  AND2X1_LVT U4920 ( .A1(n4971), .A2(n4752), .Y(n6972) );
  INVX1_LVT U4921 ( .A(ibuf_io_inst_0_bits_inst_rs1[2]), .Y(n4752) );
  IBUFFX2_LVT U4922 ( .A(n9522), .Y(n9440) );
  IBUFFX2_LVT U4923 ( .A(n5099), .Y(n5138) );
  AND3X1_LVT U4924 ( .A1(n8958), .A2(n8957), .A3(n8956), .Y(n3050) );
  NOR2X4_LVT U4925 ( .A1(n2552), .A2(n9528), .Y(n9107) );
  AOI22X1_LVT U4926 ( .A1(n2570), .A2(io_fpu_inst[13]), .A3(io_fpu_inst[5]), 
        .A4(n9107), .Y(n4844) );
  IBUFFX2_LVT U4927 ( .A(n9526), .Y(n9105) );
  IBUFFX2_LVT U4928 ( .A(n9107), .Y(n9096) );
  AO22X1_LVT U4929 ( .A1(n5173), .A2(n5174), .A3(n9107), .A4(n9097), .Y(
        id_ctrl_wfd) );
  AND3X1_LVT U4930 ( .A1(n7802), .A2(n7801), .A3(n7800), .Y(n3051) );
  AND3X1_LVT U4931 ( .A1(n7815), .A2(n7813), .A3(n7814), .Y(n3052) );
  AND3X1_LVT U4932 ( .A1(n7798), .A2(n7797), .A3(n7796), .Y(n3053) );
  AND3X1_LVT U4933 ( .A1(n7890), .A2(n7889), .A3(n7888), .Y(n3054) );
  AND3X1_LVT U4934 ( .A1(n7903), .A2(n7902), .A3(n7901), .Y(n3055) );
  AND3X1_LVT U4935 ( .A1(n7886), .A2(n7885), .A3(n7884), .Y(n3056) );
  AND3X1_LVT U4936 ( .A1(n7835), .A2(n7834), .A3(n7833), .Y(n3057) );
  AND3X1_LVT U4937 ( .A1(n7831), .A2(n7830), .A3(n7829), .Y(n3058) );
  AND3X1_LVT U4938 ( .A1(n7848), .A2(n7847), .A3(n7846), .Y(n3059) );
  XNOR2X1_LVT U4939 ( .A1(n4813), .A2(n9390), .Y(n5424) );
  AND3X1_LVT U4940 ( .A1(n7770), .A2(n7769), .A3(n7768), .Y(n3061) );
  AND3X1_LVT U4941 ( .A1(n7783), .A2(n7782), .A3(n7781), .Y(n3062) );
  AND3X1_LVT U4942 ( .A1(n7766), .A2(n7765), .A3(n7764), .Y(n3063) );
  AND3X1_LVT U4943 ( .A1(n7875), .A2(n7874), .A3(n7873), .Y(n3064) );
  AND3X1_LVT U4944 ( .A1(n7859), .A2(n7858), .A3(n7857), .Y(n3065) );
  AND3X1_LVT U4945 ( .A1(n7642), .A2(n7641), .A3(n7640), .Y(n3066) );
  AND3X1_LVT U4946 ( .A1(n7655), .A2(n7654), .A3(n7653), .Y(n3067) );
  AND3X1_LVT U4947 ( .A1(n7638), .A2(n7637), .A3(n7636), .Y(n3068) );
  AND3X1_LVT U4948 ( .A1(n7486), .A2(n7485), .A3(n7484), .Y(n3069) );
  AND3X1_LVT U4949 ( .A1(n7499), .A2(n7498), .A3(n7497), .Y(n3070) );
  AND3X1_LVT U4950 ( .A1(n7482), .A2(n7481), .A3(n7480), .Y(n3071) );
  NAND2X0_LVT U4951 ( .A1(n4844), .A2(n4845), .Y(n3073) );
  NBUFFX2_LVT U4952 ( .A(n9524), .Y(io_fpu_inst[13]) );
  NAND3X2_LVT U4953 ( .A1(n2068), .A2(n6931), .A3(n3709), .Y(n9006) );
  AND3X2_LVT U4954 ( .A1(n6975), .A2(n6931), .A3(n2068), .Y(n3692) );
  AND2X1_LVT U4955 ( .A1(n3044), .A2(n5106), .Y(n9231) );
  INVX1_LVT U4956 ( .A(n9521), .Y(n9438) );
  IBUFFX2_LVT U4957 ( .A(n2981), .Y(n3877) );
  IBUFFX2_LVT U4958 ( .A(n6877), .Y(n3878) );
  MUX21X1_LVT U4959 ( .A1(n5249), .A2(div_io_resp_bits_tag[3]), .S0(n5403), 
        .Y(n5426) );
  MUX21X1_LVT U4960 ( .A1(n5228), .A2(div_io_resp_bits_tag[4]), .S0(n5403), 
        .Y(n5428) );
  MUX21X1_LVT U4961 ( .A1(n5185), .A2(div_io_resp_bits_tag[1]), .S0(n5403), 
        .Y(n5423) );
  MUX21X1_LVT U4962 ( .A1(io_fpu_dmem_resp_tag[0]), .A2(
        div_io_resp_bits_tag[0]), .S0(n5403), .Y(n5306) );
  INVX1_LVT U4963 ( .A(n3883), .Y(n3880) );
  NAND4X1_LVT U4964 ( .A1(n9114), .A2(io_fpu_inst[5]), .A3(n9113), .A4(n9112), 
        .Y(n9115) );
  INVX1_LVT U4965 ( .A(n3803), .Y(n3801) );
  INVX1_LVT U4966 ( .A(n3803), .Y(n3802) );
  INVX1_LVT U4967 ( .A(n3803), .Y(n6764) );
  XOR2X1_LVT U4968 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n9398), .Y(
        n5429) );
  MUX21X1_LVT U4969 ( .A1(n3103), .A2(n5423), .S0(n9381), .Y(n9390) );
  IBUFFX2_LVT U4970 ( .A(n6878), .Y(n3883) );
  IBUFFX2_LVT U4971 ( .A(io_dmem_resp_bits_tag[0]), .Y(n4685) );
  IBUFFX2_LVT U4972 ( .A(n3799), .Y(n3798) );
  IBUFFX2_LVT U4973 ( .A(n9028), .Y(n3717) );
  IBUFFX2_LVT U4974 ( .A(n9028), .Y(n4014) );
  IBUFFX2_LVT U4975 ( .A(n9028), .Y(n3716) );
  NAND3X2_LVT U4976 ( .A1(n6974), .A2(n6973), .A3(n6941), .Y(n9028) );
  IBUFFX2_LVT U4977 ( .A(n2069), .Y(n3744) );
  NBUFFX2_LVT U4978 ( .A(n9518), .Y(n3078) );
  NBUFFX2_LVT U4979 ( .A(n9518), .Y(n3079) );
  INVX1_LVT U4980 ( .A(ibuf_io_inst_0_bits_inst_rs2[1]), .Y(n4813) );
  XOR2X1_LVT U4981 ( .A1(n3781), .A2(n9403), .Y(n5432) );
  IBUFFX2_LVT U4982 ( .A(n9036), .Y(n4017) );
  IBUFFX2_LVT U4983 ( .A(n3012), .Y(n3991) );
  IBUFFX2_LVT U4984 ( .A(n9036), .Y(n4016) );
  IBUFFX2_LVT U4985 ( .A(n2825), .Y(n6956) );
  IBUFFX2_LVT U4986 ( .A(n9523), .Y(n9445) );
  IBUFFX2_LVT U4987 ( .A(n9047), .Y(n3683) );
  IBUFFX2_LVT U4988 ( .A(n9047), .Y(n4053) );
  INVX1_LVT U4989 ( .A(n3658), .Y(n4007) );
  INVX1_LVT U4990 ( .A(n3658), .Y(n4006) );
  INVX1_LVT U4991 ( .A(n3715), .Y(n3747) );
  IBUFFX2_LVT U4992 ( .A(n3012), .Y(n3992) );
  IBUFFX2_LVT U4993 ( .A(n3683), .Y(n3632) );
  IBUFFX2_LVT U4994 ( .A(n3683), .Y(n3656) );
  IBUFFX2_LVT U4995 ( .A(n9529), .Y(n9104) );
  NAND3X2_LVT U4996 ( .A1(n2068), .A2(n6957), .A3(n3709), .Y(n3653) );
  AND3X2_LVT U4997 ( .A1(n3773), .A2(n6948), .A3(n6940), .Y(n9022) );
  IBUFFX2_LVT U4998 ( .A(n6763), .Y(n3799) );
  AND2X1_LVT U4999 ( .A1(n5450), .A2(ibuf_io_inst_0_bits_inst_rs2[3]), .Y(
        n6794) );
  IBUFFX2_LVT U5000 ( .A(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(n3782) );
  IBUFFX2_LVT U5001 ( .A(n4040), .Y(n4036) );
  NBUFFX2_LVT U5002 ( .A(net34650), .Y(n4080) );
  NBUFFX2_LVT U5003 ( .A(net34650), .Y(n4082) );
  NBUFFX2_LVT U5004 ( .A(net34650), .Y(n4084) );
  NBUFFX2_LVT U5005 ( .A(net34650), .Y(n4081) );
  NBUFFX2_LVT U5006 ( .A(net34650), .Y(n4083) );
  NBUFFX2_LVT U5007 ( .A(net34535), .Y(n4223) );
  NBUFFX2_LVT U5008 ( .A(net34575), .Y(n4173) );
  NBUFFX2_LVT U5009 ( .A(net34535), .Y(n4222) );
  NBUFFX2_LVT U5010 ( .A(net34535), .Y(n4219) );
  NBUFFX2_LVT U5011 ( .A(net34535), .Y(n4221) );
  NBUFFX2_LVT U5012 ( .A(net34535), .Y(n4220) );
  NBUFFX2_LVT U5013 ( .A(net34565), .Y(n4183) );
  NBUFFX2_LVT U5014 ( .A(net34525), .Y(n4234) );
  NBUFFX2_LVT U5015 ( .A(net34525), .Y(n4235) );
  NBUFFX2_LVT U5016 ( .A(net34565), .Y(n4184) );
  NBUFFX2_LVT U5017 ( .A(net34565), .Y(n4185) );
  NBUFFX2_LVT U5018 ( .A(net34565), .Y(n4187) );
  NBUFFX2_LVT U5019 ( .A(net34565), .Y(n4186) );
  NBUFFX2_LVT U5020 ( .A(net34575), .Y(n4174) );
  NBUFFX2_LVT U5021 ( .A(net34575), .Y(n4175) );
  NBUFFX2_LVT U5022 ( .A(net34525), .Y(n4231) );
  NBUFFX2_LVT U5023 ( .A(net34570), .Y(n4177) );
  NBUFFX2_LVT U5024 ( .A(net34555), .Y(n4195) );
  NBUFFX2_LVT U5025 ( .A(net34525), .Y(n4232) );
  NBUFFX2_LVT U5026 ( .A(net34570), .Y(n4178) );
  NBUFFX2_LVT U5027 ( .A(net34570), .Y(n4179) );
  NBUFFX2_LVT U5028 ( .A(net34570), .Y(n4180) );
  NBUFFX2_LVT U5029 ( .A(net34525), .Y(n4233) );
  NBUFFX2_LVT U5030 ( .A(net34570), .Y(n4181) );
  NBUFFX2_LVT U5031 ( .A(net34545), .Y(n4210) );
  NBUFFX2_LVT U5032 ( .A(net34615), .Y(n4123) );
  NBUFFX2_LVT U5033 ( .A(net34615), .Y(n4124) );
  NBUFFX2_LVT U5034 ( .A(net34615), .Y(n4125) );
  NBUFFX2_LVT U5035 ( .A(net34555), .Y(n4198) );
  NBUFFX2_LVT U5036 ( .A(net34615), .Y(n4126) );
  NBUFFX2_LVT U5037 ( .A(net34615), .Y(n4127) );
  NBUFFX2_LVT U5038 ( .A(net34555), .Y(n4197) );
  NBUFFX2_LVT U5039 ( .A(net34545), .Y(n4209) );
  NBUFFX2_LVT U5040 ( .A(net34555), .Y(n4196) );
  NBUFFX2_LVT U5041 ( .A(net34605), .Y(n4135) );
  NBUFFX2_LVT U5042 ( .A(net34605), .Y(n4136) );
  NBUFFX2_LVT U5043 ( .A(net34605), .Y(n4137) );
  NBUFFX2_LVT U5044 ( .A(net34635), .Y(n4102) );
  NBUFFX2_LVT U5045 ( .A(net34635), .Y(n4099) );
  NBUFFX2_LVT U5046 ( .A(net34635), .Y(n4103) );
  NBUFFX2_LVT U5047 ( .A(net34545), .Y(n4208) );
  NBUFFX2_LVT U5048 ( .A(net34635), .Y(n4100) );
  NBUFFX2_LVT U5049 ( .A(net34545), .Y(n4207) );
  NBUFFX2_LVT U5050 ( .A(net34625), .Y(n4111) );
  NBUFFX2_LVT U5051 ( .A(net34625), .Y(n4112) );
  NBUFFX2_LVT U5052 ( .A(net34625), .Y(n4113) );
  NBUFFX2_LVT U5053 ( .A(net34625), .Y(n4114) );
  NBUFFX2_LVT U5054 ( .A(net34625), .Y(n4115) );
  NBUFFX2_LVT U5055 ( .A(net34555), .Y(n4199) );
  NBUFFX2_LVT U5056 ( .A(net34545), .Y(n4211) );
  NBUFFX2_LVT U5057 ( .A(net34635), .Y(n4101) );
  NBUFFX2_LVT U5058 ( .A(net34595), .Y(n4151) );
  NBUFFX2_LVT U5059 ( .A(net34645), .Y(n4089) );
  NBUFFX2_LVT U5060 ( .A(net34645), .Y(n4088) );
  NBUFFX2_LVT U5061 ( .A(net34645), .Y(n4087) );
  NBUFFX2_LVT U5062 ( .A(net34645), .Y(n4086) );
  NBUFFX2_LVT U5063 ( .A(net34585), .Y(n4159) );
  NBUFFX2_LVT U5064 ( .A(net34585), .Y(n4160) );
  NBUFFX2_LVT U5065 ( .A(net34585), .Y(n4161) );
  NBUFFX2_LVT U5066 ( .A(net34585), .Y(n4162) );
  NBUFFX2_LVT U5067 ( .A(net34585), .Y(n4163) );
  NBUFFX2_LVT U5068 ( .A(net34575), .Y(n4171) );
  NBUFFX2_LVT U5069 ( .A(net34575), .Y(n4172) );
  NBUFFX2_LVT U5070 ( .A(net34595), .Y(n4150) );
  NBUFFX2_LVT U5071 ( .A(net34595), .Y(n4149) );
  NBUFFX2_LVT U5072 ( .A(net34595), .Y(n4148) );
  NBUFFX2_LVT U5073 ( .A(net34645), .Y(n4090) );
  NBUFFX2_LVT U5074 ( .A(net34605), .Y(n4138) );
  NBUFFX2_LVT U5075 ( .A(net34605), .Y(n4139) );
  NBUFFX2_LVT U5076 ( .A(net34595), .Y(n4147) );
  NBUFFX2_LVT U5077 ( .A(net34640), .Y(n4098) );
  NAND3X0_LVT U5078 ( .A1(n9244), .A2(n9243), .A3(n9242), .Y(n9245) );
  NBUFFX2_LVT U5079 ( .A(net34540), .Y(n4217) );
  NBUFFX2_LVT U5080 ( .A(net34540), .Y(n4216) );
  NBUFFX2_LVT U5081 ( .A(net34655), .Y(n4078) );
  NBUFFX2_LVT U5082 ( .A(net34520), .Y(n4239) );
  NBUFFX2_LVT U5083 ( .A(net34540), .Y(n4215) );
  NBUFFX2_LVT U5084 ( .A(net34540), .Y(n4214) );
  NBUFFX2_LVT U5085 ( .A(net34530), .Y(n4228) );
  NBUFFX2_LVT U5086 ( .A(net34530), .Y(n4227) );
  NBUFFX2_LVT U5087 ( .A(net34530), .Y(n4226) );
  NBUFFX2_LVT U5088 ( .A(net34530), .Y(n4229) );
  NBUFFX2_LVT U5089 ( .A(net34530), .Y(n4225) );
  NBUFFX2_LVT U5090 ( .A(net34655), .Y(n4076) );
  NBUFFX2_LVT U5091 ( .A(net34655), .Y(n4074) );
  NBUFFX2_LVT U5092 ( .A(net34520), .Y(n4241) );
  NBUFFX2_LVT U5093 ( .A(net34655), .Y(n4077) );
  NBUFFX2_LVT U5094 ( .A(net34655), .Y(n4075) );
  NBUFFX2_LVT U5095 ( .A(net34560), .Y(n4190) );
  NBUFFX2_LVT U5096 ( .A(net34600), .Y(n4145) );
  NBUFFX2_LVT U5097 ( .A(net34560), .Y(n4191) );
  NBUFFX2_LVT U5098 ( .A(net34600), .Y(n4144) );
  NBUFFX2_LVT U5099 ( .A(net34600), .Y(n4143) );
  NBUFFX2_LVT U5100 ( .A(net34560), .Y(n4192) );
  NBUFFX2_LVT U5101 ( .A(net34600), .Y(n4142) );
  NBUFFX2_LVT U5102 ( .A(net34600), .Y(n4141) );
  NBUFFX2_LVT U5103 ( .A(net34560), .Y(n4193) );
  NBUFFX2_LVT U5104 ( .A(net34610), .Y(n4133) );
  NBUFFX2_LVT U5105 ( .A(net34610), .Y(n4132) );
  NBUFFX2_LVT U5106 ( .A(net34610), .Y(n4131) );
  NBUFFX2_LVT U5107 ( .A(net34580), .Y(n4167) );
  NBUFFX2_LVT U5108 ( .A(net34580), .Y(n4166) );
  NBUFFX2_LVT U5109 ( .A(net34580), .Y(n4165) );
  NBUFFX2_LVT U5110 ( .A(net34630), .Y(n4105) );
  NBUFFX2_LVT U5111 ( .A(net34630), .Y(n4106) );
  NBUFFX2_LVT U5112 ( .A(net34580), .Y(n4169) );
  NBUFFX2_LVT U5113 ( .A(net34580), .Y(n4168) );
  NBUFFX2_LVT U5114 ( .A(net34630), .Y(n4107) );
  NBUFFX2_LVT U5115 ( .A(net34520), .Y(n4240) );
  NBUFFX2_LVT U5116 ( .A(net34590), .Y(n4157) );
  NBUFFX2_LVT U5117 ( .A(net34590), .Y(n4156) );
  NBUFFX2_LVT U5118 ( .A(net34590), .Y(n4155) );
  NBUFFX2_LVT U5119 ( .A(net34630), .Y(n4108) );
  NBUFFX2_LVT U5120 ( .A(net34590), .Y(n4154) );
  NBUFFX2_LVT U5121 ( .A(net34520), .Y(n4238) );
  NBUFFX2_LVT U5122 ( .A(net34630), .Y(n4109) );
  NBUFFX2_LVT U5123 ( .A(net34560), .Y(n4189) );
  NBUFFX2_LVT U5124 ( .A(net34590), .Y(n4153) );
  NBUFFX2_LVT U5125 ( .A(net34520), .Y(n4237) );
  NBUFFX2_LVT U5126 ( .A(net34550), .Y(n4204) );
  NBUFFX2_LVT U5127 ( .A(net34620), .Y(n4119) );
  NBUFFX2_LVT U5128 ( .A(net34550), .Y(n4202) );
  NBUFFX2_LVT U5129 ( .A(net34550), .Y(n4203) );
  NBUFFX2_LVT U5130 ( .A(net34620), .Y(n4120) );
  NBUFFX2_LVT U5131 ( .A(net34620), .Y(n4121) );
  NBUFFX2_LVT U5132 ( .A(net34540), .Y(n4213) );
  NBUFFX2_LVT U5133 ( .A(net34610), .Y(n4130) );
  NBUFFX2_LVT U5134 ( .A(net34610), .Y(n4129) );
  NBUFFX2_LVT U5135 ( .A(net34620), .Y(n4117) );
  NBUFFX2_LVT U5136 ( .A(net34550), .Y(n4201) );
  NBUFFX2_LVT U5137 ( .A(net34550), .Y(n4205) );
  NBUFFX2_LVT U5138 ( .A(net34620), .Y(n4118) );
  NBUFFX2_LVT U5139 ( .A(net34640), .Y(n4093) );
  NBUFFX2_LVT U5140 ( .A(net34640), .Y(n4095) );
  NBUFFX2_LVT U5141 ( .A(net34640), .Y(n4094) );
  NBUFFX2_LVT U5142 ( .A(net34640), .Y(n4096) );
  NBUFFX2_LVT U5143 ( .A(net34640), .Y(n4097) );
  NBUFFX2_LVT U5144 ( .A(net34640), .Y(n4092) );
  MUX21X1_LVT U5145 ( .A1(n9252), .A2(wb_cause[3]), .S0(wb_cause[1]), .Y(n9255) );
  INVX1_LVT U5146 ( .A(n5260), .Y(n5287) );
  OR2X1_LVT U5147 ( .A1(n5259), .A2(n5270), .Y(n5276) );
  OR2X1_LVT U5148 ( .A1(n5259), .A2(n5280), .Y(n5266) );
  INVX1_LVT U5149 ( .A(n9164), .Y(n9144) );
  OR2X1_LVT U5150 ( .A1(io_fpu_dmem_resp_tag[2]), .A2(n5244), .Y(n5237) );
  NBUFFX2_LVT U5151 ( .A(n711), .Y(n4066) );
  NBUFFX2_LVT U5152 ( .A(n711), .Y(n4067) );
  NBUFFX2_LVT U5153 ( .A(n_T_427__T_1136_data[16]), .Y(n4362) );
  NBUFFX2_LVT U5154 ( .A(n_T_427__T_1136_data[16]), .Y(n4363) );
  NBUFFX2_LVT U5155 ( .A(n_T_427__T_1136_data[54]), .Y(n4468) );
  NBUFFX2_LVT U5156 ( .A(n_T_427__T_1136_data[54]), .Y(n4467) );
  NBUFFX2_LVT U5157 ( .A(n_T_427__T_1136_data[36]), .Y(n4415) );
  NBUFFX2_LVT U5158 ( .A(n_T_427__T_1136_data[36]), .Y(n4414) );
  NBUFFX2_LVT U5159 ( .A(n_T_427__T_1136_data[49]), .Y(n4453) );
  NBUFFX2_LVT U5160 ( .A(n_T_427__T_1136_data[52]), .Y(n4462) );
  NBUFFX2_LVT U5161 ( .A(n_T_427__T_1136_data[56]), .Y(n4474) );
  NBUFFX2_LVT U5162 ( .A(n_T_427__T_1136_data[29]), .Y(n4396) );
  NBUFFX2_LVT U5163 ( .A(n_T_427__T_1136_data[30]), .Y(n4399) );
  NBUFFX2_LVT U5164 ( .A(n_T_427__T_1136_data[49]), .Y(n4452) );
  NBUFFX2_LVT U5165 ( .A(n_T_427__T_1136_data[41]), .Y(n4429) );
  NBUFFX2_LVT U5166 ( .A(n_T_427__T_1136_data[29]), .Y(n4397) );
  NBUFFX2_LVT U5167 ( .A(n_T_427__T_1136_data[56]), .Y(n4473) );
  NBUFFX2_LVT U5168 ( .A(n_T_427__T_1136_data[30]), .Y(n4400) );
  NBUFFX2_LVT U5169 ( .A(n_T_427__T_1136_data[41]), .Y(n4428) );
  NBUFFX2_LVT U5170 ( .A(n_T_427__T_1136_data[52]), .Y(n4461) );
  NBUFFX2_LVT U5171 ( .A(n_T_427__T_1136_data[27]), .Y(n4391) );
  NBUFFX2_LVT U5172 ( .A(n_T_427__T_1136_data[27]), .Y(n4392) );
  NBUFFX2_LVT U5173 ( .A(n_T_427__T_1136_data[58]), .Y(n4480) );
  NBUFFX2_LVT U5174 ( .A(n_T_427__T_1136_data[58]), .Y(n4479) );
  NBUFFX2_LVT U5175 ( .A(n_T_427__T_1136_data[62]), .Y(n4491) );
  NBUFFX2_LVT U5176 ( .A(n_T_427__T_1136_data[60]), .Y(n4485) );
  NBUFFX2_LVT U5177 ( .A(n_T_427__T_1136_data[62]), .Y(n4492) );
  NBUFFX2_LVT U5178 ( .A(n_T_427__T_1136_data[60]), .Y(n4486) );
  NBUFFX2_LVT U5179 ( .A(n_T_427__T_1136_data[53]), .Y(n4465) );
  NBUFFX2_LVT U5180 ( .A(n_T_427__T_1136_data[53]), .Y(n4464) );
  NBUFFX2_LVT U5181 ( .A(n_T_427__T_1136_data[59]), .Y(n4483) );
  NBUFFX2_LVT U5182 ( .A(n_T_427__T_1136_data[59]), .Y(n4482) );
  NBUFFX2_LVT U5183 ( .A(n_T_427__T_1136_data[1]), .Y(n4320) );
  NBUFFX2_LVT U5184 ( .A(n_T_427__T_1136_data[1]), .Y(n4319) );
  NBUFFX2_LVT U5185 ( .A(n_T_427__T_1136_data[50]), .Y(n4456) );
  NBUFFX2_LVT U5186 ( .A(n_T_427__T_1136_data[50]), .Y(n4455) );
  NBUFFX2_LVT U5187 ( .A(n_T_427__T_1136_data[61]), .Y(n4489) );
  NBUFFX2_LVT U5188 ( .A(n_T_427__T_1136_data[61]), .Y(n4488) );
  NBUFFX2_LVT U5189 ( .A(n_T_427__T_1136_data[57]), .Y(n4477) );
  NBUFFX2_LVT U5190 ( .A(n_T_427__T_1136_data[55]), .Y(n4470) );
  NBUFFX2_LVT U5191 ( .A(n_T_427__T_1136_data[55]), .Y(n4471) );
  NBUFFX2_LVT U5192 ( .A(n_T_427__T_1136_data[57]), .Y(n4476) );
  NBUFFX2_LVT U5193 ( .A(n_T_427__T_1136_data[19]), .Y(n4372) );
  NBUFFX2_LVT U5194 ( .A(n_T_427__T_1136_data[20]), .Y(n4375) );
  NBUFFX2_LVT U5195 ( .A(n_T_427__T_1136_data[19]), .Y(n4371) );
  NBUFFX2_LVT U5196 ( .A(n_T_427__T_1136_data[24]), .Y(n4385) );
  NBUFFX2_LVT U5197 ( .A(n_T_427__T_1136_data[0]), .Y(n4317) );
  NBUFFX2_LVT U5198 ( .A(n_T_427__T_1136_data[24]), .Y(n4384) );
  NBUFFX2_LVT U5199 ( .A(n_T_427__T_1136_data[0]), .Y(n4316) );
  NBUFFX2_LVT U5200 ( .A(n_T_427__T_1136_data[18]), .Y(n4368) );
  NBUFFX2_LVT U5201 ( .A(n_T_427__T_1136_data[18]), .Y(n4369) );
  NBUFFX2_LVT U5202 ( .A(n_T_427__T_1136_data[20]), .Y(n4374) );
  NBUFFX2_LVT U5203 ( .A(n_T_427__T_1136_data[63]), .Y(n4495) );
  NBUFFX2_LVT U5204 ( .A(n_T_427__T_1136_data[63]), .Y(n4494) );
  NBUFFX2_LVT U5205 ( .A(n_T_427__T_1136_data[37]), .Y(n4417) );
  NBUFFX2_LVT U5206 ( .A(n_T_427__T_1136_data[37]), .Y(n4418) );
  NBUFFX2_LVT U5207 ( .A(n_T_427__T_1136_data[44]), .Y(n4437) );
  NBUFFX2_LVT U5208 ( .A(n_T_427__T_1136_data[32]), .Y(n4404) );
  NBUFFX2_LVT U5209 ( .A(n_T_427__T_1136_data[34]), .Y(n4410) );
  NBUFFX2_LVT U5210 ( .A(n_T_427__T_1136_data[46]), .Y(n4444) );
  NBUFFX2_LVT U5211 ( .A(n_T_427__T_1136_data[46]), .Y(n4443) );
  NBUFFX2_LVT U5212 ( .A(n_T_427__T_1136_data[39]), .Y(n4423) );
  NBUFFX2_LVT U5213 ( .A(n_T_427__T_1136_data[32]), .Y(n4405) );
  NBUFFX2_LVT U5214 ( .A(n_T_427__T_1136_data[44]), .Y(n4438) );
  NBUFFX2_LVT U5215 ( .A(n_T_427__T_1136_data[34]), .Y(n4409) );
  NBUFFX2_LVT U5216 ( .A(n_T_427__T_1136_data[39]), .Y(n4422) );
  NBUFFX2_LVT U5217 ( .A(n_T_427__T_1136_data[17]), .Y(n4365) );
  NBUFFX2_LVT U5218 ( .A(n_T_427__T_1136_data[23]), .Y(n4381) );
  NBUFFX2_LVT U5219 ( .A(n_T_427__T_1136_data[23]), .Y(n4382) );
  NBUFFX2_LVT U5220 ( .A(n_T_427__T_1136_data[17]), .Y(n4366) );
  NBUFFX2_LVT U5221 ( .A(n_T_427__T_1136_data[40]), .Y(n4425) );
  NBUFFX2_LVT U5222 ( .A(n_T_427__T_1136_data[47]), .Y(n4447) );
  NBUFFX2_LVT U5223 ( .A(n_T_427__T_1136_data[48]), .Y(n4450) );
  NBUFFX2_LVT U5224 ( .A(n_T_427__T_1136_data[48]), .Y(n4449) );
  NBUFFX2_LVT U5225 ( .A(n_T_427__T_1136_data[47]), .Y(n4446) );
  NBUFFX2_LVT U5226 ( .A(n_T_427__T_1136_data[40]), .Y(n4426) );
  NBUFFX2_LVT U5227 ( .A(n_T_427__T_1136_data[45]), .Y(n4441) );
  NBUFFX2_LVT U5228 ( .A(n_T_427__T_1136_data[45]), .Y(n4440) );
  NBUFFX2_LVT U5229 ( .A(n_T_427__T_1136_data[51]), .Y(n4458) );
  NBUFFX2_LVT U5230 ( .A(n_T_427__T_1136_data[43]), .Y(n4434) );
  NBUFFX2_LVT U5231 ( .A(n_T_427__T_1136_data[42]), .Y(n4431) );
  NBUFFX2_LVT U5232 ( .A(n_T_427__T_1136_data[51]), .Y(n4459) );
  NBUFFX2_LVT U5233 ( .A(n_T_427__T_1136_data[43]), .Y(n4435) );
  NBUFFX2_LVT U5234 ( .A(n_T_427__T_1136_data[42]), .Y(n4432) );
  AND3X1_LVT U5235 ( .A1(io_imem_bht_update_bits_mispredict), .A2(
        io_imem_bht_update_valid), .A3(n9329), .Y(io_imem_btb_update_valid) );
  NAND3X0_LVT U5236 ( .A1(n9231), .A2(n2618), .A3(n9079), .Y(n9080) );
  XOR2X1_LVT U5237 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n591), .Y(n5032)
         );
  XOR2X1_LVT U5238 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n589), .Y(n5030)
         );
  XOR2X1_LVT U5239 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n592), .Y(n5035)
         );
  XOR2X1_LVT U5240 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n3201), .Y(n5017) );
  XOR2X1_LVT U5241 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n3103), .Y(n5018) );
  XOR2X1_LVT U5242 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n3199), .Y(n5014) );
  XOR2X1_LVT U5243 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n3198), .Y(n5015) );
  XOR2X1_LVT U5244 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n3102), .Y(n5016) );
  NAND4X0_LVT U5245 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n5437), .Y(n4910) );
  NAND4X0_LVT U5246 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n5437), .Y(n4914) );
  OA21X1_LVT U5247 ( .A1(n3264), .A2(n6422), .A3(n5434), .Y(n4883) );
  MUX21X1_LVT U5248 ( .A1(n4812), .A2(n4811), .S0(n2494), .Y(n4839) );
  NAND2X0_LVT U5249 ( .A1(n4782), .A2(ibuf_io_inst_0_bits_raw[27]), .Y(n4803)
         );
  NAND2X0_LVT U5250 ( .A1(n4781), .A2(ibuf_io_inst_0_bits_raw[28]), .Y(n4801)
         );
  XOR2X1_LVT U5251 ( .A1(n2674), .A2(n3200), .Y(n4624) );
  XOR2X1_LVT U5252 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n596), .Y(n4619)
         );
  XOR2X1_LVT U5253 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n595), .Y(n4620)
         );
  XOR2X1_LVT U5254 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n3200), .Y(n4621) );
  INVX1_LVT U5255 ( .A(ibuf_io_pc[34]), .Y(n4557) );
  XOR2X1_LVT U5256 ( .A1(n9484), .A2(ibuf_io_pc[5]), .Y(n4541) );
  XOR2X1_LVT U5257 ( .A1(n9334), .A2(n4532), .Y(n4535) );
  XOR2X1_LVT U5258 ( .A1(n9503), .A2(ibuf_io_pc[3]), .Y(n4537) );
  XOR2X1_LVT U5259 ( .A1(n9499), .A2(ibuf_io_pc[7]), .Y(n4543) );
  INVX1_LVT U5260 ( .A(ibuf_io_pc[16]), .Y(n4518) );
  NBUFFX2_LVT U5261 ( .A(n711), .Y(n4065) );
  OR2X1_LVT U5262 ( .A1(csr_io_exception), .A2(csr_io_eret), .Y(n711) );
  NBUFFX2_LVT U5263 ( .A(n6898), .Y(n3957) );
  NBUFFX2_LVT U5264 ( .A(n6886), .Y(n3908) );
  NBUFFX2_LVT U5265 ( .A(n6838), .Y(n3840) );
  NBUFFX2_LVT U5266 ( .A(n6865), .Y(n3859) );
  NBUFFX2_LVT U5267 ( .A(n6868), .Y(n3867) );
  NBUFFX2_LVT U5268 ( .A(n6870), .Y(n3871) );
  NBUFFX2_LVT U5269 ( .A(n6898), .Y(n3958) );
  INVX1_LVT U5270 ( .A(n5546), .Y(n6870) );
  INVX1_LVT U5271 ( .A(n4814), .Y(n4901) );
  NAND2X0_LVT U5272 ( .A1(n5452), .A2(n2878), .Y(n3083) );
  NBUFFX2_LVT U5273 ( .A(n6715), .Y(n3796) );
  NBUFFX2_LVT U5274 ( .A(n6869), .Y(n3868) );
  NBUFFX2_LVT U5275 ( .A(n6837), .Y(n3836) );
  NAND2X0_LVT U5276 ( .A1(n5449), .A2(n5436), .Y(n6766) );
  NBUFFX2_LVT U5277 ( .A(n6795), .Y(n3812) );
  AND2X1_LVT U5278 ( .A1(n4027), .A2(n2135), .Y(n3661) );
  NBUFFX2_LVT U5279 ( .A(n9038), .Y(n4027) );
  NBUFFX2_LVT U5280 ( .A(n8900), .Y(n3960) );
  NBUFFX2_LVT U5281 ( .A(n8981), .Y(n3979) );
  NBUFFX2_LVT U5282 ( .A(n8932), .Y(n3972) );
  NBUFFX2_LVT U5283 ( .A(n8931), .Y(n3968) );
  NBUFFX2_LVT U5284 ( .A(n8982), .Y(n3983) );
  NBUFFX2_LVT U5285 ( .A(n8980), .Y(n3976) );
  NAND2X0_LVT U5286 ( .A1(n6939), .A2(n6936), .Y(n3625) );
  NBUFFX2_LVT U5287 ( .A(n9042), .Y(n4051) );
  INVX1_LVT U5288 ( .A(n3184), .Y(n4026) );
  INVX1_LVT U5289 ( .A(n6945), .Y(n9042) );
  INVX1_LVT U5290 ( .A(n4017), .Y(n4015) );
  XOR2X1_LVT U5291 ( .A1(ibuf_io_inst_0_bits_inst_rs1[3]), .A2(n9403), .Y(
        n6908) );
  XOR2X1_LVT U5292 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n9398), .Y(
        n6909) );
  XOR2X1_LVT U5293 ( .A1(n3040), .A2(n2098), .Y(n6910) );
  XOR2X1_LVT U5294 ( .A1(n3042), .A2(n2038), .Y(n6911) );
  XOR2X1_LVT U5295 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n588), .Y(n5010) );
  XOR2X1_LVT U5296 ( .A1(ibuf_io_inst_0_bits_inst_rs1[2]), .A2(n590), .Y(n5012) );
  XOR2X1_LVT U5297 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n595), .Y(n4617) );
  OAI21X1_LVT U5298 ( .A1(n2618), .A2(n3079), .A3(n9522), .Y(n3180) );
  XOR2X1_LVT U5299 ( .A1(n9495), .A2(ibuf_io_pc[4]), .Y(n4540) );
  INVX1_LVT U5300 ( .A(ibuf_io_pc[2]), .Y(n4532) );
  XOR2X1_LVT U5301 ( .A1(n9512), .A2(ibuf_io_pc[1]), .Y(n4534) );
  NBUFFX2_LVT U5302 ( .A(n8901), .Y(n3964) );
  OA22X1_LVT U5303 ( .A1(n3269), .A2(n5906), .A3(n3128), .A4(n5905), .Y(n4882)
         );
  AO22X1_LVT U5304 ( .A1(n_T_698[3]), .A2(n9101), .A3(io_fpu_fromint_data[3]), 
        .A4(n9103), .Y(alu_io_in1[3]) );
  AO22X1_LVT U5305 ( .A1(n_T_698[4]), .A2(n9101), .A3(io_fpu_fromint_data[4]), 
        .A4(n9103), .Y(alu_io_in1[4]) );
  AO22X1_LVT U5306 ( .A1(n_T_698[2]), .A2(n4054), .A3(io_fpu_fromint_data[2]), 
        .A4(n9103), .Y(alu_io_in1[2]) );
  AO22X1_LVT U5307 ( .A1(n_T_698[6]), .A2(n4054), .A3(io_fpu_fromint_data[6]), 
        .A4(n9103), .Y(alu_io_in1[6]) );
  AO22X1_LVT U5308 ( .A1(n_T_698[0]), .A2(n9101), .A3(io_fpu_fromint_data[0]), 
        .A4(n9103), .Y(alu_io_in1[0]) );
  AO22X1_LVT U5309 ( .A1(n_T_698[7]), .A2(n4054), .A3(io_fpu_fromint_data[7]), 
        .A4(n9103), .Y(alu_io_in1[7]) );
  AO22X1_LVT U5310 ( .A1(n_T_698[10]), .A2(n4054), .A3(io_fpu_fromint_data[10]), .A4(n9103), .Y(alu_io_in1[10]) );
  AO22X1_LVT U5311 ( .A1(n_T_698[12]), .A2(n4054), .A3(io_fpu_fromint_data[12]), .A4(n9103), .Y(alu_io_in1[12]) );
  AO22X1_LVT U5312 ( .A1(n_T_698[13]), .A2(n4054), .A3(io_fpu_fromint_data[13]), .A4(n9103), .Y(alu_io_in1[13]) );
  AO22X1_LVT U5313 ( .A1(n_T_698[14]), .A2(n4054), .A3(io_fpu_fromint_data[14]), .A4(n9103), .Y(alu_io_in1[14]) );
  AO22X1_LVT U5314 ( .A1(n_T_698[15]), .A2(n4054), .A3(io_fpu_fromint_data[15]), .A4(n9103), .Y(alu_io_in1[15]) );
  AO22X1_LVT U5315 ( .A1(n_T_698[16]), .A2(n4054), .A3(io_fpu_fromint_data[16]), .A4(n9103), .Y(alu_io_in1[16]) );
  AO22X1_LVT U5316 ( .A1(n4054), .A2(n_T_698[17]), .A3(io_fpu_fromint_data[17]), .A4(n9103), .Y(alu_io_in1[17]) );
  AO22X1_LVT U5317 ( .A1(n_T_698[18]), .A2(n4054), .A3(io_fpu_fromint_data[18]), .A4(n9103), .Y(alu_io_in1[18]) );
  AO22X1_LVT U5318 ( .A1(n_T_698[19]), .A2(n4054), .A3(io_fpu_fromint_data[19]), .A4(n9103), .Y(alu_io_in1[19]) );
  AO22X1_LVT U5319 ( .A1(n9101), .A2(n_T_698[20]), .A3(io_fpu_fromint_data[20]), .A4(n9103), .Y(alu_io_in1[20]) );
  AO22X1_LVT U5320 ( .A1(n_T_698[21]), .A2(n9101), .A3(io_fpu_fromint_data[21]), .A4(n9103), .Y(alu_io_in1[21]) );
  AO22X1_LVT U5321 ( .A1(n_T_698[22]), .A2(n9101), .A3(io_fpu_fromint_data[22]), .A4(n9103), .Y(alu_io_in1[22]) );
  AO22X1_LVT U5322 ( .A1(n_T_698[29]), .A2(n4054), .A3(io_fpu_fromint_data[29]), .A4(n9103), .Y(alu_io_in1[29]) );
  AO22X1_LVT U5323 ( .A1(n9101), .A2(n_T_698[30]), .A3(io_fpu_fromint_data[30]), .A4(n9103), .Y(alu_io_in1[30]) );
  AO22X1_LVT U5324 ( .A1(n_T_698[23]), .A2(n9101), .A3(io_fpu_fromint_data[23]), .A4(n9103), .Y(alu_io_in1[23]) );
  AO22X1_LVT U5325 ( .A1(n_T_698[24]), .A2(n9101), .A3(io_fpu_fromint_data[24]), .A4(n9103), .Y(alu_io_in1[24]) );
  AO22X1_LVT U5326 ( .A1(n4054), .A2(n_T_698[33]), .A3(io_fpu_fromint_data[33]), .A4(n9103), .Y(alu_io_in1[33]) );
  AO22X1_LVT U5327 ( .A1(n_T_698[35]), .A2(n9101), .A3(io_fpu_fromint_data[35]), .A4(n9103), .Y(alu_io_in1[35]) );
  AO22X1_LVT U5328 ( .A1(n_T_698[32]), .A2(n9101), .A3(io_fpu_fromint_data[32]), .A4(n9103), .Y(alu_io_in1[32]) );
  AO22X1_LVT U5329 ( .A1(n_T_698[34]), .A2(n4054), .A3(io_fpu_fromint_data[34]), .A4(n9103), .Y(alu_io_in1[34]) );
  AO22X1_LVT U5330 ( .A1(n4054), .A2(n_T_698[36]), .A3(io_fpu_fromint_data[36]), .A4(n9103), .Y(alu_io_in1[36]) );
  AO22X1_LVT U5331 ( .A1(n9101), .A2(n_T_698[37]), .A3(io_fpu_fromint_data[37]), .A4(n9103), .Y(alu_io_in1[37]) );
  AO22X1_LVT U5332 ( .A1(n4054), .A2(n_T_698[38]), .A3(io_fpu_fromint_data[38]), .A4(n9103), .Y(alu_io_in1[38]) );
  NAND2X0_LVT U5333 ( .A1(mem_br_target[39]), .A2(n6249), .Y(n6857) );
  AND2X1_LVT U5334 ( .A1(n5409), .A2(n5410), .Y(n6855) );
  INVX1_LVT U5335 ( .A(n5410), .Y(n6856) );
  AND2X1_LVT U5336 ( .A1(n5407), .A2(n5406), .Y(n6249) );
  INVX1_LVT U5337 ( .A(n9292), .Y(n9301) );
  INVX1_LVT U5338 ( .A(n3234), .Y(n4058) );
  NAND2X0_LVT U5339 ( .A1(io_dmem_req_bits_size[0]), .A2(
        io_dmem_req_bits_size[1]), .Y(n3234) );
  NOR2X0_LVT U5340 ( .A1(io_dmem_req_bits_size[1]), .A2(
        io_dmem_req_bits_size[0]), .Y(n9291) );
  OR2X1_LVT U5341 ( .A1(io_fpu_sboard_clra[4]), .A2(io_fpu_sboard_clra[3]), 
        .Y(n5193) );
  MUX21X1_LVT U5342 ( .A1(n7016), .A2(io_fpu_dmem_resp_data[0]), .S0(n9064), 
        .Y(io_fpu_fromint_data[0]) );
  OR2X1_LVT U5343 ( .A1(n9201), .A2(n9173), .Y(n9164) );
  OR2X1_LVT U5344 ( .A1(n9201), .A2(n9172), .Y(n9163) );
  OR2X1_LVT U5345 ( .A1(ex_ctrl_sel_imm[2]), .A2(n546), .Y(n9178) );
  AND3X1_LVT U5346 ( .A1(n9173), .A2(n9179), .A3(ex_reg_inst_31_), .Y(n9226)
         );
  AND2X1_LVT U5347 ( .A1(n9101), .A2(n_T_698[39]), .Y(n9102) );
  NOR2X0_LVT U5348 ( .A1(ex_ctrl_sel_alu1_0_), .A2(n561), .Y(n9101) );
  AND2X1_LVT U5349 ( .A1(n561), .A2(ex_ctrl_sel_alu1_0_), .Y(n9103) );
  MUX21X1_LVT U5350 ( .A1(io_fpu_inst[3]), .A2(io_fpu_inst[2]), .S0(n2553), 
        .Y(id_ctrl_sel_imm[1]) );
  INVX1_LVT U5351 ( .A(n5282), .Y(n5381) );
  INVX1_LVT U5352 ( .A(n5272), .Y(n5365) );
  AND2X1_LVT U5353 ( .A1(n5210), .A2(n3043), .Y(n5317) );
  AND2X1_LVT U5354 ( .A1(n5227), .A2(wb_waddr[3]), .Y(n5382) );
  INVX1_LVT U5355 ( .A(n5298), .Y(n5362) );
  INVX1_LVT U5356 ( .A(ex_reg_rs_bypass_1), .Y(n6901) );
  AND2X1_LVT U5357 ( .A1(n5484), .A2(ex_reg_rs_bypass_1), .Y(n6900) );
  AND2X1_LVT U5358 ( .A1(n7017), .A2(n569), .Y(n9065) );
  OR2X1_LVT U5359 ( .A1(mem_reg_xcpt), .A2(mem_reg_xcpt_interrupt), .Y(n1279)
         );
  MUX21X1_LVT U5360 ( .A1(io_fpu_inst[13]), .A2(n5421), .S0(n9287), .Y(N370)
         );
  MUX21X1_LVT U5361 ( .A1(n2618), .A2(n9288), .S0(n9287), .Y(N369) );
  MUX21X1_LVT U5362 ( .A1(n3226), .A2(n4592), .S0(n3792), .Y(n9505) );
  MUX21X1_LVT U5363 ( .A1(n3219), .A2(n4586), .S0(n3792), .Y(n9492) );
  MUX21X1_LVT U5364 ( .A1(n3110), .A2(n4581), .S0(n3792), .Y(n9497) );
  MUX21X1_LVT U5365 ( .A1(n3210), .A2(n4580), .S0(n4591), .Y(n9493) );
  MUX21X1_LVT U5366 ( .A1(n3216), .A2(n4579), .S0(n3792), .Y(n9501) );
  MUX21X1_LVT U5367 ( .A1(n3224), .A2(n4578), .S0(n3792), .Y(n9486) );
  MUX21X1_LVT U5368 ( .A1(n_T_918[28]), .A2(mem_br_target[28]), .S0(n3792), 
        .Y(n9368) );
  MUX21X1_LVT U5369 ( .A1(n_T_918[24]), .A2(mem_br_target[24]), .S0(n3792), 
        .Y(n9364) );
  MUX21X1_LVT U5370 ( .A1(n4573), .A2(mem_br_target[39]), .S0(n3792), .Y(n9377) );
  MUX21X1_LVT U5371 ( .A1(n3212), .A2(n4572), .S0(n3792), .Y(n9510) );
  MUX21X1_LVT U5372 ( .A1(n_T_918[21]), .A2(mem_br_target[21]), .S0(n3792), 
        .Y(n9361) );
  MUX21X1_LVT U5373 ( .A1(n3211), .A2(n4571), .S0(n3792), .Y(n9490) );
  MUX21X1_LVT U5374 ( .A1(n3106), .A2(n4570), .S0(n3792), .Y(n9500) );
  MUX21X1_LVT U5375 ( .A1(n3225), .A2(n4569), .S0(n3792), .Y(n9509) );
  MUX21X1_LVT U5376 ( .A1(n_T_918[15]), .A2(mem_br_target[15]), .S0(n3792), 
        .Y(n9355) );
  MUX21X1_LVT U5377 ( .A1(n3111), .A2(n4568), .S0(n3792), .Y(n9504) );
  MUX21X1_LVT U5378 ( .A1(n3528), .A2(n4567), .S0(n3792), .Y(n9494) );
  MUX21X1_LVT U5379 ( .A1(n3105), .A2(n4562), .S0(n4591), .Y(n9502) );
  MUX21X1_LVT U5380 ( .A1(n_T_918[34]), .A2(mem_br_target[34]), .S0(n3792), 
        .Y(n9373) );
  MUX21X1_LVT U5381 ( .A1(n3107), .A2(n4550), .S0(n4591), .Y(n9487) );
  MUX21X1_LVT U5382 ( .A1(n3207), .A2(n4533), .S0(n4591), .Y(n9512) );
  MUX21X1_LVT U5383 ( .A1(n3221), .A2(n4527), .S0(n4591), .Y(n9491) );
  MUX21X1_LVT U5384 ( .A1(n3223), .A2(n4526), .S0(n3792), .Y(n9506) );
  MUX21X1_LVT U5385 ( .A1(n3220), .A2(n4525), .S0(n4591), .Y(n9496) );
  MUX21X1_LVT U5386 ( .A1(n3213), .A2(n4524), .S0(n3792), .Y(n9488) );
  MUX21X1_LVT U5387 ( .A1(n3209), .A2(n4523), .S0(n4591), .Y(n9489) );
  MUX21X1_LVT U5388 ( .A1(n3227), .A2(n4522), .S0(n3792), .Y(n9508) );
  MUX21X1_LVT U5389 ( .A1(n3218), .A2(n4517), .S0(n3792), .Y(n9483) );
  NBUFFX2_LVT U5390 ( .A(n4591), .Y(n3792) );
  MUX21X1_LVT U5391 ( .A1(n3205), .A2(n4516), .S0(n4591), .Y(n9498) );
  AND2X1_LVT U5392 ( .A1(n3230), .A2(n5080), .Y(n5083) );
  AND2X1_LVT U5393 ( .A1(n_T_844_10_), .A2(n5082), .Y(n9427) );
  NAND3X2_LVT U5394 ( .A1(n2068), .A2(n6972), .A3(n3709), .Y(n3684) );
  NAND3X2_LVT U5395 ( .A1(n6975), .A2(n6957), .A3(n2068), .Y(n3658) );
  NAND3X2_LVT U5396 ( .A1(n3773), .A2(n6954), .A3(n2068), .Y(n3601) );
  OR2X2_LVT U5397 ( .A1(n9113), .A2(n9104), .Y(n1699) );
  OR2X2_LVT U5398 ( .A1(n4848), .A2(n4847), .Y(n6991) );
  NAND2X0_LVT U5399 ( .A1(n5408), .A2(n3251), .Y(n5410) );
  NBUFFX2_LVT U5400 ( .A(net34475), .Y(n4311) );
  NBUFFX2_LVT U5401 ( .A(n9276), .Y(n4056) );
  NBUFFX2_LVT U5402 ( .A(n9276), .Y(n4057) );
  NBUFFX2_LVT U5403 ( .A(n9276), .Y(n4055) );
  NBUFFX2_LVT U5404 ( .A(n5296), .Y(n3794) );
  NBUFFX2_LVT U5405 ( .A(n5296), .Y(n3793) );
  AND2X1_LVT U5406 ( .A1(n4498), .A2(n9379), .Y(n5296) );
  NBUFFX2_LVT U5407 ( .A(n9378), .Y(n4059) );
  NBUFFX2_LVT U5408 ( .A(n9414), .Y(n4062) );
  NBUFFX2_LVT U5409 ( .A(n9378), .Y(n4060) );
  NBUFFX2_LVT U5410 ( .A(n9414), .Y(n4063) );
  NBUFFX2_LVT U5411 ( .A(n9378), .Y(n4061) );
  NBUFFX2_LVT U5412 ( .A(n9414), .Y(n4064) );
  NAND2X0_LVT U5413 ( .A1(n5481), .A2(n_T_635[1]), .Y(n5483) );
  OR2X1_LVT U5414 ( .A1(n9330), .A2(n4065), .Y(n9332) );
  NBUFFX2_LVT U5415 ( .A(n6860), .Y(n3853) );
  AND3X2_LVT U5416 ( .A1(n3709), .A2(n6957), .A3(n6940), .Y(n3770) );
  NBUFFX2_LVT U5417 ( .A(n6861), .Y(n3857) );
  NBUFFX2_LVT U5418 ( .A(n6859), .Y(n3847) );
  NBUFFX2_LVT U5419 ( .A(n6861), .Y(n3854) );
  NBUFFX2_LVT U5420 ( .A(n6859), .Y(n3846) );
  NBUFFX2_LVT U5421 ( .A(n6861), .Y(n3856) );
  NBUFFX2_LVT U5422 ( .A(n6860), .Y(n3852) );
  NBUFFX2_LVT U5423 ( .A(n6861), .Y(n3855) );
  AND2X1_LVT U5424 ( .A1(n5411), .A2(n5415), .Y(n6858) );
  AND2X1_LVT U5425 ( .A1(n5412), .A2(n5413), .Y(n5411) );
  OR3X1_LVT U5426 ( .A1(wb_ctrl_csr[1]), .A2(wb_ctrl_csr[0]), .A3(
        wb_ctrl_csr[2]), .Y(n5412) );
  AO21X1_LVT U5427 ( .A1(n9249), .A2(n4515), .A3(n9240), .Y(csr_io_exception)
         );
  AO21X1_LVT U5428 ( .A1(n4514), .A2(n9249), .A3(n3262), .Y(n9240) );
  NBUFFX2_LVT U5429 ( .A(n9525), .Y(n3593) );
  NBUFFX2_LVT U5430 ( .A(clock), .Y(n4499) );
  AND2X1_LVT U5431 ( .A1(n5416), .A2(n5415), .Y(n6859) );
  NBUFFX2_LVT U5432 ( .A(n9526), .Y(n3590) );
  NBUFFX2_LVT U5433 ( .A(n9526), .Y(io_fpu_inst[5]) );
  NOR4X1_LVT U5434 ( .A1(n_T_904[6]), .A2(n_T_904[4]), .A3(n_T_904[7]), .A4(
        n3104), .Y(n9513) );
  NBUFFX2_LVT U5435 ( .A(net34660), .Y(n4073) );
  NBUFFX2_LVT U5436 ( .A(net34660), .Y(n4071) );
  NBUFFX2_LVT U5437 ( .A(net34660), .Y(n4072) );
  NBUFFX2_LVT U5438 ( .A(net34480), .Y(n4294) );
  NBUFFX2_LVT U5439 ( .A(net34480), .Y(n4296) );
  NBUFFX2_LVT U5440 ( .A(net34480), .Y(n4292) );
  NBUFFX2_LVT U5441 ( .A(net34480), .Y(n4293) );
  NBUFFX2_LVT U5442 ( .A(net34480), .Y(n4297) );
  NBUFFX2_LVT U5443 ( .A(net34480), .Y(n4295) );
  NBUFFX2_LVT U5444 ( .A(net34480), .Y(n4299) );
  NBUFFX2_LVT U5445 ( .A(net34469), .Y(n4315) );
  NBUFFX2_LVT U5446 ( .A(net34510), .Y(n4254) );
  NBUFFX2_LVT U5447 ( .A(net34500), .Y(n4266) );
  NBUFFX2_LVT U5448 ( .A(net34515), .Y(n4248) );
  NBUFFX2_LVT U5449 ( .A(net34495), .Y(n4272) );
  NBUFFX2_LVT U5450 ( .A(net34505), .Y(n4260) );
  NBUFFX2_LVT U5451 ( .A(net34490), .Y(n4278) );
  NBUFFX2_LVT U5452 ( .A(net34485), .Y(n4284) );
  NBUFFX2_LVT U5453 ( .A(net34665), .Y(n4070) );
  NBUFFX2_LVT U5454 ( .A(net34665), .Y(n4069) );
  NBUFFX2_LVT U5455 ( .A(net34665), .Y(n4068) );
  NBUFFX2_LVT U5456 ( .A(net34645), .Y(n4091) );
  NBUFFX2_LVT U5457 ( .A(net34570), .Y(n4182) );
  NBUFFX2_LVT U5458 ( .A(net34525), .Y(n4236) );
  NBUFFX2_LVT U5459 ( .A(net34535), .Y(n4224) );
  NBUFFX2_LVT U5460 ( .A(net34635), .Y(n4104) );
  NBUFFX2_LVT U5461 ( .A(net34555), .Y(n4200) );
  NBUFFX2_LVT U5462 ( .A(net34575), .Y(n4176) );
  NBUFFX2_LVT U5463 ( .A(net34565), .Y(n4188) );
  NBUFFX2_LVT U5464 ( .A(net34585), .Y(n4164) );
  NBUFFX2_LVT U5465 ( .A(net34605), .Y(n4140) );
  NBUFFX2_LVT U5466 ( .A(net34545), .Y(n4212) );
  NBUFFX2_LVT U5467 ( .A(net34625), .Y(n4116) );
  NBUFFX2_LVT U5468 ( .A(net34615), .Y(n4128) );
  NBUFFX2_LVT U5469 ( .A(net34595), .Y(n4152) );
  NBUFFX2_LVT U5470 ( .A(net34469), .Y(n4313) );
  NBUFFX2_LVT U5471 ( .A(net34469), .Y(n4314) );
  NBUFFX2_LVT U5472 ( .A(net34469), .Y(n4312) );
  NBUFFX2_LVT U5473 ( .A(net34490), .Y(n4273) );
  NBUFFX2_LVT U5474 ( .A(net34510), .Y(n4249) );
  NBUFFX2_LVT U5475 ( .A(net34495), .Y(n4267) );
  NBUFFX2_LVT U5476 ( .A(net34510), .Y(n4253) );
  NBUFFX2_LVT U5477 ( .A(net34510), .Y(n4252) );
  NBUFFX2_LVT U5478 ( .A(net34510), .Y(n4251) );
  NBUFFX2_LVT U5479 ( .A(net34510), .Y(n4250) );
  NBUFFX2_LVT U5480 ( .A(net34500), .Y(n4261) );
  NBUFFX2_LVT U5481 ( .A(net34490), .Y(n4277) );
  NBUFFX2_LVT U5482 ( .A(net34500), .Y(n4263) );
  NBUFFX2_LVT U5483 ( .A(net34485), .Y(n4281) );
  NBUFFX2_LVT U5484 ( .A(net34505), .Y(n4258) );
  NBUFFX2_LVT U5485 ( .A(net34505), .Y(n4257) );
  NBUFFX2_LVT U5486 ( .A(net34505), .Y(n4256) );
  NBUFFX2_LVT U5487 ( .A(net34515), .Y(n4243) );
  NBUFFX2_LVT U5488 ( .A(net34505), .Y(n4255) );
  NBUFFX2_LVT U5489 ( .A(net34515), .Y(n4244) );
  NBUFFX2_LVT U5490 ( .A(net34500), .Y(n4264) );
  NBUFFX2_LVT U5491 ( .A(net34515), .Y(n4245) );
  NBUFFX2_LVT U5492 ( .A(net34505), .Y(n4259) );
  NBUFFX2_LVT U5493 ( .A(net34515), .Y(n4247) );
  NBUFFX2_LVT U5494 ( .A(net34495), .Y(n4271) );
  NBUFFX2_LVT U5495 ( .A(net34485), .Y(n4279) );
  NBUFFX2_LVT U5496 ( .A(net34500), .Y(n4262) );
  NBUFFX2_LVT U5497 ( .A(net34485), .Y(n4282) );
  NBUFFX2_LVT U5498 ( .A(net34485), .Y(n4283) );
  NBUFFX2_LVT U5499 ( .A(net34500), .Y(n4265) );
  NBUFFX2_LVT U5500 ( .A(net34490), .Y(n4274) );
  NBUFFX2_LVT U5501 ( .A(net34490), .Y(n4276) );
  NBUFFX2_LVT U5502 ( .A(net34495), .Y(n4268) );
  NBUFFX2_LVT U5503 ( .A(net34490), .Y(n4275) );
  NBUFFX2_LVT U5504 ( .A(net34515), .Y(n4246) );
  NBUFFX2_LVT U5505 ( .A(net34495), .Y(n4270) );
  NBUFFX2_LVT U5506 ( .A(net34495), .Y(n4269) );
  NBUFFX2_LVT U5507 ( .A(net34485), .Y(n4280) );
  NBUFFX2_LVT U5508 ( .A(n4285), .Y(n4288) );
  NBUFFX2_LVT U5509 ( .A(n4285), .Y(n4289) );
  NBUFFX2_LVT U5510 ( .A(n4285), .Y(n4290) );
  NBUFFX2_LVT U5511 ( .A(n4285), .Y(n4287) );
  NBUFFX2_LVT U5512 ( .A(n4285), .Y(n4291) );
  NBUFFX2_LVT U5513 ( .A(n4285), .Y(n4298) );
  NBUFFX2_LVT U5514 ( .A(n4285), .Y(n4286) );
  NBUFFX2_LVT U5515 ( .A(net34655), .Y(n4079) );
  NBUFFX2_LVT U5516 ( .A(net34630), .Y(n4110) );
  NBUFFX2_LVT U5517 ( .A(net34590), .Y(n4158) );
  NBUFFX2_LVT U5518 ( .A(net34530), .Y(n4230) );
  NBUFFX2_LVT U5519 ( .A(net34560), .Y(n4194) );
  NBUFFX2_LVT U5520 ( .A(net34600), .Y(n4146) );
  NBUFFX2_LVT U5521 ( .A(net34610), .Y(n4134) );
  NBUFFX2_LVT U5522 ( .A(net34520), .Y(n4242) );
  NBUFFX2_LVT U5523 ( .A(net34540), .Y(n4218) );
  NBUFFX2_LVT U5524 ( .A(net34620), .Y(n4122) );
  NBUFFX2_LVT U5525 ( .A(net34550), .Y(n4206) );
  NBUFFX2_LVT U5526 ( .A(net34580), .Y(n4170) );
  XOR2X1_LVT U5527 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(n592), .Y(n5038) );
  XOR2X1_LVT U5528 ( .A1(n2494), .A2(n588), .Y(n5039) );
  XOR2X1_LVT U5529 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(n591), .Y(n5040) );
  XOR2X1_LVT U5530 ( .A1(n1859), .A2(io_dmem_req_bits_tag[4]), .Y(n5042) );
  XOR2X1_LVT U5531 ( .A1(n2674), .A2(io_dmem_req_bits_tag[3]), .Y(n5043) );
  XOR2X1_LVT U5532 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n3102), .Y(
        n5025) );
  XOR2X1_LVT U5533 ( .A1(n3781), .A2(n3199), .Y(n5026) );
  XOR2X1_LVT U5534 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n3198), .Y(
        n5022) );
  XOR2X1_LVT U5535 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n3103), .Y(
        n5023) );
  XOR2X1_LVT U5536 ( .A1(n2072), .A2(n3201), .Y(n5024) );
  XOR2X1_LVT U5537 ( .A1(n2876), .A2(n5423), .Y(n5000) );
  XOR2X1_LVT U5538 ( .A1(n2825), .A2(n5426), .Y(n5001) );
  XOR2X1_LVT U5539 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n5428), .Y(
        n5002) );
  XOR2X1_LVT U5540 ( .A1(n2098), .A2(n5306), .Y(n5004) );
  XOR2X1_LVT U5541 ( .A1(n2038), .A2(n5313), .Y(n5005) );
  XOR2X1_LVT U5542 ( .A1(n2876), .A2(n3103), .Y(n4937) );
  XOR2X1_LVT U5543 ( .A1(n2825), .A2(n3199), .Y(n4938) );
  XOR2X1_LVT U5544 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n3198), .Y(
        n4939) );
  XOR2X1_LVT U5545 ( .A1(n2038), .A2(n3043), .Y(n4941) );
  XOR2X1_LVT U5546 ( .A1(n2098), .A2(n3041), .Y(n4942) );
  XOR2X1_LVT U5547 ( .A1(n2674), .A2(n3102), .Y(n4920) );
  XOR2X1_LVT U5548 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(n3201), .Y(n4921)
         );
  XOR2X1_LVT U5549 ( .A1(n2494), .A2(n3198), .Y(n4922) );
  XOR2X1_LVT U5550 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(wb_waddr[1]), .Y(
        n4924) );
  XOR2X1_LVT U5551 ( .A1(n1859), .A2(wb_waddr[3]), .Y(n4925) );
  XOR2X1_LVT U5552 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n5423), .Y(
        n4871) );
  XOR2X1_LVT U5553 ( .A1(n3781), .A2(n5426), .Y(n4872) );
  XOR2X1_LVT U5554 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n5428), .Y(
        n4868) );
  XOR2X1_LVT U5555 ( .A1(n2072), .A2(n5427), .Y(n4869) );
  XOR2X1_LVT U5556 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n2575), .Y(
        n4870) );
  XOR2X1_LVT U5557 ( .A1(ibuf_io_inst_0_bits_inst_rd[3]), .A2(n5426), .Y(n4688) );
  XOR2X1_LVT U5558 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n5428), .Y(n4689) );
  XOR2X1_LVT U5559 ( .A1(ibuf_io_inst_0_bits_inst_rd[0]), .A2(n5427), .Y(n4690) );
  XOR2X1_LVT U5560 ( .A1(ibuf_io_inst_0_bits_inst_rd[2]), .A2(n2575), .Y(n4686) );
  XOR2X1_LVT U5561 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n5423), .Y(n4687) );
  XOR2X1_LVT U5562 ( .A1(ibuf_io_inst_0_bits_raw[27]), .A2(n3202), .Y(n4623)
         );
  XOR2X1_LVT U5563 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(n598), .Y(n4625) );
  XOR2X1_LVT U5564 ( .A1(n1859), .A2(n2566), .Y(n4627) );
  XOR2X1_LVT U5565 ( .A1(n2494), .A2(n_T_849[4]), .Y(n4628) );
  XOR2X1_LVT U5566 ( .A1(ibuf_io_inst_0_bits_inst_rd[1]), .A2(n598), .Y(n4622)
         );
  XOR2X1_LVT U5567 ( .A1(n9377), .A2(n_T_698[39]), .Y(n4606) );
  XOR2X1_LVT U5568 ( .A1(n9355), .A2(n124), .Y(n4602) );
  XOR2X1_LVT U5569 ( .A1(n9374), .A2(n104), .Y(n4605) );
  XOR2X1_LVT U5570 ( .A1(n9373), .A2(n_T_698[34]), .Y(n4609) );
  XOR2X1_LVT U5571 ( .A1(n9368), .A2(n_T_698[28]), .Y(n4597) );
  XOR2X1_LVT U5572 ( .A1(n9364), .A2(n_T_698[24]), .Y(n4598) );
  NOR4X1_LVT U5573 ( .A1(n_T_918[39]), .A2(n_T_918[40]), .A3(n_T_918[47]), 
        .A4(n_T_918[60]), .Y(n9464) );
  NOR4X1_LVT U5574 ( .A1(n_T_918[59]), .A2(n_T_918[48]), .A3(n_T_918[62]), 
        .A4(n_T_918[56]), .Y(n9465) );
  NOR4X1_LVT U5575 ( .A1(n_T_918[63]), .A2(n_T_918[46]), .A3(n_T_918[42]), 
        .A4(n_T_918[52]), .Y(n9460) );
  NOR4X1_LVT U5576 ( .A1(n_T_918[41]), .A2(n_T_918[53]), .A3(n_T_918[54]), 
        .A4(n_T_918[50]), .Y(n9461) );
  NOR4X1_LVT U5577 ( .A1(n_T_918[49]), .A2(n_T_918[45]), .A3(n_T_918[61]), 
        .A4(n_T_918[57]), .Y(n9462) );
  NOR4X1_LVT U5578 ( .A1(n_T_918[55]), .A2(n_T_918[58]), .A3(n_T_918[44]), 
        .A4(n_T_918[43]), .Y(n9463) );
  NOR4X1_LVT U5579 ( .A1(n9457), .A2(n9456), .A3(n9455), .A4(n9454), .Y(n9458)
         );
  NBUFFX2_LVT U5580 ( .A(n6830), .Y(n3835) );
  NBUFFX2_LVT U5581 ( .A(n6884), .Y(n3903) );
  NBUFFX2_LVT U5582 ( .A(n6897), .Y(n3956) );
  NBUFFX2_LVT U5583 ( .A(n6895), .Y(n3946) );
  NBUFFX2_LVT U5584 ( .A(n6893), .Y(n3936) );
  NBUFFX2_LVT U5585 ( .A(n6891), .Y(n3926) );
  NBUFFX2_LVT U5586 ( .A(n6812), .Y(n3821) );
  NBUFFX2_LVT U5587 ( .A(n6883), .Y(n3902) );
  NBUFFX2_LVT U5588 ( .A(n6897), .Y(n3955) );
  NBUFFX2_LVT U5589 ( .A(n6895), .Y(n3945) );
  NBUFFX2_LVT U5590 ( .A(n6893), .Y(n3935) );
  NBUFFX2_LVT U5591 ( .A(n6891), .Y(n3925) );
  NBUFFX2_LVT U5592 ( .A(n6882), .Y(n3895) );
  NBUFFX2_LVT U5593 ( .A(n6773), .Y(n3806) );
  NBUFFX2_LVT U5594 ( .A(n6880), .Y(n3893) );
  NBUFFX2_LVT U5595 ( .A(n6795), .Y(n3814) );
  NBUFFX2_LVT U5596 ( .A(n6883), .Y(n3901) );
  NBUFFX2_LVT U5597 ( .A(n6870), .Y(n3873) );
  NBUFFX2_LVT U5598 ( .A(n6829), .Y(n3833) );
  NBUFFX2_LVT U5599 ( .A(n6884), .Y(n3904) );
  NBUFFX2_LVT U5600 ( .A(n6869), .Y(n3870) );
  NBUFFX2_LVT U5601 ( .A(n6812), .Y(n3820) );
  NBUFFX2_LVT U5602 ( .A(n6880), .Y(n3894) );
  NBUFFX2_LVT U5603 ( .A(n6837), .Y(n3838) );
  NBUFFX2_LVT U5604 ( .A(n6811), .Y(n3819) );
  NBUFFX2_LVT U5605 ( .A(n6896), .Y(n3951) );
  NBUFFX2_LVT U5606 ( .A(n6894), .Y(n3941) );
  NBUFFX2_LVT U5607 ( .A(n6892), .Y(n3931) );
  NBUFFX2_LVT U5608 ( .A(n6774), .Y(n3810) );
  NBUFFX2_LVT U5609 ( .A(n6813), .Y(n3823) );
  NBUFFX2_LVT U5610 ( .A(n6884), .Y(n3905) );
  NBUFFX2_LVT U5611 ( .A(n6882), .Y(n3896) );
  NBUFFX2_LVT U5612 ( .A(n6893), .Y(n3933) );
  NBUFFX2_LVT U5613 ( .A(n6774), .Y(n3809) );
  NBUFFX2_LVT U5614 ( .A(n6887), .Y(n3912) );
  NBUFFX2_LVT U5615 ( .A(n6795), .Y(n3813) );
  NBUFFX2_LVT U5616 ( .A(n6868), .Y(n3866) );
  NBUFFX2_LVT U5617 ( .A(n6715), .Y(n3795) );
  NBUFFX2_LVT U5618 ( .A(n6869), .Y(n3869) );
  NBUFFX2_LVT U5619 ( .A(n6882), .Y(n3897) );
  NBUFFX2_LVT U5620 ( .A(n6773), .Y(n3807) );
  NBUFFX2_LVT U5621 ( .A(n6883), .Y(n3899) );
  NBUFFX2_LVT U5622 ( .A(n6897), .Y(n3952) );
  NBUFFX2_LVT U5623 ( .A(n6895), .Y(n3942) );
  NBUFFX2_LVT U5624 ( .A(n6891), .Y(n3922) );
  NBUFFX2_LVT U5625 ( .A(n6880), .Y(n3890) );
  NBUFFX2_LVT U5626 ( .A(n6888), .Y(n3913) );
  NBUFFX2_LVT U5627 ( .A(n6887), .Y(n3911) );
  NBUFFX2_LVT U5628 ( .A(n6773), .Y(n3808) );
  OR2X1_LVT U5629 ( .A1(n8803), .A2(n2645), .Y(n8804) );
  NBUFFX2_LVT U5630 ( .A(n_T_427__T_1136_data[57]), .Y(n4478) );
  NBUFFX2_LVT U5631 ( .A(n6715), .Y(n3797) );
  NBUFFX2_LVT U5632 ( .A(n6837), .Y(n3837) );
  NBUFFX2_LVT U5633 ( .A(n6813), .Y(n3822) );
  NBUFFX2_LVT U5634 ( .A(n6890), .Y(n3917) );
  NBUFFX2_LVT U5635 ( .A(n6891), .Y(n3923) );
  NBUFFX2_LVT U5636 ( .A(n6893), .Y(n3932) );
  NBUFFX2_LVT U5637 ( .A(n6880), .Y(n3891) );
  NBUFFX2_LVT U5638 ( .A(n6879), .Y(n3885) );
  NBUFFX2_LVT U5639 ( .A(n6829), .Y(n3831) );
  NBUFFX2_LVT U5640 ( .A(n6896), .Y(n3947) );
  NBUFFX2_LVT U5641 ( .A(n6897), .Y(n3953) );
  NBUFFX2_LVT U5642 ( .A(n6883), .Y(n3898) );
  NBUFFX2_LVT U5643 ( .A(n6895), .Y(n3943) );
  NBUFFX2_LVT U5644 ( .A(n6894), .Y(n3937) );
  NBUFFX2_LVT U5645 ( .A(n_T_427__T_1136_data[51]), .Y(n4460) );
  NBUFFX2_LVT U5646 ( .A(n_T_427__T_1136_data[53]), .Y(n4466) );
  NBUFFX2_LVT U5647 ( .A(n_T_427__T_1136_data[54]), .Y(n4469) );
  NBUFFX2_LVT U5648 ( .A(n_T_427__T_1136_data[60]), .Y(n4487) );
  OR2X1_LVT U5649 ( .A1(n8878), .A2(n2155), .Y(n8879) );
  NBUFFX2_LVT U5650 ( .A(n_T_427__T_1136_data[59]), .Y(n4484) );
  NBUFFX2_LVT U5651 ( .A(n_T_427__T_1136_data[45]), .Y(n4442) );
  NBUFFX2_LVT U5652 ( .A(n_T_427__T_1136_data[16]), .Y(n4364) );
  NBUFFX2_LVT U5653 ( .A(n_T_427__T_1136_data[24]), .Y(n4386) );
  NAND3X0_LVT U5654 ( .A1(n3731), .A2(n3732), .A3(n3733), .Y(N738) );
  NBUFFX2_LVT U5655 ( .A(n_T_427__T_1136_data[58]), .Y(n4481) );
  NBUFFX2_LVT U5656 ( .A(n_T_427__T_1136_data[47]), .Y(n4448) );
  OA21X1_LVT U5657 ( .A1(n3477), .A2(n3753), .A3(n8442), .Y(n8445) );
  NBUFFX2_LVT U5658 ( .A(n_T_427__T_1136_data[49]), .Y(n4454) );
  NBUFFX2_LVT U5659 ( .A(n6829), .Y(n3832) );
  NBUFFX2_LVT U5660 ( .A(n6883), .Y(n3900) );
  NBUFFX2_LVT U5661 ( .A(n6896), .Y(n3949) );
  AND2X1_LVT U5662 ( .A1(n5457), .A2(n5455), .Y(n6896) );
  NBUFFX2_LVT U5663 ( .A(n6897), .Y(n3954) );
  NBUFFX2_LVT U5664 ( .A(n6894), .Y(n3939) );
  AND2X1_LVT U5665 ( .A1(n5457), .A2(n2034), .Y(n6894) );
  NBUFFX2_LVT U5666 ( .A(n6895), .Y(n3944) );
  NBUFFX2_LVT U5667 ( .A(n6892), .Y(n3929) );
  AND2X1_LVT U5668 ( .A1(n5457), .A2(n5451), .Y(n6892) );
  NBUFFX2_LVT U5669 ( .A(n6893), .Y(n3934) );
  NBUFFX2_LVT U5670 ( .A(n6890), .Y(n3919) );
  AND2X1_LVT U5671 ( .A1(n5457), .A2(n5449), .Y(n6890) );
  NBUFFX2_LVT U5672 ( .A(n6891), .Y(n3924) );
  NBUFFX2_LVT U5673 ( .A(n6879), .Y(n3886) );
  AND2X1_LVT U5674 ( .A1(n5446), .A2(n5454), .Y(n6879) );
  NBUFFX2_LVT U5675 ( .A(n6880), .Y(n3892) );
  AND2X1_LVT U5676 ( .A1(n5437), .A2(n5449), .Y(n3579) );
  NBUFFX2_LVT U5677 ( .A(n6870), .Y(n3872) );
  NBUFFX2_LVT U5678 ( .A(n6865), .Y(n3860) );
  NBUFFX2_LVT U5679 ( .A(n6889), .Y(n3915) );
  NBUFFX2_LVT U5680 ( .A(n6811), .Y(n3818) );
  NBUFFX2_LVT U5681 ( .A(n6887), .Y(n3910) );
  NBUFFX2_LVT U5682 ( .A(n6830), .Y(n3834) );
  XOR2X1_LVT U5683 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n592), .Y(n4861) );
  XOR2X1_LVT U5684 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n588), .Y(n4862) );
  XOR2X1_LVT U5685 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n590), .Y(n4863) );
  XOR2X1_LVT U5686 ( .A1(n3781), .A2(n589), .Y(n4864) );
  XOR2X1_LVT U5687 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n591), .Y(n5044) );
  XOR2X1_LVT U5688 ( .A1(ibuf_io_inst_0_bits_inst_rs2[2]), .A2(n3200), .Y(
        n4629) );
  XOR2X1_LVT U5689 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n598), .Y(n4630) );
  XOR2X1_LVT U5690 ( .A1(ibuf_io_inst_0_bits_inst_rs2[4]), .A2(n595), .Y(n4631) );
  XOR2X1_LVT U5691 ( .A1(n3781), .A2(n596), .Y(n4632) );
  XOR2X1_LVT U5692 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n_T_849[11]), 
        .Y(n4860) );
  NBUFFX2_LVT U5693 ( .A(n_T_427__T_1136_data[55]), .Y(n4472) );
  NBUFFX2_LVT U5694 ( .A(n_T_427__T_1136_data[32]), .Y(n4406) );
  NBUFFX2_LVT U5695 ( .A(n_T_427__T_1136_data[50]), .Y(n4457) );
  NBUFFX2_LVT U5696 ( .A(n_T_427__T_1136_data[40]), .Y(n4427) );
  NBUFFX2_LVT U5697 ( .A(n_T_427__T_1136_data[1]), .Y(n4321) );
  NBUFFX2_LVT U5698 ( .A(n_T_427__T_1136_data[43]), .Y(n4436) );
  NAND3X0_LVT U5699 ( .A1(n3735), .A2(n3736), .A3(n3737), .Y(N732) );
  OR2X1_LVT U5700 ( .A1(n8624), .A2(n3656), .Y(n8625) );
  NBUFFX2_LVT U5701 ( .A(n_T_427__T_1136_data[52]), .Y(n4463) );
  NAND3X0_LVT U5702 ( .A1(n3748), .A2(n3749), .A3(n3750), .Y(N743) );
  OR2X1_LVT U5703 ( .A1(n9048), .A2(n3632), .Y(n9049) );
  NBUFFX2_LVT U5704 ( .A(n_T_427__T_1136_data[63]), .Y(n4496) );
  NBUFFX2_LVT U5705 ( .A(n_T_427__T_1136_data[19]), .Y(n4373) );
  NBUFFX2_LVT U5706 ( .A(n_T_427__T_1136_data[56]), .Y(n4475) );
  NBUFFX2_LVT U5707 ( .A(n_T_427__T_1136_data[44]), .Y(n4439) );
  NBUFFX2_LVT U5708 ( .A(n_T_427__T_1136_data[37]), .Y(n4419) );
  NBUFFX2_LVT U5709 ( .A(n_T_427__T_1136_data[48]), .Y(n4451) );
  NBUFFX2_LVT U5710 ( .A(n8932), .Y(n3975) );
  OR2X1_LVT U5711 ( .A1(n8987), .A2(n2155), .Y(n8988) );
  NBUFFX2_LVT U5712 ( .A(n_T_427__T_1136_data[62]), .Y(n4493) );
  NBUFFX2_LVT U5713 ( .A(n_T_427__T_1136_data[41]), .Y(n4430) );
  OA21X1_LVT U5714 ( .A1(n3475), .A2(n3601), .A3(n8246), .Y(n8249) );
  NBUFFX2_LVT U5715 ( .A(n3182), .Y(n4048) );
  NBUFFX2_LVT U5716 ( .A(n_T_427__T_1136_data[39]), .Y(n4424) );
  NBUFFX2_LVT U5717 ( .A(n_T_427__T_1136_data[36]), .Y(n4416) );
  NBUFFX2_LVT U5718 ( .A(n8901), .Y(n3967) );
  NBUFFX2_LVT U5719 ( .A(n_T_427__T_1136_data[46]), .Y(n4445) );
  NBUFFX2_LVT U5720 ( .A(n6858), .Y(n3845) );
  NBUFFX2_LVT U5721 ( .A(n9037), .Y(n4021) );
  NBUFFX2_LVT U5722 ( .A(n9041), .Y(n4044) );
  NBUFFX2_LVT U5723 ( .A(n8982), .Y(n3986) );
  NBUFFX2_LVT U5724 ( .A(n_T_427__T_1136_data[34]), .Y(n4411) );
  AND2X1_LVT U5725 ( .A1(n3712), .A2(n_T_427[993]), .Y(n3763) );
  NBUFFX2_LVT U5726 ( .A(n9029), .Y(n3641) );
  NBUFFX2_LVT U5727 ( .A(n_T_427__T_1136_data[61]), .Y(n4490) );
  NBUFFX2_LVT U5728 ( .A(n9016), .Y(n4001) );
  NBUFFX2_LVT U5729 ( .A(n_T_427__T_1136_data[17]), .Y(n4367) );
  NBUFFX2_LVT U5730 ( .A(n_T_427__T_1136_data[20]), .Y(n4376) );
  NBUFFX2_LVT U5731 ( .A(n9042), .Y(n4052) );
  NBUFFX2_LVT U5732 ( .A(n8931), .Y(n3971) );
  NBUFFX2_LVT U5733 ( .A(n9037), .Y(n4022) );
  NBUFFX2_LVT U5734 ( .A(n9039), .Y(n4035) );
  NBUFFX2_LVT U5735 ( .A(n_T_427__T_1136_data[42]), .Y(n4433) );
  NBUFFX2_LVT U5736 ( .A(n9016), .Y(n4002) );
  INVX1_LVT U5737 ( .A(n9014), .Y(n3995) );
  NBUFFX2_LVT U5738 ( .A(n9039), .Y(n4031) );
  NBUFFX2_LVT U5739 ( .A(n8900), .Y(n3961) );
  NBUFFX2_LVT U5740 ( .A(n8981), .Y(n3980) );
  INVX1_LVT U5741 ( .A(n9006), .Y(n3990) );
  NBUFFX2_LVT U5742 ( .A(n9015), .Y(n4000) );
  NBUFFX2_LVT U5743 ( .A(n_T_427__T_1136_data[0]), .Y(n4318) );
  NBUFFX2_LVT U5744 ( .A(n6858), .Y(n3841) );
  NBUFFX2_LVT U5745 ( .A(n9041), .Y(n4041) );
  NBUFFX2_LVT U5746 ( .A(n3182), .Y(n4045) );
  NBUFFX2_LVT U5747 ( .A(n9039), .Y(n4032) );
  NBUFFX2_LVT U5748 ( .A(n9038), .Y(n4030) );
  NBUFFX2_LVT U5749 ( .A(n9037), .Y(n4018) );
  NBUFFX2_LVT U5750 ( .A(n9042), .Y(n4049) );
  NBUFFX2_LVT U5751 ( .A(n_T_427__T_1136_data[30]), .Y(n4401) );
  NBUFFX2_LVT U5752 ( .A(n8900), .Y(n3963) );
  NBUFFX2_LVT U5753 ( .A(n8981), .Y(n3982) );
  NBUFFX2_LVT U5754 ( .A(n6859), .Y(n3848) );
  NBUFFX2_LVT U5755 ( .A(n_T_427__T_1136_data[27]), .Y(n4393) );
  NBUFFX2_LVT U5756 ( .A(n_T_427__T_1136_data[23]), .Y(n4383) );
  NBUFFX2_LVT U5757 ( .A(n6861), .Y(n3858) );
  NBUFFX2_LVT U5758 ( .A(n6858), .Y(n3844) );
  NBUFFX2_LVT U5759 ( .A(n9041), .Y(n4043) );
  NBUFFX2_LVT U5760 ( .A(n3182), .Y(n4047) );
  NBUFFX2_LVT U5761 ( .A(n8932), .Y(n3974) );
  NBUFFX2_LVT U5762 ( .A(n8901), .Y(n3966) );
  NBUFFX2_LVT U5763 ( .A(n8931), .Y(n3970) );
  NBUFFX2_LVT U5764 ( .A(n8982), .Y(n3985) );
  NBUFFX2_LVT U5765 ( .A(n9039), .Y(n4034) );
  NBUFFX2_LVT U5766 ( .A(n9038), .Y(n4028) );
  NBUFFX2_LVT U5767 ( .A(n9037), .Y(n4020) );
  NBUFFX2_LVT U5768 ( .A(n_T_427__T_1136_data[29]), .Y(n4398) );
  NBUFFX2_LVT U5769 ( .A(n6860), .Y(n3851) );
  NBUFFX2_LVT U5770 ( .A(n9016), .Y(n4003) );
  NBUFFX2_LVT U5771 ( .A(n9015), .Y(n3998) );
  NBUFFX2_LVT U5772 ( .A(n9041), .Y(n4042) );
  NBUFFX2_LVT U5773 ( .A(n8900), .Y(n3962) );
  NBUFFX2_LVT U5774 ( .A(n3182), .Y(n4046) );
  NBUFFX2_LVT U5775 ( .A(n8981), .Y(n3981) );
  NBUFFX2_LVT U5776 ( .A(n8932), .Y(n3973) );
  NBUFFX2_LVT U5777 ( .A(n8901), .Y(n3965) );
  NBUFFX2_LVT U5778 ( .A(n8931), .Y(n3969) );
  NBUFFX2_LVT U5779 ( .A(n8982), .Y(n3984) );
  NBUFFX2_LVT U5780 ( .A(n9039), .Y(n4033) );
  NBUFFX2_LVT U5781 ( .A(n9038), .Y(n4029) );
  NBUFFX2_LVT U5782 ( .A(n8980), .Y(n3977) );
  NBUFFX2_LVT U5783 ( .A(n9037), .Y(n4019) );
  NBUFFX2_LVT U5784 ( .A(n9042), .Y(n4050) );
  NBUFFX2_LVT U5785 ( .A(n_T_427__T_1136_data[18]), .Y(n4370) );
  NBUFFX2_LVT U5786 ( .A(n6859), .Y(n3849) );
  NBUFFX2_LVT U5787 ( .A(n6858), .Y(n3843) );
  INVX1_LVT U5788 ( .A(n9008), .Y(n3993) );
  XOR2X1_LVT U5789 ( .A1(io_fpu_inst[20]), .A2(n9522), .Y(n5142) );
  INVX1_LVT U5790 ( .A(n5394), .Y(n3567) );
  OA21X1_LVT U5791 ( .A1(n5118), .A2(n3039), .A3(n5111), .Y(n5112) );
  XOR2X1_LVT U5792 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n592), .Y(n5011) );
  XOR2X1_LVT U5793 ( .A1(n2876), .A2(n598), .Y(n4615) );
  XOR2X1_LVT U5794 ( .A1(ibuf_io_inst_0_bits_inst_rs1[2]), .A2(n3200), .Y(
        n4616) );
  OA21X1_LVT U5795 ( .A1(io_fpu_inst[2]), .A2(n3076), .A3(n5165), .Y(n5109) );
  NBUFFX2_LVT U5796 ( .A(n6888), .Y(n3914) );
  NBUFFX2_LVT U5797 ( .A(n6885), .Y(n3907) );
  NBUFFX2_LVT U5798 ( .A(n6885), .Y(n3906) );
  NBUFFX2_LVT U5799 ( .A(n6838), .Y(n3839) );
  AND3X1_LVT U5800 ( .A1(n6118), .A2(n6117), .A3(n6116), .Y(n3091) );
  NAND2X0_LVT U5801 ( .A1(wb_cause[3]), .A2(n9252), .Y(n3100) );
  NBUFFX2_LVT U5802 ( .A(n9015), .Y(n3997) );
  NBUFFX2_LVT U5803 ( .A(n9015), .Y(n3996) );
  NBUFFX2_LVT U5804 ( .A(n9015), .Y(n3999) );
  NBUFFX2_LVT U5805 ( .A(n9016), .Y(n4004) );
  NBUFFX2_LVT U5806 ( .A(n9016), .Y(n4005) );
  NBUFFX2_LVT U5807 ( .A(n6886), .Y(n3909) );
  NBUFFX2_LVT U5808 ( .A(n6889), .Y(n3916) );
  AND4X1_LVT U5809 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .Y(n3181)
         );
  NBUFFX2_LVT U5810 ( .A(n6796), .Y(n3816) );
  NBUFFX2_LVT U5811 ( .A(n6796), .Y(n3815) );
  NBUFFX2_LVT U5812 ( .A(n6898), .Y(n3959) );
  NBUFFX2_LVT U5813 ( .A(n6892), .Y(n3927) );
  NBUFFX2_LVT U5814 ( .A(n6892), .Y(n3930) );
  NBUFFX2_LVT U5815 ( .A(n6892), .Y(n3928) );
  NBUFFX2_LVT U5816 ( .A(n6890), .Y(n3920) );
  NBUFFX2_LVT U5817 ( .A(n6890), .Y(n3918) );
  NBUFFX2_LVT U5818 ( .A(n6890), .Y(n3921) );
  NBUFFX2_LVT U5819 ( .A(n6894), .Y(n3938) );
  NBUFFX2_LVT U5820 ( .A(n6894), .Y(n3940) );
  NBUFFX2_LVT U5821 ( .A(n6896), .Y(n3948) );
  NBUFFX2_LVT U5822 ( .A(n6896), .Y(n3950) );
  NBUFFX2_LVT U5823 ( .A(n6879), .Y(n3889) );
  NBUFFX2_LVT U5824 ( .A(n6879), .Y(n3888) );
  NBUFFX2_LVT U5825 ( .A(n6879), .Y(n3887) );
  NBUFFX2_LVT U5826 ( .A(n8980), .Y(n3978) );
  AND3X1_LVT U5827 ( .A1(n6166), .A2(n6165), .A3(n6164), .Y(n3183) );
  NAND2X0_LVT U5828 ( .A1(n6946), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n3184) );
  NBUFFX2_LVT U5829 ( .A(n6810), .Y(n3817) );
  NBUFFX2_LVT U5830 ( .A(n6859), .Y(n3850) );
  NBUFFX2_LVT U5831 ( .A(n6858), .Y(n3842) );
  NBUFFX2_LVT U5832 ( .A(n9101), .Y(n4054) );
  AND4X1_LVT U5833 ( .A1(n9481), .A2(n9480), .A3(n9479), .A4(n9478), .Y(n3204)
         );
  AND2X1_LVT U5834 ( .A1(n3078), .A2(n9105), .Y(n3566) );
  OA22X1_LVT U5835 ( .A1(n5115), .A2(n3571), .A3(n3570), .A4(n1699), .Y(n3576)
         );
  OR2X1_LVT U5836 ( .A1(csr_io_status_isa[3]), .A2(n3039), .Y(n3571) );
  AND4X1_LVT U5837 ( .A1(n3576), .A2(n5112), .A3(n5121), .A4(n5120), .Y(n3572)
         );
  AND2X1_LVT U5838 ( .A1(n3574), .A2(n5113), .Y(n3573) );
  NAND2X0_LVT U5839 ( .A1(n9231), .A2(n3575), .Y(n9413) );
  AO22X1_LVT U5840 ( .A1(n1853), .A2(n3577), .A3(n1867), .A4(n1891), .Y(
        id_ctrl_sel_imm[0]) );
  NAND4X0_LVT U5841 ( .A1(n4616), .A2(n4615), .A3(n4617), .A4(n3581), .Y(n4847) );
  NAND2X0_LVT U5842 ( .A1(n5446), .A2(n5450), .Y(n6878) );
  AND2X1_LVT U5843 ( .A1(n9446), .A2(io_fpu_inst[12]), .Y(n9230) );
  AND2X1_LVT U5844 ( .A1(n9446), .A2(n3077), .Y(n5101) );
  NAND2X0_LVT U5845 ( .A1(n3583), .A2(io_fpu_inst[14]), .Y(n5105) );
  NAND2X0_LVT U5846 ( .A1(n2547), .A2(n2131), .Y(n5122) );
  NAND2X0_LVT U5847 ( .A1(n5077), .A2(n5076), .Y(n3584) );
  AND2X1_LVT U5848 ( .A1(n9440), .A2(io_fpu_inst[28]), .Y(n3585) );
  OA22X1_LVT U5849 ( .A1(n5443), .A2(n3586), .A3(n3490), .A4(n3880), .Y(n5445)
         );
  OA22X1_LVT U5850 ( .A1(n6695), .A2(n3586), .A3(n3491), .A4(n3882), .Y(n6698)
         );
  OA22X1_LVT U5851 ( .A1(n6720), .A2(n3586), .A3(n3492), .A4(n3882), .Y(n6723)
         );
  OA22X1_LVT U5852 ( .A1(n6739), .A2(n3586), .A3(n3493), .A4(n3882), .Y(n6743)
         );
  OA22X1_LVT U5853 ( .A1(n6801), .A2(n3586), .A3(n3483), .A4(n3882), .Y(n6805)
         );
  OA22X1_LVT U5854 ( .A1(n6843), .A2(n3586), .A3(n3484), .A4(n3882), .Y(n6846)
         );
  NBUFFX2_LVT U5855 ( .A(net34650), .Y(n4085) );
  NAND2X0_LVT U5856 ( .A1(n9253), .A2(csr_io_exception), .Y(n9254) );
  AND2X1_LVT U5857 ( .A1(n3100), .A2(n3589), .Y(n9253) );
  INVX1_LVT U5858 ( .A(wb_cause[63]), .Y(n3589) );
  AND3X1_LVT U5918 ( .A1(n7138), .A2(n7137), .A3(n7136), .Y(n3598) );
  AND3X1_LVT U5919 ( .A1(n7131), .A2(n7130), .A3(n7129), .Y(n3599) );
  NBUFFX2_LVT U5920 ( .A(n9053), .Y(n3789) );
  NBUFFX2_LVT U5921 ( .A(n3613), .Y(n3602) );
  NBUFFX2_LVT U5922 ( .A(n9004), .Y(n3603) );
  NBUFFX2_LVT U5923 ( .A(n9004), .Y(n3604) );
  NBUFFX2_LVT U5924 ( .A(n9004), .Y(n3605) );
  NBUFFX2_LVT U5925 ( .A(n3613), .Y(n3606) );
  NBUFFX2_LVT U5926 ( .A(n9004), .Y(n3607) );
  NBUFFX2_LVT U5927 ( .A(n3613), .Y(n3608) );
  NBUFFX2_LVT U5928 ( .A(n3613), .Y(n3609) );
  NBUFFX2_LVT U5929 ( .A(n9004), .Y(n3611) );
  NBUFFX2_LVT U5930 ( .A(n9047), .Y(n3612) );
  NBUFFX2_LVT U5931 ( .A(n9021), .Y(n3615) );
  NBUFFX2_LVT U5932 ( .A(n9021), .Y(n3616) );
  NBUFFX2_LVT U5933 ( .A(n9021), .Y(n3617) );
  NBUFFX2_LVT U5934 ( .A(n9021), .Y(n3618) );
  NBUFFX2_LVT U5935 ( .A(n9021), .Y(n3619) );
  NBUFFX2_LVT U5936 ( .A(n9021), .Y(n3620) );
  NBUFFX2_LVT U5937 ( .A(n9021), .Y(n3621) );
  AND3X1_LVT U5938 ( .A1(n8006), .A2(n8007), .A3(n8008), .Y(n3622) );
  AND3X1_LVT U5939 ( .A1(n8005), .A2(n8004), .A3(n8003), .Y(n3623) );
  NBUFFX2_LVT U5940 ( .A(n9058), .Y(n3624) );
  NBUFFX2_LVT U5941 ( .A(n9007), .Y(n3626) );
  NBUFFX2_LVT U5942 ( .A(n9007), .Y(n3627) );
  NBUFFX2_LVT U5943 ( .A(n9007), .Y(n3628) );
  NBUFFX2_LVT U5944 ( .A(n9007), .Y(n3629) );
  NBUFFX2_LVT U5945 ( .A(n9007), .Y(n3630) );
  AND3X1_LVT U5946 ( .A1(n8942), .A2(n8941), .A3(n8940), .Y(n3634) );
  NBUFFX2_LVT U5947 ( .A(n9029), .Y(n3635) );
  NBUFFX2_LVT U5948 ( .A(n9029), .Y(n3636) );
  NBUFFX2_LVT U5949 ( .A(n9029), .Y(n3638) );
  NBUFFX2_LVT U5950 ( .A(n9029), .Y(n3639) );
  NBUFFX2_LVT U5951 ( .A(n9029), .Y(n3640) );
  OR2X1_LVT U5952 ( .A1(n4016), .A2(n3644), .Y(n8753) );
  OR2X1_LVT U5953 ( .A1(n2090), .A2(n3645), .Y(n7874) );
  OR2X1_LVT U5954 ( .A1(n9412), .A2(n3646), .Y(n6971) );
  NBUFFX2_LVT U5955 ( .A(n8944), .Y(n3647) );
  NBUFFX2_LVT U5956 ( .A(n9022), .Y(n3648) );
  NBUFFX2_LVT U5957 ( .A(n9022), .Y(n3650) );
  NBUFFX2_LVT U5958 ( .A(n9022), .Y(n3651) );
  NBUFFX2_LVT U5959 ( .A(n9022), .Y(n3652) );
  OR2X1_LVT U5960 ( .A1(n2069), .A2(n3655), .Y(n7966) );
  NBUFFX2_LVT U5961 ( .A(n9012), .Y(n3657) );
  OR2X1_LVT U5962 ( .A1(n2089), .A2(n3659), .Y(n8389) );
  OR2X1_LVT U5963 ( .A1(n2090), .A2(n3660), .Y(n8426) );
  OR2X1_LVT U5964 ( .A1(n4016), .A2(n3090), .Y(n7814) );
  AND3X1_LVT U5965 ( .A1(n8725), .A2(n8724), .A3(n8723), .Y(n3662) );
  NBUFFX2_LVT U5966 ( .A(n9030), .Y(n3668) );
  NBUFFX2_LVT U5967 ( .A(n9030), .Y(n3669) );
  NBUFFX2_LVT U5968 ( .A(n3666), .Y(n3670) );
  NBUFFX2_LVT U5969 ( .A(n3666), .Y(n3671) );
  NBUFFX2_LVT U5970 ( .A(n3666), .Y(n3672) );
  NBUFFX2_LVT U5971 ( .A(n9030), .Y(n3673) );
  NBUFFX2_LVT U5972 ( .A(n9030), .Y(n3674) );
  NBUFFX2_LVT U5973 ( .A(n9030), .Y(n3675) );
  AND3X1_LVT U5974 ( .A1(n8037), .A2(n8036), .A3(n8038), .Y(n3676) );
  AND3X1_LVT U5975 ( .A1(n8041), .A2(n8040), .A3(n8039), .Y(n3677) );
  AND3X1_LVT U5976 ( .A1(n8736), .A2(n8735), .A3(n8737), .Y(n3678) );
  OR2X1_LVT U5977 ( .A1(n4016), .A2(n3679), .Y(n6943) );
  AND3X1_LVT U5978 ( .A1(n7532), .A2(n7531), .A3(n7530), .Y(n3680) );
  AND3X1_LVT U5979 ( .A1(n7515), .A2(n7514), .A3(n7513), .Y(n3681) );
  AND3X1_LVT U5980 ( .A1(n7517), .A2(n7518), .A3(n7519), .Y(n3682) );
  OR2X1_LVT U5981 ( .A1(n2069), .A2(n3685), .Y(n8131) );
  OA21X1_LVT U5982 ( .A1(n3412), .A2(n3753), .A3(n8591), .Y(n8594) );
  OA21X1_LVT U5983 ( .A1(n3413), .A2(n3751), .A3(n8374), .Y(n8377) );
  OR2X1_LVT U5984 ( .A1(n2090), .A2(n3686), .Y(n6997) );
  OR2X1_LVT U5985 ( .A1(n2089), .A2(n3687), .Y(n8072) );
  OR2X1_LVT U5986 ( .A1(n2090), .A2(n3688), .Y(n8321) );
  OA21X1_LVT U5987 ( .A1(n3414), .A2(n3753), .A3(n8488), .Y(n8491) );
  OA21X1_LVT U5988 ( .A1(n3415), .A2(n3753), .A3(n8358), .Y(n8361) );
  AND3X1_LVT U5989 ( .A1(n8024), .A2(n8025), .A3(n8026), .Y(n3690) );
  NBUFFX2_LVT U5990 ( .A(n3708), .Y(n3691) );
  AND3X1_LVT U5991 ( .A1(n7705), .A2(n7704), .A3(n7703), .Y(n3693) );
  AND3X1_LVT U5992 ( .A1(n7701), .A2(n7700), .A3(n7699), .Y(n3694) );
  AND3X1_LVT U5993 ( .A1(n7718), .A2(n7717), .A3(n7716), .Y(n3695) );
  AND3X1_LVT U5994 ( .A1(n7454), .A2(n7453), .A3(n7452), .Y(n3696) );
  AND3X1_LVT U5995 ( .A1(n7470), .A2(n7469), .A3(n7468), .Y(n3697) );
  AND3X1_LVT U5996 ( .A1(n7738), .A2(n7737), .A3(n7736), .Y(n3698) );
  AND3X1_LVT U5997 ( .A1(n7734), .A2(n7733), .A3(n7732), .Y(n3699) );
  AND3X1_LVT U5998 ( .A1(n7751), .A2(n7750), .A3(n7749), .Y(n3700) );
  AND3X1_LVT U5999 ( .A1(n7607), .A2(n7606), .A3(n7605), .Y(n3701) );
  AND3X1_LVT U6000 ( .A1(n7622), .A2(n7621), .A3(n7620), .Y(n3702) );
  AND3X1_LVT U6001 ( .A1(n7544), .A2(n7543), .A3(n7542), .Y(n3703) );
  AND3X1_LVT U6002 ( .A1(n7559), .A2(n7558), .A3(n7557), .Y(n3704) );
  AND3X1_LVT U6003 ( .A1(n7575), .A2(n7574), .A3(n7573), .Y(n3705) );
  AND3X1_LVT U6004 ( .A1(n7591), .A2(n7590), .A3(n7589), .Y(n3706) );
  NBUFFX2_LVT U6005 ( .A(n8994), .Y(n3707) );
  NAND2X0_LVT U6006 ( .A1(n3182), .A2(n8105), .Y(n3708) );
  OR2X1_LVT U6007 ( .A1(n4016), .A2(n3710), .Y(n7441) );
  OR2X1_LVT U6008 ( .A1(n4016), .A2(n3711), .Y(n7847) );
  NBUFFX2_LVT U6009 ( .A(n9059), .Y(n3713) );
  NBUFFX2_LVT U6010 ( .A(n9059), .Y(n3714) );
  NBUFFX2_LVT U6011 ( .A(n9059), .Y(n3791) );
  AND3X1_LVT U6012 ( .A1(n8696), .A2(n8695), .A3(n8694), .Y(n3718) );
  AND3X1_LVT U6013 ( .A1(n8692), .A2(n8691), .A3(n8690), .Y(n3720) );
  AND3X1_LVT U6014 ( .A1(n8660), .A2(n8659), .A3(n8658), .Y(n3721) );
  AND3X1_LVT U6015 ( .A1(n8654), .A2(n8653), .A3(n8652), .Y(n3722) );
  AND2X1_LVT U6016 ( .A1(n8910), .A2(n8909), .Y(n3723) );
  AND3X1_LVT U6017 ( .A1(n8908), .A2(n8907), .A3(n8906), .Y(n3724) );
  AND2X1_LVT U6018 ( .A1(n8588), .A2(n8587), .Y(n3726) );
  AND3X1_LVT U6019 ( .A1(n8586), .A2(n8585), .A3(n8584), .Y(n3727) );
  NAND3X0_LVT U6020 ( .A1(n3728), .A2(n3729), .A3(n3730), .Y(N739) );
  NOR3X0_LVT U6021 ( .A1(n8849), .A2(n8850), .A3(n8851), .Y(n3733) );
  NOR3X0_LVT U6022 ( .A1(n8813), .A2(n8814), .A3(n8815), .Y(n3734) );
  NAND3X0_LVT U6023 ( .A1(n3738), .A2(n3739), .A3(n3740), .Y(N729) );
  NAND3X0_LVT U6024 ( .A1(n3741), .A2(n3742), .A3(n3743), .Y(N727) );
  NBUFFX2_LVT U6025 ( .A(n9058), .Y(n3745) );
  XOR2X1_LVT U6026 ( .A1(n2876), .A2(n9390), .Y(n6907) );
  NBUFFX2_LVT U6027 ( .A(n9014), .Y(n3751) );
  NBUFFX2_LVT U6028 ( .A(n9028), .Y(n3752) );
  NBUFFX2_LVT U6029 ( .A(n9014), .Y(n3753) );
  AND3X1_LVT U6030 ( .A1(n8241), .A2(n8240), .A3(n8239), .Y(n3754) );
  NBUFFX2_LVT U6031 ( .A(n9026), .Y(n3755) );
  AND3X1_LVT U6032 ( .A1(n7993), .A2(n7992), .A3(n7991), .Y(n3762) );
  AOI21X1_LVT U6033 ( .A1(n3716), .A2(n_T_427[1057]), .A3(n3763), .Y(n8008) );
  INVX1_LVT U6034 ( .A(n9006), .Y(n3764) );
  AND2X1_LVT U6035 ( .A1(n6962), .A2(n6965), .Y(n3765) );
  AND3X1_LVT U6036 ( .A1(n7989), .A2(n7988), .A3(n7987), .Y(n3766) );
  NBUFFX2_LVT U6037 ( .A(n9006), .Y(n3767) );
  OR2X1_LVT U6038 ( .A1(n3653), .A2(n3774), .Y(n8492) );
  AOI21X1_LVT U6039 ( .A1(n4014), .A2(n_T_427[1058]), .A3(n3775), .Y(n8041) );
  AND2X1_LVT U6040 ( .A1(n3712), .A2(n_T_427[994]), .Y(n3775) );
  AND2X1_LVT U6041 ( .A1(n3712), .A2(n_T_427[1014]), .Y(n3776) );
  AND2X1_LVT U6042 ( .A1(n3712), .A2(n_T_427[1000]), .Y(n3777) );
  AND3X1_LVT U6043 ( .A1(n8237), .A2(n8236), .A3(n8235), .Y(n3778) );
  AND3X1_LVT U6044 ( .A1(n8022), .A2(n8021), .A3(n8020), .Y(n3779) );
  AND3X1_LVT U6045 ( .A1(n8720), .A2(n8719), .A3(n8718), .Y(n3780) );
  NBUFFX2_LVT U6046 ( .A(n9035), .Y(n3786) );
  NBUFFX2_LVT U6047 ( .A(n9035), .Y(n3787) );
  NBUFFX2_LVT U6048 ( .A(n9035), .Y(n3788) );
  NBUFFX2_LVT U6049 ( .A(n9053), .Y(n3790) );
  NBUFFX2_LVT U6050 ( .A(net34475), .Y(n4300) );
  NBUFFX2_LVT U6051 ( .A(net34475), .Y(n4301) );
  NBUFFX2_LVT U6052 ( .A(net34475), .Y(n4302) );
  NBUFFX2_LVT U6053 ( .A(net34475), .Y(n4303) );
  NBUFFX2_LVT U6054 ( .A(net34475), .Y(n4304) );
  NBUFFX2_LVT U6055 ( .A(net34475), .Y(n4305) );
  NBUFFX2_LVT U6056 ( .A(net34475), .Y(n4306) );
  NBUFFX2_LVT U6057 ( .A(net34475), .Y(n4307) );
  NBUFFX2_LVT U6058 ( .A(net34475), .Y(n4308) );
  NBUFFX2_LVT U6059 ( .A(net34475), .Y(n4309) );
  NBUFFX2_LVT U6060 ( .A(net34475), .Y(n4310) );
  AND2X1_LVT U6061 ( .A1(n9529), .A2(n3590), .Y(n4507) );
  INVX1_LVT U6062 ( .A(n9520), .Y(n9437) );
  NAND2X0_LVT U6063 ( .A1(n3593), .A2(io_fpu_inst[4]), .Y(n9111) );
  INVX1_LVT U6064 ( .A(io_fpu_inst[10]), .Y(n9447) );
  AO21X1_LVT U6065 ( .A1(n9446), .A2(n9105), .A3(n9445), .Y(n4505) );
  NAND2X0_LVT U6066 ( .A1(n9529), .A2(n9446), .Y(n5086) );
  AND2X1_LVT U6067 ( .A1(n2137), .A2(n4507), .Y(n4510) );
  NAND2X0_LVT U6068 ( .A1(n9435), .A2(n9524), .Y(n4508) );
  NAND2X0_LVT U6069 ( .A1(n9438), .A2(n5394), .Y(n5149) );
  AND2X1_LVT U6070 ( .A1(wb_ctrl_mem), .A2(wb_reg_valid), .Y(n9249) );
  OR2X1_LVT U6071 ( .A1(io_dmem_s2_xcpt_pf_st), .A2(io_dmem_s2_xcpt_pf_ld), 
        .Y(n9239) );
  OR3X1_LVT U6072 ( .A1(io_dmem_s2_xcpt_ae_ld), .A2(io_dmem_s2_xcpt_ae_st), 
        .A3(n9239), .Y(n4515) );
  OR2X1_LVT U6073 ( .A1(io_dmem_s2_xcpt_ma_st), .A2(io_dmem_s2_xcpt_ma_ld), 
        .Y(n4514) );
  INVX1_LVT U6074 ( .A(mem_br_target[38]), .Y(n4516) );
  INVX1_LVT U6075 ( .A(mem_br_target[26]), .Y(n4517) );
  MUX21X1_LVT U6076 ( .A1(n_T_918[16]), .A2(mem_br_target[16]), .S0(n4591), 
        .Y(n9356) );
  AND3X1_LVT U6077 ( .A1(n4521), .A2(n4520), .A3(n4519), .Y(n4566) );
  INVX1_LVT U6078 ( .A(mem_br_target[36]), .Y(n4522) );
  INVX1_LVT U6079 ( .A(mem_br_target[27]), .Y(n4523) );
  INVX1_LVT U6080 ( .A(mem_br_target[23]), .Y(n4524) );
  INVX1_LVT U6081 ( .A(mem_br_target[18]), .Y(n4525) );
  INVX1_LVT U6082 ( .A(mem_br_target[14]), .Y(n4526) );
  INVX1_LVT U6083 ( .A(mem_br_target[12]), .Y(n4527) );
  INVX1_LVT U6084 ( .A(mem_br_target[8]), .Y(n4528) );
  MUX21X1_LVT U6085 ( .A1(n3222), .A2(n4528), .S0(n3792), .Y(n9511) );
  INVX1_LVT U6086 ( .A(mem_br_target[7]), .Y(n4529) );
  MUX21X1_LVT U6087 ( .A1(n3214), .A2(n4529), .S0(n4591), .Y(n9499) );
  INVX1_LVT U6088 ( .A(mem_br_target[3]), .Y(n4530) );
  MUX21X1_LVT U6089 ( .A1(n3208), .A2(n4530), .S0(n4591), .Y(n9503) );
  INVX1_LVT U6090 ( .A(ibuf_io_pc[0]), .Y(n4531) );
  OA21X1_LVT U6091 ( .A1(io_imem_resp_valid), .A2(ibuf_io_inst_0_valid), .A3(
        n4531), .Y(n4536) );
  MUX21X1_LVT U6092 ( .A1(n_T_918[2]), .A2(mem_br_target[2]), .S0(n3792), .Y(
        n9334) );
  INVX1_LVT U6093 ( .A(mem_br_target[1]), .Y(n4533) );
  AND4X1_LVT U6094 ( .A1(n4537), .A2(n4536), .A3(n4535), .A4(n4534), .Y(n4542)
         );
  INVX1_LVT U6095 ( .A(mem_br_target[5]), .Y(n4538) );
  MUX21X1_LVT U6096 ( .A1(n3109), .A2(n4538), .S0(n4591), .Y(n9484) );
  INVX1_LVT U6097 ( .A(mem_br_target[4]), .Y(n4539) );
  MUX21X1_LVT U6098 ( .A1(n3112), .A2(n4539), .S0(n3792), .Y(n9495) );
  AND4X1_LVT U6099 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .Y(n4548)
         );
  INVX1_LVT U6100 ( .A(mem_br_target[9]), .Y(n4544) );
  MUX21X1_LVT U6101 ( .A1(n3108), .A2(n4544), .S0(n4591), .Y(n9507) );
  INVX1_LVT U6102 ( .A(mem_br_target[6]), .Y(n4545) );
  MUX21X1_LVT U6103 ( .A1(n3217), .A2(n4545), .S0(n3792), .Y(n9485) );
  AND4X1_LVT U6104 ( .A1(n4549), .A2(n4548), .A3(n4547), .A4(n4546), .Y(n4552)
         );
  INVX1_LVT U6105 ( .A(mem_br_target[17]), .Y(n4550) );
  AND2X1_LVT U6106 ( .A1(n4552), .A2(n4551), .Y(n4553) );
  AND4X1_LVT U6107 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .Y(n4559)
         );
  AND4X1_LVT U6108 ( .A1(n4561), .A2(n4560), .A3(n4559), .A4(n4558), .Y(n4564)
         );
  INVX1_LVT U6109 ( .A(mem_br_target[31]), .Y(n4562) );
  AND4X1_LVT U6110 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .Y(n4596)
         );
  INVX1_LVT U6111 ( .A(mem_br_target[37]), .Y(n4567) );
  MUX21X1_LVT U6112 ( .A1(n_T_918[35]), .A2(mem_br_target[35]), .S0(n4591), 
        .Y(n9374) );
  INVX1_LVT U6113 ( .A(mem_br_target[29]), .Y(n4568) );
  INVX1_LVT U6114 ( .A(mem_br_target[10]), .Y(n4569) );
  INVX1_LVT U6115 ( .A(mem_br_target[13]), .Y(n4570) );
  INVX1_LVT U6116 ( .A(mem_br_target[11]), .Y(n4571) );
  INVX1_LVT U6117 ( .A(mem_br_target[19]), .Y(n4572) );
  MUX21X1_LVT U6118 ( .A1(n_T_918[39]), .A2(n3205), .S0(n9470), .Y(n4573) );
  NOR4X1_LVT U6119 ( .A1(n4577), .A2(n4576), .A3(n4575), .A4(n4574), .Y(n4595)
         );
  INVX1_LVT U6120 ( .A(mem_br_target[20]), .Y(n4578) );
  INVX1_LVT U6121 ( .A(mem_br_target[22]), .Y(n4579) );
  INVX1_LVT U6122 ( .A(mem_br_target[33]), .Y(n4580) );
  INVX1_LVT U6123 ( .A(mem_br_target[25]), .Y(n4581) );
  NAND4X0_LVT U6124 ( .A1(n4585), .A2(n4584), .A3(n4583), .A4(n4582), .Y(n4588) );
  INVX1_LVT U6125 ( .A(mem_br_target[30]), .Y(n4586) );
  NOR4X1_LVT U6126 ( .A1(n4590), .A2(n4589), .A3(n4588), .A4(n4587), .Y(n4594)
         );
  INVX1_LVT U6127 ( .A(mem_br_target[32]), .Y(n4592) );
  NAND4X0_LVT U6128 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .Y(n4614) );
  NOR3X0_LVT U6129 ( .A1(n4598), .A2(n4597), .A3(n9482), .Y(n4612) );
  OA21X1_LVT U6130 ( .A1(n_T_698[31]), .A2(n9502), .A3(n4600), .Y(n4601) );
  OA21X1_LVT U6131 ( .A1(n_T_698[32]), .A2(n9505), .A3(n4601), .Y(n4611) );
  OAI22X1_LVT U6132 ( .A1(n_T_698[27]), .A2(n9489), .A3(n_T_698[29]), .A4(
        n9504), .Y(n4608) );
  OA22X1_LVT U6133 ( .A1(n_T_698[19]), .A2(n9510), .A3(n_T_698[25]), .A4(n9497), .Y(n4604) );
  NAND4X0_LVT U6134 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .Y(n4607) );
  NOR4X1_LVT U6135 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .Y(n4610)
         );
  NAND4X0_LVT U6136 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n3204), .Y(n4613) );
  NOR3X0_LVT U6137 ( .A1(ex_reg_valid), .A2(ex_reg_replay), .A3(
        ex_reg_xcpt_interrupt), .Y(n9426) );
  INVX1_LVT U6138 ( .A(n9426), .Y(n5089) );
  MUX21X1_LVT U6139 ( .A1(n4614), .A2(n4613), .S0(n5089), .Y(
        io_imem_bht_update_bits_mispredict) );
  AND2X1_LVT U6140 ( .A1(ibuf_io_inst_0_valid), .A2(n9418), .Y(n9417) );
  NAND3X0_LVT U6141 ( .A1(n4618), .A2(io_fpu_dec_ren1), .A3(n4846), .Y(n4638)
         );
  AND4X1_LVT U6142 ( .A1(n4622), .A2(n4621), .A3(n4620), .A4(n4619), .Y(n4947)
         );
  NAND3X0_LVT U6143 ( .A1(n4947), .A2(io_fpu_dec_wen), .A3(n4946), .Y(n4637)
         );
  NAND4X0_LVT U6144 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(io_fpu_dec_ren3), 
        .Y(n4626) );
  OR3X1_LVT U6145 ( .A1(n4628), .A2(n4627), .A3(n4626), .Y(n4636) );
  NAND4X0_LVT U6146 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .Y(n4858) );
  NAND3X0_LVT U6147 ( .A1(n4634), .A2(io_fpu_dec_ren2), .A3(n4633), .Y(n4635)
         );
  NAND4X0_LVT U6148 ( .A1(n4638), .A2(n4637), .A3(n4636), .A4(n4635), .Y(n4639) );
  AO21X1_LVT U6149 ( .A1(mem_ctrl_wfd), .A2(n4639), .A3(csr_io_singleStep), 
        .Y(n4640) );
  NAND2X0_LVT U6150 ( .A1(n4640), .A2(mem_reg_valid), .Y(n4746) );
  OA22X1_LVT U6151 ( .A1(n3124), .A2(n4708), .A3(n3086), .A4(n4675), .Y(n4645)
         );
  NAND2X0_LVT U6152 ( .A1(n4729), .A2(n_T_1298[2]), .Y(n4644) );
  NAND2X0_LVT U6153 ( .A1(n4731), .A2(n_T_1298[0]), .Y(n4643) );
  NAND3X0_LVT U6154 ( .A1(n4645), .A2(n4644), .A3(n4643), .Y(n4650) );
  OA22X1_LVT U6155 ( .A1(n3125), .A2(n4708), .A3(n3088), .A4(n4675), .Y(n4648)
         );
  NAND2X0_LVT U6156 ( .A1(n4729), .A2(n_T_1298[6]), .Y(n4647) );
  NAND2X0_LVT U6157 ( .A1(n4731), .A2(n_T_1298[4]), .Y(n4646) );
  NAND3X0_LVT U6158 ( .A1(n4648), .A2(n4647), .A3(n4646), .Y(n4649) );
  MUX21X1_LVT U6159 ( .A1(n4650), .A2(n4649), .S0(
        ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4661) );
  NAND2X0_LVT U6160 ( .A1(n4731), .A2(n_T_1298[8]), .Y(n4652) );
  NAND2X0_LVT U6161 ( .A1(n4732), .A2(n_T_1298[9]), .Y(n4651) );
  NAND4X0_LVT U6162 ( .A1(n4652), .A2(n4651), .A3(n4733), .A4(n4719), .Y(n4659) );
  AO22X1_LVT U6163 ( .A1(n_T_1298[11]), .A2(n4730), .A3(n4729), .A4(
        n_T_1298[10]), .Y(n4658) );
  AO22X1_LVT U6164 ( .A1(n_T_1298[15]), .A2(n4730), .A3(n4731), .A4(
        n_T_1298[12]), .Y(n4656) );
  NAND2X0_LVT U6165 ( .A1(n4732), .A2(n_T_1298[13]), .Y(n4654) );
  NAND2X0_LVT U6166 ( .A1(n4729), .A2(n_T_1298[14]), .Y(n4653) );
  NAND3X0_LVT U6167 ( .A1(n4654), .A2(ibuf_io_inst_0_bits_inst_rd[2]), .A3(
        n4653), .Y(n4655) );
  OA21X1_LVT U6168 ( .A1(n4656), .A2(n4655), .A3(
        ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4657) );
  OA22X1_LVT U6169 ( .A1(n4659), .A2(n4658), .A3(
        ibuf_io_inst_0_bits_inst_rd[4]), .A4(n4657), .Y(n4660) );
  AO21X1_LVT U6170 ( .A1(n4662), .A2(n4661), .A3(n4660), .Y(n4683) );
  OA22X1_LVT U6171 ( .A1(n3126), .A2(n4708), .A3(n3087), .A4(n4675), .Y(n4665)
         );
  AND2X1_LVT U6172 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(n4662), .Y(n4666) );
  AND2X1_LVT U6173 ( .A1(n4666), .A2(n4733), .Y(n4717) );
  NAND2X0_LVT U6174 ( .A1(n4731), .A2(n_T_1298[16]), .Y(n4664) );
  NAND2X0_LVT U6175 ( .A1(n4729), .A2(n_T_1298[18]), .Y(n4663) );
  NAND4X0_LVT U6176 ( .A1(n4665), .A2(n4717), .A3(n4664), .A4(n4663), .Y(n4671) );
  OA22X1_LVT U6177 ( .A1(n3239), .A2(n4708), .A3(n3114), .A4(n4675), .Y(n4669)
         );
  AND2X1_LVT U6178 ( .A1(n4666), .A2(ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4698) );
  NAND2X0_LVT U6179 ( .A1(n4731), .A2(n_T_1298[20]), .Y(n4668) );
  NAND2X0_LVT U6180 ( .A1(n4729), .A2(n_T_1298[22]), .Y(n4667) );
  NAND4X0_LVT U6181 ( .A1(n4669), .A2(n4698), .A3(n4668), .A4(n4667), .Y(n4670) );
  NAND2X0_LVT U6182 ( .A1(n1699), .A2(n3039), .Y(n9286) );
  AND4X1_LVT U6183 ( .A1(n4671), .A2(n4670), .A3(io_fpu_dec_wen), .A4(n9286), 
        .Y(n4682) );
  OA22X1_LVT U6184 ( .A1(n3085), .A2(n4708), .A3(n3116), .A4(n4675), .Y(n4674)
         );
  AND2X1_LVT U6185 ( .A1(ibuf_io_inst_0_bits_inst_rd[4]), .A2(
        ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4676) );
  AND2X1_LVT U6186 ( .A1(n4733), .A2(n4676), .Y(n4711) );
  NAND2X0_LVT U6187 ( .A1(n4731), .A2(n_T_1298[24]), .Y(n4673) );
  NAND2X0_LVT U6188 ( .A1(n4729), .A2(n_T_1298[26]), .Y(n4672) );
  NAND4X0_LVT U6189 ( .A1(n4674), .A2(n4711), .A3(n4673), .A4(n4672), .Y(n4681) );
  OA22X1_LVT U6190 ( .A1(n3241), .A2(n4708), .A3(n3084), .A4(n4675), .Y(n4679)
         );
  AND2X1_LVT U6191 ( .A1(n4676), .A2(ibuf_io_inst_0_bits_inst_rd[2]), .Y(n4727) );
  NAND2X0_LVT U6192 ( .A1(n4731), .A2(n_T_1298[28]), .Y(n4678) );
  NAND2X0_LVT U6193 ( .A1(n4729), .A2(n_T_1298[30]), .Y(n4677) );
  NAND4X0_LVT U6194 ( .A1(n4679), .A2(n4727), .A3(n4678), .A4(n4677), .Y(n4680) );
  NAND4X0_LVT U6195 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .Y(n4745) );
  AND2X1_LVT U6196 ( .A1(n4700), .A2(n4733), .Y(n4691) );
  NAND2X0_LVT U6197 ( .A1(n4691), .A2(n4731), .Y(n4684) );
  AND2X1_LVT U6198 ( .A1(id_ctrl_wxd), .A2(n4684), .Y(n5054) );
  NAND2X0_LVT U6199 ( .A1(n4687), .A2(n4686), .Y(n4696) );
  NAND2X0_LVT U6200 ( .A1(wb_ctrl_wxd), .A2(wb_reg_valid), .Y(n5402) );
  NAND2X0_LVT U6201 ( .A1(div_io_resp_valid), .A2(n5402), .Y(n5415) );
  AO21X1_LVT U6202 ( .A1(n_T_1187[3]), .A2(n4730), .A3(n4692), .Y(n4694) );
  AO22X1_LVT U6203 ( .A1(n4729), .A2(n_T_1187[2]), .A3(n_T_1187[1]), .A4(n4732), .Y(n4693) );
  OA22X1_LVT U6204 ( .A1(n4696), .A2(n4695), .A3(n4694), .A4(n4693), .Y(n4715)
         );
  AO22X1_LVT U6205 ( .A1(n_T_1187[23]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[22]), .Y(n4706) );
  NAND2X0_LVT U6206 ( .A1(n4731), .A2(n_T_1187[20]), .Y(n4699) );
  NAND2X0_LVT U6207 ( .A1(n4732), .A2(n_T_1187[21]), .Y(n4697) );
  NAND3X0_LVT U6208 ( .A1(n4699), .A2(n4698), .A3(n4697), .Y(n4705) );
  AO22X1_LVT U6209 ( .A1(n_T_1187[7]), .A2(n4730), .A3(n4729), .A4(n_T_1187[6]), .Y(n4704) );
  NAND2X0_LVT U6210 ( .A1(n4731), .A2(n_T_1187[4]), .Y(n4702) );
  NAND2X0_LVT U6211 ( .A1(n4732), .A2(n_T_1187[5]), .Y(n4701) );
  NAND4X0_LVT U6212 ( .A1(n4702), .A2(n4701), .A3(
        ibuf_io_inst_0_bits_inst_rd[2]), .A4(n4700), .Y(n4703) );
  OA22X1_LVT U6213 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .Y(n4714)
         );
  OA22X1_LVT U6214 ( .A1(n3135), .A2(n4708), .A3(n3265), .A4(n4707), .Y(n4712)
         );
  NAND2X0_LVT U6215 ( .A1(n4732), .A2(n_T_1187[25]), .Y(n4710) );
  NAND2X0_LVT U6216 ( .A1(n4731), .A2(n_T_1187[24]), .Y(n4709) );
  NAND4X0_LVT U6217 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .Y(n4713) );
  AND4X1_LVT U6218 ( .A1(n5054), .A2(n4715), .A3(n4714), .A4(n4713), .Y(n4743)
         );
  AO22X1_LVT U6219 ( .A1(n_T_1187[19]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[18]), .Y(n4725) );
  NAND2X0_LVT U6220 ( .A1(n4731), .A2(n_T_1187[16]), .Y(n4718) );
  NAND2X0_LVT U6221 ( .A1(n4732), .A2(n_T_1187[17]), .Y(n4716) );
  NAND3X0_LVT U6222 ( .A1(n4718), .A2(n4717), .A3(n4716), .Y(n4724) );
  AO22X1_LVT U6223 ( .A1(n_T_1187[15]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[14]), .Y(n4723) );
  NAND2X0_LVT U6224 ( .A1(n4731), .A2(n_T_1187[12]), .Y(n4721) );
  NAND2X0_LVT U6225 ( .A1(n4732), .A2(n_T_1187[13]), .Y(n4720) );
  AND2X1_LVT U6226 ( .A1(n4719), .A2(ibuf_io_inst_0_bits_inst_rd[3]), .Y(n4734) );
  NAND4X0_LVT U6227 ( .A1(n4721), .A2(n4720), .A3(
        ibuf_io_inst_0_bits_inst_rd[2]), .A4(n4734), .Y(n4722) );
  OA22X1_LVT U6228 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .Y(n4742)
         );
  AO22X1_LVT U6229 ( .A1(n_T_1187[31]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[30]), .Y(n4740) );
  NAND2X0_LVT U6230 ( .A1(n4731), .A2(n_T_1187[28]), .Y(n4728) );
  NAND2X0_LVT U6231 ( .A1(n4732), .A2(n_T_1187[29]), .Y(n4726) );
  NAND3X0_LVT U6232 ( .A1(n4728), .A2(n4727), .A3(n4726), .Y(n4739) );
  AO22X1_LVT U6233 ( .A1(n_T_1187[11]), .A2(n4730), .A3(n4729), .A4(
        n_T_1187[10]), .Y(n4738) );
  NAND2X0_LVT U6234 ( .A1(n4731), .A2(n_T_1187[8]), .Y(n4736) );
  NAND2X0_LVT U6235 ( .A1(n4732), .A2(n_T_1187[9]), .Y(n4735) );
  NAND4X0_LVT U6236 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .Y(n4737) );
  OA22X1_LVT U6237 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .Y(n4741)
         );
  NAND3X0_LVT U6238 ( .A1(n4743), .A2(n4742), .A3(n4741), .Y(n4744) );
  NAND3X0_LVT U6239 ( .A1(n4746), .A2(n4745), .A3(n4744), .Y(n9285) );
  AND2X1_LVT U6240 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n2877), .Y(
        n4971) );
  NAND2X0_LVT U6241 ( .A1(ibuf_io_inst_0_bits_inst_rs1[0]), .A2(n2790), .Y(
        n4968) );
  INVX1_LVT U6242 ( .A(n4968), .Y(n4749) );
  AO22X1_LVT U6243 ( .A1(n6972), .A2(n_T_1298[3]), .A3(n6974), .A4(n_T_1298[1]), .Y(n4756) );
  AND2X1_LVT U6244 ( .A1(n4747), .A2(n2876), .Y(n4970) );
  AO22X1_LVT U6245 ( .A1(n6946), .A2(n_T_1298[7]), .A3(n6931), .A4(n_T_1298[6]), .Y(n4755) );
  NAND2X0_LVT U6246 ( .A1(n6957), .A2(n_T_1298[0]), .Y(n4751) );
  NAND2X0_LVT U6247 ( .A1(n6954), .A2(n_T_1298[5]), .Y(n4750) );
  NAND4X0_LVT U6248 ( .A1(n4751), .A2(n6963), .A3(n4750), .A4(n6956), .Y(n4754) );
  AO22X1_LVT U6249 ( .A1(n6926), .A2(n_T_1298[4]), .A3(n6948), .A4(n_T_1298[2]), .Y(n4753) );
  AO22X1_LVT U6250 ( .A1(n6972), .A2(n_T_1298[11]), .A3(n6946), .A4(
        n_T_1298[15]), .Y(n4762) );
  AO22X1_LVT U6251 ( .A1(n6974), .A2(n_T_1298[9]), .A3(n6926), .A4(
        n_T_1298[12]), .Y(n4761) );
  AO22X1_LVT U6252 ( .A1(n6957), .A2(n_T_1298[8]), .A3(n6948), .A4(
        n_T_1298[10]), .Y(n4760) );
  NAND2X0_LVT U6253 ( .A1(n6931), .A2(n_T_1298[14]), .Y(n4758) );
  NAND2X0_LVT U6254 ( .A1(n6954), .A2(n_T_1298[13]), .Y(n4757) );
  AO22X1_LVT U6255 ( .A1(n6946), .A2(n_T_1298[23]), .A3(n6957), .A4(
        n_T_1298[16]), .Y(n4768) );
  AO22X1_LVT U6256 ( .A1(n6974), .A2(n_T_1298[17]), .A3(n6954), .A4(
        n_T_1298[21]), .Y(n4767) );
  OA22X1_LVT U6257 ( .A1(n3238), .A2(n6955), .A3(n3117), .A4(n6947), .Y(n4765)
         );
  AND2X1_LVT U6258 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n6956), .Y(
        n6924) );
  NAND2X0_LVT U6259 ( .A1(n6948), .A2(n_T_1298[18]), .Y(n4764) );
  NAND2X0_LVT U6260 ( .A1(n6972), .A2(n_T_1298[19]), .Y(n4763) );
  OR3X1_LVT U6261 ( .A1(n4766), .A2(n4767), .A3(n4768), .Y(n4780) );
  NAND2X0_LVT U6262 ( .A1(n6974), .A2(n_T_1298[25]), .Y(n4770) );
  AND2X1_LVT U6263 ( .A1(ibuf_io_inst_0_bits_inst_rs1[4]), .A2(n2825), .Y(
        n6917) );
  NAND2X0_LVT U6264 ( .A1(n6946), .A2(n_T_1298[31]), .Y(n4769) );
  AND3X1_LVT U6265 ( .A1(n4770), .A2(n6917), .A3(n4769), .Y(n4778) );
  OA22X1_LVT U6266 ( .A1(n3237), .A2(n4771), .A3(n3123), .A4(n6955), .Y(n4777)
         );
  OA22X1_LVT U6267 ( .A1(n3084), .A2(n4772), .A3(n3118), .A4(n6947), .Y(n4776)
         );
  OA22X1_LVT U6268 ( .A1(n4774), .A2(n3085), .A3(n3232), .A4(n4773), .Y(n4775)
         );
  NAND4X0_LVT U6269 ( .A1(n4778), .A2(n4777), .A3(n4776), .A4(n4775), .Y(n4779) );
  NAND2X0_LVT U6270 ( .A1(ibuf_io_inst_0_bits_raw[28]), .A2(
        ibuf_io_inst_0_bits_raw[27]), .Y(n4802) );
  OA22X1_LVT U6271 ( .A1(n3124), .A2(n4802), .A3(n3247), .A4(n4801), .Y(n4784)
         );
  OA22X1_LVT U6272 ( .A1(n3254), .A2(n4804), .A3(n3086), .A4(n4803), .Y(n4783)
         );
  AND2X1_LVT U6273 ( .A1(n4784), .A2(n4783), .Y(n4794) );
  OA22X1_LVT U6274 ( .A1(n3240), .A2(n4802), .A3(n3115), .A4(n4801), .Y(n4786)
         );
  OA22X1_LVT U6275 ( .A1(n3242), .A2(n4804), .A3(n3119), .A4(n4803), .Y(n4785)
         );
  AND2X1_LVT U6276 ( .A1(n4786), .A2(n4785), .Y(n4793) );
  OA22X1_LVT U6277 ( .A1(n3125), .A2(n4802), .A3(n3248), .A4(n4801), .Y(n4788)
         );
  OA22X1_LVT U6278 ( .A1(n3253), .A2(n4804), .A3(n3088), .A4(n4803), .Y(n4787)
         );
  AND2X1_LVT U6279 ( .A1(n4788), .A2(n4787), .Y(n4792) );
  OA22X1_LVT U6280 ( .A1(n3236), .A2(n4802), .A3(n3121), .A4(n4801), .Y(n4790)
         );
  OA22X1_LVT U6281 ( .A1(n3235), .A2(n4804), .A3(n3120), .A4(n4803), .Y(n4789)
         );
  AND2X1_LVT U6282 ( .A1(n4790), .A2(n4789), .Y(n4791) );
  MUX41X1_LVT U6283 ( .A1(n4794), .A3(n4793), .A2(n4792), .A4(n4791), .S0(
        n1859), .S1(n2674), .Y(n4812) );
  OA22X1_LVT U6284 ( .A1(n3126), .A2(n4802), .A3(n3250), .A4(n4801), .Y(n4796)
         );
  OA22X1_LVT U6285 ( .A1(n3252), .A2(n4804), .A3(n3087), .A4(n4803), .Y(n4795)
         );
  AND2X1_LVT U6286 ( .A1(n4796), .A2(n4795), .Y(n4810) );
  OA22X1_LVT U6287 ( .A1(n3085), .A2(n4802), .A3(n3232), .A4(n4801), .Y(n4798)
         );
  OA22X1_LVT U6288 ( .A1(n3237), .A2(n4804), .A3(n3116), .A4(n4803), .Y(n4797)
         );
  AND2X1_LVT U6289 ( .A1(n4798), .A2(n4797), .Y(n4809) );
  OA22X1_LVT U6290 ( .A1(n3239), .A2(n4802), .A3(n3117), .A4(n4801), .Y(n4800)
         );
  OA22X1_LVT U6291 ( .A1(n3238), .A2(n4804), .A3(n3114), .A4(n4803), .Y(n4799)
         );
  AND2X1_LVT U6292 ( .A1(n4800), .A2(n4799), .Y(n4808) );
  OA22X1_LVT U6293 ( .A1(n3241), .A2(n4802), .A3(n3118), .A4(n4801), .Y(n4806)
         );
  OA22X1_LVT U6294 ( .A1(n3123), .A2(n4804), .A3(n3084), .A4(n4803), .Y(n4805)
         );
  AND2X1_LVT U6295 ( .A1(n4806), .A2(n4805), .Y(n4807) );
  MUX41X1_LVT U6296 ( .A1(n4810), .A3(n4809), .A2(n4808), .A4(n4807), .S0(
        n1859), .S1(ibuf_io_inst_0_bits_raw[29]), .Y(n4811) );
  AND2X1_LVT U6297 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(
        ibuf_io_inst_0_bits_inst_rs2[0]), .Y(n4889) );
  AO22X1_LVT U6298 ( .A1(n_T_1298[3]), .A2(n5452), .A3(n5455), .A4(n_T_1298[0]), .Y(n4820) );
  AND2X1_LVT U6299 ( .A1(ibuf_io_inst_0_bits_inst_rs2[0]), .A2(n4813), .Y(
        n4890) );
  AO22X1_LVT U6300 ( .A1(n_T_1298[7]), .A2(n5450), .A3(n5456), .A4(n_T_1298[1]), .Y(n4819) );
  AND2X1_LVT U6301 ( .A1(ibuf_io_inst_0_bits_inst_rs2[1]), .A2(n4815), .Y(
        n4900) );
  AO22X1_LVT U6302 ( .A1(n2034), .A2(n_T_1298[4]), .A3(n_T_1298[6]), .A4(n5449), .Y(n4818) );
  AO22X1_LVT U6303 ( .A1(n5451), .A2(n_T_1298[5]), .A3(n_T_1298[2]), .A4(n5454), .Y(n4817) );
  NOR4X1_LVT U6304 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .Y(n4835)
         );
  OA22X1_LVT U6305 ( .A1(n3236), .A2(n5438), .A3(n3119), .A4(n4905), .Y(n4824)
         );
  INVX1_LVT U6306 ( .A(n5453), .Y(n4880) );
  OA22X1_LVT U6307 ( .A1(n3235), .A2(n4880), .A3(n3115), .A4(n4873), .Y(n4823)
         );
  OA22X1_LVT U6308 ( .A1(n3240), .A2(n4906), .A3(n3120), .A4(n4894), .Y(n4822)
         );
  OA22X1_LVT U6309 ( .A1(n3242), .A2(n5435), .A3(n3121), .A4(n4874), .Y(n4821)
         );
  AO22X1_LVT U6310 ( .A1(n_T_1298[19]), .A2(n5452), .A3(n5454), .A4(
        n_T_1298[18]), .Y(n4828) );
  AO22X1_LVT U6311 ( .A1(n_T_1298[23]), .A2(n5450), .A3(n2034), .A4(
        n_T_1298[20]), .Y(n4827) );
  AO22X1_LVT U6312 ( .A1(n5455), .A2(n_T_1298[16]), .A3(n_T_1298[22]), .A4(
        n5449), .Y(n4826) );
  AO22X1_LVT U6313 ( .A1(n5451), .A2(n_T_1298[21]), .A3(n_T_1298[17]), .A4(
        n5456), .Y(n4825) );
  NOR4X1_LVT U6314 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), .Y(n4834)
         );
  AO22X1_LVT U6315 ( .A1(n_T_1298[27]), .A2(n5452), .A3(n5456), .A4(
        n_T_1298[25]), .Y(n4832) );
  AO22X1_LVT U6316 ( .A1(n_T_1298[31]), .A2(n5450), .A3(n5455), .A4(
        n_T_1298[24]), .Y(n4831) );
  AO22X1_LVT U6317 ( .A1(n2034), .A2(n_T_1298[28]), .A3(n_T_1298[30]), .A4(
        n5449), .Y(n4830) );
  AO22X1_LVT U6318 ( .A1(n5451), .A2(n_T_1298[29]), .A3(n_T_1298[26]), .A4(
        n5454), .Y(n4829) );
  NOR4X1_LVT U6319 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), .Y(n4833)
         );
  MUX41X1_LVT U6320 ( .A1(n4835), .A3(n3181), .A2(n4834), .A4(n4833), .S0(
        n3781), .S1(ibuf_io_inst_0_bits_inst_rs2[4]), .Y(n4836) );
  OA22X1_LVT U6321 ( .A1(n4839), .A2(n4838), .A3(n4837), .A4(n4836), .Y(n4849)
         );
  NAND2X0_LVT U6322 ( .A1(mem_ctrl_mem), .A2(mem_reg_slow_bypass), .Y(n4840)
         );
  NAND3X0_LVT U6323 ( .A1(n4840), .A2(n370), .A3(n3246), .Y(n4841) );
  NOR4X1_LVT U6324 ( .A1(mem_ctrl_csr[0]), .A2(mem_ctrl_csr[2]), .A3(n3279), 
        .A4(n4841), .Y(n4949) );
  NAND2X0_LVT U6325 ( .A1(n5163), .A2(io_fpu_inst[14]), .Y(n4842) );
  NAND2X0_LVT U6326 ( .A1(n2538), .A2(n9288), .Y(n9280) );
  AND2X1_LVT U6327 ( .A1(mem_ctrl_wxd), .A2(mem_reg_valid), .Y(n4948) );
  NAND2X0_LVT U6328 ( .A1(n4846), .A2(n4948), .Y(n4848) );
  OA22X1_LVT U6329 ( .A1(n2512), .A2(n4849), .A3(n4949), .A4(n5094), .Y(n4851)
         );
  NAND2X0_LVT U6330 ( .A1(n1612), .A2(n9432), .Y(n5087) );
  NAND3X0_LVT U6331 ( .A1(n5087), .A2(blocked), .A3(n5065), .Y(n4850) );
  AND3X1_LVT U6332 ( .A1(n4850), .A2(n4851), .A3(n4852), .Y(n4955) );
  AND2X1_LVT U6333 ( .A1(n5396), .A2(n2618), .Y(n1828) );
  NAND2X0_LVT U6334 ( .A1(n5087), .A2(id_reg_fence), .Y(n4854) );
  AND2X1_LVT U6335 ( .A1(ex_ctrl_mem), .A2(ex_reg_valid), .Y(io_dmem_req_valid) );
  INVX1_LVT U6336 ( .A(io_dmem_req_valid), .Y(n4853) );
  AND2X1_LVT U6337 ( .A1(n4853), .A2(io_dmem_ordered), .Y(n5063) );
  AO21X1_LVT U6338 ( .A1(n4855), .A2(n4854), .A3(n5063), .Y(n4954) );
  NAND2X0_LVT U6339 ( .A1(n4856), .A2(n3597), .Y(n4857) );
  NAND2X0_LVT U6340 ( .A1(n1531), .A2(n1532), .Y(n5466) );
  AND2X1_LVT U6341 ( .A1(n5466), .A2(n5421), .Y(n5021) );
  NOR3X0_LVT U6342 ( .A1(n4860), .A2(n4859), .A3(n4858), .Y(n5420) );
  NAND2X0_LVT U6343 ( .A1(n5021), .A2(n5420), .Y(n5093) );
  INVX1_LVT U6344 ( .A(n5044), .Y(n4867) );
  AND2X1_LVT U6345 ( .A1(ex_reg_valid), .A2(ex_ctrl_wxd), .Y(n5009) );
  AND4X1_LVT U6346 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .Y(n5045)
         );
  INVX1_LVT U6347 ( .A(n5045), .Y(n4865) );
  OR3X1_LVT U6348 ( .A1(n4867), .A2(n4866), .A3(n4865), .Y(n5419) );
  NAND2X0_LVT U6349 ( .A1(n4872), .A2(n4871), .Y(n4887) );
  OA22X1_LVT U6350 ( .A1(n3272), .A2(n4894), .A3(n3129), .A4(n4873), .Y(n4878)
         );
  OA22X1_LVT U6351 ( .A1(n3260), .A2(n4880), .A3(n3127), .A4(n4874), .Y(n4877)
         );
  OA22X1_LVT U6352 ( .A1(n4906), .A2(n3259), .A3(n3133), .A4(n4905), .Y(n4876)
         );
  OA22X1_LVT U6353 ( .A1(n5438), .A2(n3266), .A3(n3134), .A4(n5435), .Y(n4875)
         );
  NAND4X0_LVT U6354 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .Y(n4879) );
  AND2X1_LVT U6355 ( .A1(n4879), .A2(n2878), .Y(n4886) );
  NAND2X0_LVT U6356 ( .A1(n5451), .A2(n5436), .Y(n5546) );
  OA22X1_LVT U6357 ( .A1(n3271), .A2(n5546), .A3(n3136), .A4(n6766), .Y(n4884)
         );
  NAND2X0_LVT U6358 ( .A1(n5454), .A2(n5436), .Y(n6422) );
  NAND2X0_LVT U6359 ( .A1(n5452), .A2(n5436), .Y(n5906) );
  NAND2X0_LVT U6360 ( .A1(n5456), .A2(n5436), .Y(n5905) );
  NAND2X0_LVT U6361 ( .A1(n5450), .A2(n5436), .Y(n6767) );
  OA22X1_LVT U6362 ( .A1(n3270), .A2(n6767), .A3(n3132), .A4(n6423), .Y(n4881)
         );
  NAND4X0_LVT U6363 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n4881), .Y(n4885) );
  OAI22X1_LVT U6364 ( .A1(n4888), .A2(n4887), .A3(n4886), .A4(n4885), .Y(n4916) );
  OA22X1_LVT U6365 ( .A1(n4899), .A2(n3267), .A3(n3131), .A4(n4898), .Y(n4893)
         );
  NAND2X0_LVT U6366 ( .A1(n4901), .A2(n_T_1187[28]), .Y(n4892) );
  NAND2X0_LVT U6367 ( .A1(n4900), .A2(n_T_1187[30]), .Y(n4891) );
  OA22X1_LVT U6368 ( .A1(n5438), .A2(n3268), .A3(n3130), .A4(n4894), .Y(n4897)
         );
  NAND2X0_LVT U6369 ( .A1(n2034), .A2(n_T_1187[20]), .Y(n4896) );
  NAND2X0_LVT U6370 ( .A1(n5449), .A2(n_T_1187[22]), .Y(n4895) );
  NAND3X0_LVT U6371 ( .A1(n4897), .A2(n4896), .A3(n4895), .Y(n4913) );
  OA22X1_LVT U6372 ( .A1(n4899), .A2(n3135), .A3(n3089), .A4(n4898), .Y(n4904)
         );
  NAND2X0_LVT U6373 ( .A1(n4900), .A2(n_T_1187[26]), .Y(n4903) );
  NAND2X0_LVT U6374 ( .A1(n4901), .A2(n_T_1187[24]), .Y(n4902) );
  MUX21X1_LVT U6375 ( .A1(n4910), .A2(n4914), .S0(
        ibuf_io_inst_0_bits_inst_rs2[2]), .Y(n4912) );
  OA22X1_LVT U6376 ( .A1(n4906), .A2(n3258), .A3(n3113), .A4(n4905), .Y(n4909)
         );
  NAND2X0_LVT U6377 ( .A1(n5455), .A2(n_T_1187[16]), .Y(n4908) );
  NAND2X0_LVT U6378 ( .A1(n5454), .A2(n_T_1187[18]), .Y(n4907) );
  NAND3X0_LVT U6379 ( .A1(n4909), .A2(n4908), .A3(n4907), .Y(n4911) );
  AOI222X1_LVT U6380 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n5447), .A5(
        n4911), .A6(n4910), .Y(n4915) );
  OA22X1_LVT U6381 ( .A1(n5051), .A2(n5419), .A3(n4916), .A4(n4915), .Y(n4935)
         );
  AND2X1_LVT U6382 ( .A1(ex_reg_valid), .A2(ex_ctrl_div), .Y(n9422) );
  AO21X1_LVT U6383 ( .A1(n5415), .A2(n4917), .A3(n9422), .Y(n4932) );
  NOR2X0_LVT U6384 ( .A1(id_reg_pause), .A2(csr_io_csr_stall), .Y(n4928) );
  AND3X1_LVT U6385 ( .A1(wb_ctrl_wfd), .A2(wb_reg_valid), .A3(io_fpu_dec_ren3), 
        .Y(n4919) );
  NAND4X0_LVT U6386 ( .A1(n4922), .A2(n4921), .A3(n4920), .A4(n4919), .Y(n4923) );
  OR3X1_LVT U6387 ( .A1(n4925), .A2(n4924), .A3(n4923), .Y(n4927) );
  NAND2X0_LVT U6388 ( .A1(csr_io_singleStep), .A2(wb_reg_valid), .Y(n4926) );
  NAND4X0_LVT U6389 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .Y(n4930) );
  AOI21X1_LVT U6390 ( .A1(n4932), .A2(n4931), .A3(n4930), .Y(n4933) );
  OA21X1_LVT U6391 ( .A1(n4935), .A2(n4934), .A3(n4933), .Y(n4936) );
  OA21X1_LVT U6392 ( .A1(n4949), .A2(n5093), .A3(n4936), .Y(n4953) );
  NAND4X0_LVT U6393 ( .A1(n4939), .A2(n4938), .A3(n4937), .A4(wb_reg_valid), 
        .Y(n4940) );
  OR3X1_LVT U6394 ( .A1(n4942), .A2(n4941), .A3(n4940), .Y(n4951) );
  AND2X1_LVT U6395 ( .A1(n4943), .A2(wb_ctrl_mem), .Y(n5175) );
  OA21X1_LVT U6396 ( .A1(wb_ctrl_div), .A2(n5175), .A3(wb_ctrl_wxd), .Y(n5301)
         );
  OA22X1_LVT U6397 ( .A1(n4945), .A2(n3229), .A3(n4944), .A4(n9280), .Y(n4950)
         );
  NAND4X0_LVT U6398 ( .A1(n5054), .A2(n4948), .A3(n4947), .A4(n4946), .Y(n5092) );
  OA22X1_LVT U6399 ( .A1(n4951), .A2(n4950), .A3(n4949), .A4(n5092), .Y(n4952)
         );
  OA22X1_LVT U6400 ( .A1(n3261), .A2(n4969), .A3(n3113), .A4(n4968), .Y(n4958)
         );
  NAND2X0_LVT U6401 ( .A1(n4970), .A2(n_T_1187[18]), .Y(n4957) );
  NAND2X0_LVT U6402 ( .A1(n4971), .A2(n_T_1187[19]), .Y(n4956) );
  NAND3X0_LVT U6403 ( .A1(n4958), .A2(n4957), .A3(n4956), .Y(n4963) );
  OA22X1_LVT U6404 ( .A1(n3275), .A2(n4969), .A3(n3089), .A4(n4968), .Y(n4961)
         );
  NAND2X0_LVT U6405 ( .A1(n4970), .A2(n_T_1187[26]), .Y(n4960) );
  NAND2X0_LVT U6406 ( .A1(n4971), .A2(n_T_1187[27]), .Y(n4959) );
  NAND3X0_LVT U6407 ( .A1(n4961), .A2(n4960), .A3(n4959), .Y(n4962) );
  MUX21X1_LVT U6408 ( .A1(n4963), .A2(n4962), .S0(n2825), .Y(n4964) );
  OR2X1_LVT U6409 ( .A1(n6963), .A2(n4964), .Y(n4979) );
  OA22X1_LVT U6410 ( .A1(n3273), .A2(n4969), .A3(n3130), .A4(n4968), .Y(n4967)
         );
  NAND2X0_LVT U6411 ( .A1(n4970), .A2(n_T_1187[22]), .Y(n4966) );
  NAND2X0_LVT U6412 ( .A1(n4971), .A2(n_T_1187[23]), .Y(n4965) );
  NAND3X0_LVT U6413 ( .A1(n4967), .A2(n4966), .A3(n4965), .Y(n4976) );
  OA22X1_LVT U6414 ( .A1(n3274), .A2(n4969), .A3(n3131), .A4(n4968), .Y(n4974)
         );
  NAND2X0_LVT U6415 ( .A1(n4970), .A2(n_T_1187[30]), .Y(n4973) );
  NAND2X0_LVT U6416 ( .A1(n4971), .A2(n_T_1187[31]), .Y(n4972) );
  NAND3X0_LVT U6417 ( .A1(n4974), .A2(n4973), .A3(n4972), .Y(n4975) );
  MUX21X1_LVT U6418 ( .A1(n4976), .A2(n4975), .S0(n2825), .Y(n4977) );
  OR2X1_LVT U6419 ( .A1(n6963), .A2(n4977), .Y(n4978) );
  MUX21X1_LVT U6420 ( .A1(n4979), .A2(n4978), .S0(n2038), .Y(n5008) );
  OA21X1_LVT U6421 ( .A1(n3132), .A2(n6949), .A3(n6963), .Y(n4982) );
  NAND2X0_LVT U6422 ( .A1(n4044), .A2(n_T_1187[2]), .Y(n4981) );
  AND2X1_LVT U6423 ( .A1(n6946), .A2(n6956), .Y(n8931) );
  NAND2X0_LVT U6424 ( .A1(n3968), .A2(n_T_1187[7]), .Y(n4980) );
  NAND3X0_LVT U6425 ( .A1(n4982), .A2(n4980), .A3(n4981), .Y(n4999) );
  NAND2X0_LVT U6426 ( .A1(n6974), .A2(n6956), .Y(n6945) );
  NAND2X0_LVT U6427 ( .A1(n3972), .A2(n_T_1187[3]), .Y(n4983) );
  OA21X1_LVT U6428 ( .A1(n3128), .A2(n6945), .A3(n4983), .Y(n4986) );
  AND2X1_LVT U6429 ( .A1(n6954), .A2(n6956), .Y(n8901) );
  NAND2X0_LVT U6430 ( .A1(n3967), .A2(n_T_1187[5]), .Y(n4985) );
  NAND2X0_LVT U6431 ( .A1(n9040), .A2(n_T_1187[6]), .Y(n4984) );
  NAND3X0_LVT U6432 ( .A1(n4986), .A2(n4984), .A3(n4985), .Y(n4998) );
  NAND2X0_LVT U6433 ( .A1(n6972), .A2(n_T_1187[11]), .Y(n4987) );
  OA21X1_LVT U6434 ( .A1(n3127), .A2(n6947), .A3(n4987), .Y(n4990) );
  NAND2X0_LVT U6435 ( .A1(n6948), .A2(n_T_1187[10]), .Y(n4989) );
  NAND2X0_LVT U6436 ( .A1(n6974), .A2(n_T_1187[9]), .Y(n4988) );
  NAND3X0_LVT U6437 ( .A1(n4990), .A2(n4989), .A3(n4988), .Y(n4996) );
  NAND2X0_LVT U6438 ( .A1(n6946), .A2(n_T_1187[15]), .Y(n4991) );
  OA21X1_LVT U6439 ( .A1(n3260), .A2(n6955), .A3(n4991), .Y(n4994) );
  NAND2X0_LVT U6440 ( .A1(n6954), .A2(n_T_1187[13]), .Y(n4993) );
  NAND2X0_LVT U6441 ( .A1(n6957), .A2(n_T_1187[8]), .Y(n4992) );
  NAND3X0_LVT U6442 ( .A1(n4994), .A2(n4993), .A3(n4992), .Y(n4995) );
  OR3X1_LVT U6443 ( .A1(n4999), .A2(n4998), .A3(n4997), .Y(n5007) );
  OR3X1_LVT U6444 ( .A1(n5005), .A2(n5004), .A3(n5003), .Y(n5006) );
  NAND2X0_LVT U6445 ( .A1(n5037), .A2(n5009), .Y(n5013) );
  OA21X1_LVT U6446 ( .A1(n9280), .A2(n9281), .A3(n9385), .Y(n5029) );
  AO22X1_LVT U6447 ( .A1(wb_ctrl_wfd), .A2(io_fpu_dec_wen), .A3(n5054), .A4(
        n5301), .Y(n5020) );
  AND4X1_LVT U6448 ( .A1(n5016), .A2(wb_reg_valid), .A3(n5015), .A4(n5014), 
        .Y(n5019) );
  NAND4X0_LVT U6449 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .Y(n9278) );
  AO22X1_LVT U6450 ( .A1(io_fpu_dec_ren2), .A2(wb_ctrl_wfd), .A3(n5021), .A4(
        n5301), .Y(n5028) );
  AND4X1_LVT U6451 ( .A1(n5024), .A2(n5023), .A3(wb_reg_valid), .A4(n5022), 
        .Y(n5027) );
  NAND4X0_LVT U6452 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .Y(n9277) );
  AND3X1_LVT U6453 ( .A1(n5029), .A2(n9278), .A3(n9277), .Y(n5059) );
  AND2X1_LVT U6454 ( .A1(n5031), .A2(n5030), .Y(n5034) );
  AND4X1_LVT U6455 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5032), .Y(n5053)
         );
  NAND2X0_LVT U6456 ( .A1(n5053), .A2(io_fpu_dec_wen), .Y(n5049) );
  NAND3X0_LVT U6457 ( .A1(n2567), .A2(io_fpu_dec_ren1), .A3(n5037), .Y(n5048)
         );
  NAND4X0_LVT U6458 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(io_fpu_dec_ren3), 
        .Y(n5041) );
  OR3X1_LVT U6459 ( .A1(n5043), .A2(n5042), .A3(n5041), .Y(n5047) );
  NAND3X0_LVT U6460 ( .A1(n5045), .A2(io_fpu_dec_ren2), .A3(n5044), .Y(n5046)
         );
  NAND4X0_LVT U6461 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .Y(n5050) );
  NAND2X0_LVT U6462 ( .A1(n5050), .A2(ex_ctrl_wfd), .Y(n5057) );
  INVX1_LVT U6463 ( .A(csr_io_singleStep), .Y(n5056) );
  NAND4X0_LVT U6464 ( .A1(n5054), .A2(ex_ctrl_wxd), .A3(n5053), .A4(n5052), 
        .Y(n5055) );
  NAND3X0_LVT U6465 ( .A1(n5057), .A2(n5056), .A3(n5055), .Y(n5058) );
  NAND2X0_LVT U6466 ( .A1(n5058), .A2(ex_reg_valid), .Y(n9279) );
  NAND3X0_LVT U6467 ( .A1(n9279), .A2(n5059), .A3(n5060), .Y(n5061) );
  NOR3X0_LVT U6468 ( .A1(n5061), .A2(n9282), .A3(n9285), .Y(n5062) );
  NAND2X0_LVT U6469 ( .A1(io_dmem_req_valid), .A2(n5064), .Y(n5095) );
  NAND2X0_LVT U6470 ( .A1(n9521), .A2(io_fpu_inst[28]), .Y(n5154) );
  AND2X1_LVT U6471 ( .A1(n5066), .A2(io_fpu_inst[5]), .Y(n9431) );
  NAND2X0_LVT U6472 ( .A1(io_fpu_inst[3]), .A2(n5067), .Y(n9110) );
  AO21X1_LVT U6473 ( .A1(n9431), .A2(n5070), .A3(n5123), .Y(n9287) );
  NAND2X0_LVT U6474 ( .A1(n5071), .A2(n3597), .Y(n1628) );
  NAND2X0_LVT U6475 ( .A1(io_fpu_inst[13]), .A2(io_fpu_inst[4]), .Y(n9089) );
  AND2X1_LVT U6476 ( .A1(n2618), .A2(n5088), .Y(N286) );
  OA21X1_LVT U6477 ( .A1(n9105), .A2(n9520), .A3(n5072), .Y(n5073) );
  AND2X1_LVT U6478 ( .A1(n559), .A2(io_dmem_req_bits_cmd[0]), .Y(n5078) );
  NAND4X0_LVT U6479 ( .A1(ex_ctrl_mem), .A2(n5078), .A3(n3122), .A4(n3244), 
        .Y(n996) );
  AND3X1_LVT U6480 ( .A1(ex_ctrl_mem), .A2(n560), .A3(n3122), .Y(n5090) );
  OR2X1_LVT U6481 ( .A1(n559), .A2(io_dmem_req_bits_cmd[2]), .Y(n5079) );
  NAND3X0_LVT U6482 ( .A1(n5090), .A2(n3245), .A3(n5079), .Y(n882) );
  NAND2X0_LVT U6483 ( .A1(io_imem_bht_update_bits_branch), .A2(
        io_imem_bht_update_bits_taken), .Y(n5080) );
  AND2X1_LVT U6484 ( .A1(n555), .A2(n5080), .Y(n5084) );
  INVX1_LVT U6485 ( .A(n5080), .Y(n5085) );
  AND2X1_LVT U6486 ( .A1(n5085), .A2(n_T_844_10_), .Y(n5081) );
  AO21X1_LVT U6487 ( .A1(n5083), .A2(n_T_904[7]), .A3(n5081), .Y(n_T_914[19])
         );
  AO21X1_LVT U6488 ( .A1(n5083), .A2(n_T_904[6]), .A3(n5081), .Y(n_T_914[18])
         );
  AO21X1_LVT U6489 ( .A1(n5083), .A2(n_T_904[5]), .A3(n5081), .Y(n_T_914[17])
         );
  AO21X1_LVT U6490 ( .A1(n5083), .A2(n_T_904[4]), .A3(n5081), .Y(n_T_914[16])
         );
  AO21X1_LVT U6491 ( .A1(n5083), .A2(n_T_904[3]), .A3(n5081), .Y(n_T_914[15])
         );
  AO21X1_LVT U6492 ( .A1(n5083), .A2(n_T_904[2]), .A3(n5081), .Y(n_T_914[14])
         );
  AO21X1_LVT U6493 ( .A1(n5083), .A2(n_T_904[1]), .A3(n5081), .Y(n_T_914[13])
         );
  AO21X1_LVT U6494 ( .A1(n5083), .A2(n_T_904[0]), .A3(n5081), .Y(n_T_914[12])
         );
  AO22X1_LVT U6495 ( .A1(n5085), .A2(n_T_849[11]), .A3(n5083), .A4(n_T_911_11), 
        .Y(n_T_914[11]) );
  AND2X1_LVT U6496 ( .A1(n_T_849[10]), .A2(n5082), .Y(n_T_914[10]) );
  AND2X1_LVT U6497 ( .A1(n_T_849[9]), .A2(n5082), .Y(n_T_914[9]) );
  AND2X1_LVT U6498 ( .A1(n_T_849[8]), .A2(n5082), .Y(n_T_914[8]) );
  AND2X1_LVT U6499 ( .A1(n_T_849[7]), .A2(n5082), .Y(n_T_914[7]) );
  AND2X1_LVT U6500 ( .A1(n_T_849[6]), .A2(n5082), .Y(n_T_914[6]) );
  AND2X1_LVT U6501 ( .A1(n_T_849[5]), .A2(n5082), .Y(n_T_914[5]) );
  AO22X1_LVT U6502 ( .A1(n_T_911[4]), .A2(n5083), .A3(n5085), .A4(n_T_849[4]), 
        .Y(n_T_914[4]) );
  INVX1_LVT U6503 ( .A(io_fpu_inst[23]), .Y(n9441) );
  AO22X1_LVT U6504 ( .A1(n_T_911[3]), .A2(n5083), .A3(n5085), .A4(n2566), .Y(
        n_T_914[3]) );
  INVX1_LVT U6505 ( .A(io_fpu_inst[22]), .Y(n9442) );
  AO222X1_LVT U6506 ( .A1(n570), .A2(n5084), .A3(n_T_911[2]), .A4(n5083), .A5(
        n_T_849[2]), .A6(n5085), .Y(n_T_914[2]) );
  INVX1_LVT U6507 ( .A(io_fpu_inst[21]), .Y(n9443) );
  AO222X1_LVT U6508 ( .A1(n_T_849[1]), .A2(n5085), .A3(n5084), .A4(mem_reg_rvc), .A5(n5083), .A6(n_T_911[1]), .Y(n_T_914[1]) );
  NAND2X0_LVT U6509 ( .A1(mem_reg_valid), .A2(mem_reg_flush_pipe), .Y(n5091)
         );
  AND2X1_LVT U6510 ( .A1(n5089), .A2(n5091), .Y(N290) );
  AND2X1_LVT U6511 ( .A1(io_imem_req_bits_speculative), .A2(mem_reg_valid), 
        .Y(io_imem_bht_update_valid) );
  NAND2X0_LVT U6512 ( .A1(mem_ctrl_wxd), .A2(io_dmem_replay_next), .Y(n5404)
         );
  NAND2X0_LVT U6513 ( .A1(n2498), .A2(io_fpu_nack_mem), .Y(n5096) );
  AND2X1_LVT U6514 ( .A1(n5404), .A2(n5096), .Y(n5169) );
  NAND3X0_LVT U6515 ( .A1(n5102), .A2(n9075), .A3(n3578), .Y(n5103) );
  NAND2X0_LVT U6516 ( .A1(csr_io_decode_0_read_illegal), .A2(n5119), .Y(n5113)
         );
  NOR2X0_LVT U6517 ( .A1(io_fpu_illegal_rm), .A2(csr_io_decode_0_fp_illegal), 
        .Y(n5118) );
  OA21X1_LVT U6518 ( .A1(io_fpu_inst[28]), .A2(n5114), .A3(n9440), .Y(n5115)
         );
  NAND2X0_LVT U6519 ( .A1(csr_io_status_isa[0]), .A2(n5116), .Y(n5117) );
  OA21X1_LVT U6520 ( .A1(n5118), .A2(n1699), .A3(n5117), .Y(n5121) );
  OR2X1_LVT U6521 ( .A1(io_fpu_inst[18]), .A2(io_fpu_inst[17]), .Y(n5128) );
  OR2X1_LVT U6522 ( .A1(io_fpu_inst[15]), .A2(io_fpu_inst[16]), .Y(n5127) );
  OR3X1_LVT U6523 ( .A1(io_fpu_inst[10]), .A2(io_fpu_inst[19]), .A3(
        io_fpu_inst[11]), .Y(n5125) );
  OR3X1_LVT U6524 ( .A1(io_fpu_inst[8]), .A2(io_fpu_inst[9]), .A3(n5125), .Y(
        n5126) );
  OR3X1_LVT U6525 ( .A1(n5128), .A2(n5127), .A3(n5126), .Y(n5158) );
  INVX1_LVT U6526 ( .A(io_fpu_inst[24]), .Y(n5148) );
  NAND3X0_LVT U6527 ( .A1(n5132), .A2(n2565), .A3(n5131), .Y(n5141) );
  AND2X1_LVT U6528 ( .A1(io_fpu_inst[31]), .A2(n9445), .Y(n5136) );
  NAND4X0_LVT U6529 ( .A1(n5139), .A2(n3567), .A3(n5138), .A4(n5137), .Y(n5140) );
  OR3X1_LVT U6530 ( .A1(n5394), .A2(n5154), .A3(n5144), .Y(n5145) );
  NAND2X0_LVT U6531 ( .A1(n2537), .A2(n5146), .Y(n5147) );
  NAND2X0_LVT U6532 ( .A1(io_fpu_inst[22]), .A2(io_fpu_inst[21]), .Y(n5153) );
  OA21X1_LVT U6533 ( .A1(io_fpu_inst[22]), .A2(n9444), .A3(n5153), .Y(n5157)
         );
  NAND2X0_LVT U6534 ( .A1(n5154), .A2(n3079), .Y(n5155) );
  NAND3X0_LVT U6535 ( .A1(n5157), .A2(n5156), .A3(n5155), .Y(n5159) );
  OR3X1_LVT U6536 ( .A1(n5160), .A2(n5159), .A3(n5158), .Y(n5161) );
  NAND2X0_LVT U6537 ( .A1(n9430), .A2(n9118), .Y(n9243) );
  AND3X1_LVT U6538 ( .A1(n9418), .A2(ex_reg_valid), .A3(n9421), .Y(n407) );
  INVX1_LVT U6539 ( .A(n407), .Y(io_fpu_killx) );
  OR3X1_LVT U6540 ( .A1(mem_reg_sfence), .A2(csr_io_status_isa[2]), .A3(n9512), 
        .Y(n5405) );
  INVX1_LVT U6541 ( .A(n1279), .Y(n5168) );
  OA21X1_LVT U6542 ( .A1(n3206), .A2(n5405), .A3(n5168), .Y(n9425) );
  NAND3X0_LVT U6543 ( .A1(io_imem_bht_update_valid), .A2(n5169), .A3(n3251), 
        .Y(n5171) );
  AO22X1_LVT U6544 ( .A1(mem_reg_store), .A2(bpu_io_xcpt_st), .A3(
        bpu_io_xcpt_ld), .A4(mem_reg_load), .Y(n5170) );
  AO22X1_LVT U6545 ( .A1(mem_reg_store), .A2(bpu_io_debug_st), .A3(
        bpu_io_debug_ld), .A4(mem_reg_load), .Y(n9237) );
  OR2X1_LVT U6546 ( .A1(n5170), .A2(n9237), .Y(n5172) );
  OR2X1_LVT U6547 ( .A1(n5171), .A2(n5172), .Y(io_dmem_s1_kill) );
  NOR2X0_LVT U6548 ( .A1(n1281), .A2(io_dmem_s1_kill), .Y(n1829) );
  AO22X1_LVT U6549 ( .A1(io_imem_req_bits_speculative), .A2(n1281), .A3(n5172), 
        .A4(io_imem_bht_update_valid), .Y(N529) );
  AND2X1_LVT U6550 ( .A1(n3198), .A2(n3043), .Y(n5227) );
  AND2X1_LVT U6551 ( .A1(n5227), .A2(n3199), .Y(n5354) );
  AND2X1_LVT U6552 ( .A1(n3103), .A2(n3041), .Y(n5272) );
  AO21X1_LVT U6553 ( .A1(n5175), .A2(wb_ctrl_wfd), .A3(io_fpu_sboard_set), .Y(
        n5176) );
  AO21X1_LVT U6554 ( .A1(n5354), .A2(n5275), .A3(n_T_1298[5]), .Y(n5179) );
  AND3X1_LVT U6555 ( .A1(io_dmem_resp_bits_has_data), .A2(
        io_dmem_resp_bits_tag[0]), .A3(n2030), .Y(io_fpu_dmem_resp_val) );
  NAND2X0_LVT U6556 ( .A1(io_fpu_dmem_resp_val), .A2(io_dmem_resp_bits_replay), 
        .Y(n5191) );
  NAND3X0_LVT U6557 ( .A1(n5254), .A2(n5191), .A3(n5177), .Y(n9379) );
  NAND2X0_LVT U6558 ( .A1(n5183), .A2(io_fpu_sboard_clra[0]), .Y(n5271) );
  OR2X1_LVT U6559 ( .A1(n5257), .A2(n5271), .Y(n5277) );
  OA22X1_LVT U6560 ( .A1(n5277), .A2(n5193), .A3(n5192), .A4(n5276), .Y(n5178)
         );
  AND3X1_LVT U6561 ( .A1(n5179), .A2(n3794), .A3(n5178), .Y(N784) );
  AND2X1_LVT U6562 ( .A1(n3199), .A2(n3102), .Y(n5255) );
  AND2X1_LVT U6563 ( .A1(n5255), .A2(n3198), .Y(n5355) );
  AND2X1_LVT U6564 ( .A1(n3201), .A2(wb_waddr[1]), .Y(n5303) );
  AO21X1_LVT U6565 ( .A1(n5355), .A2(n5248), .A3(n_T_1298[2]), .Y(n5181) );
  AND2X1_LVT U6566 ( .A1(io_fpu_sboard_clr), .A2(io_fpu_sboard_clra[1]), .Y(
        n5190) );
  NAND2X0_LVT U6567 ( .A1(n5190), .A2(n5182), .Y(n5262) );
  OR2X1_LVT U6568 ( .A1(io_fpu_sboard_clra[2]), .A2(n5193), .Y(n5201) );
  OR2X1_LVT U6569 ( .A1(io_fpu_dmem_resp_tag[2]), .A2(n5192), .Y(n5200) );
  OA22X1_LVT U6570 ( .A1(n5262), .A2(n5201), .A3(n5200), .A4(n5261), .Y(n5180)
         );
  AND3X1_LVT U6571 ( .A1(n5181), .A2(n3793), .A3(n5180), .Y(N781) );
  AND2X1_LVT U6572 ( .A1(n3103), .A2(n3201), .Y(n5282) );
  AO21X1_LVT U6573 ( .A1(n5354), .A2(n5265), .A3(n_T_1298[4]), .Y(n5187) );
  NAND2X0_LVT U6574 ( .A1(n5183), .A2(n5182), .Y(n5281) );
  OR2X1_LVT U6575 ( .A1(n5257), .A2(n5281), .Y(n5267) );
  OA22X1_LVT U6576 ( .A1(n5193), .A2(n5267), .A3(n5192), .A4(n5266), .Y(n5186)
         );
  AND3X1_LVT U6577 ( .A1(n5187), .A2(n3793), .A3(n5186), .Y(N783) );
  AO21X1_LVT U6578 ( .A1(n5354), .A2(n5248), .A3(n_T_1298[6]), .Y(n5189) );
  OR2X1_LVT U6579 ( .A1(n5257), .A2(n5262), .Y(n5251) );
  OR2X1_LVT U6580 ( .A1(n5259), .A2(n5261), .Y(n5250) );
  OA22X1_LVT U6581 ( .A1(n5193), .A2(n5251), .A3(n5192), .A4(n5250), .Y(n5188)
         );
  AND3X1_LVT U6582 ( .A1(n5189), .A2(n3794), .A3(n5188), .Y(N785) );
  AND2X1_LVT U6583 ( .A1(n3041), .A2(wb_waddr[1]), .Y(n5298) );
  AO21X1_LVT U6584 ( .A1(n5354), .A2(n5285), .A3(n_T_1298[7]), .Y(n5195) );
  NAND2X0_LVT U6585 ( .A1(n5190), .A2(io_fpu_sboard_clra[0]), .Y(n5295) );
  OR2X1_LVT U6586 ( .A1(n5257), .A2(n5295), .Y(n5288) );
  OR2X1_LVT U6587 ( .A1(n5259), .A2(n5292), .Y(n5286) );
  OA22X1_LVT U6588 ( .A1(n5193), .A2(n5288), .A3(n5192), .A4(n5286), .Y(n5194)
         );
  AND3X1_LVT U6589 ( .A1(n5195), .A2(n3793), .A3(n5194), .Y(N786) );
  AO21X1_LVT U6590 ( .A1(n5355), .A2(n5275), .A3(n_T_1298[1]), .Y(n5197) );
  OA22X1_LVT U6591 ( .A1(n5271), .A2(n5201), .A3(n5200), .A4(n5270), .Y(n5196)
         );
  AND3X1_LVT U6592 ( .A1(n5197), .A2(n3793), .A3(n5196), .Y(N780) );
  AO21X1_LVT U6593 ( .A1(n5355), .A2(n5265), .A3(n_T_1298[0]), .Y(n5199) );
  OA22X1_LVT U6594 ( .A1(n5281), .A2(n5201), .A3(n5200), .A4(n5280), .Y(n5198)
         );
  AND3X1_LVT U6595 ( .A1(n5199), .A2(n3794), .A3(n5198), .Y(N779) );
  AO21X1_LVT U6596 ( .A1(n5355), .A2(n5285), .A3(n_T_1298[3]), .Y(n5203) );
  OA22X1_LVT U6597 ( .A1(n5295), .A2(n5201), .A3(n5200), .A4(n5292), .Y(n5202)
         );
  AND3X1_LVT U6598 ( .A1(n5203), .A2(n3794), .A3(n5202), .Y(N782) );
  AND2X1_LVT U6599 ( .A1(wb_waddr[4]), .A2(wb_waddr[3]), .Y(n5210) );
  AND2X1_LVT U6600 ( .A1(n5210), .A2(n3102), .Y(n5305) );
  AO21X1_LVT U6601 ( .A1(n5305), .A2(n5248), .A3(n_T_1298[26]), .Y(n5205) );
  AND2X1_LVT U6602 ( .A1(io_fpu_sboard_clra[3]), .A2(io_fpu_sboard_clra[4]), 
        .Y(n5211) );
  NAND2X0_LVT U6603 ( .A1(n5211), .A2(n5257), .Y(n5218) );
  AND2X1_LVT U6604 ( .A1(io_fpu_dmem_resp_tag[3]), .A2(io_fpu_dmem_resp_tag[4]), .Y(n5212) );
  NAND2X0_LVT U6605 ( .A1(n5212), .A2(n5259), .Y(n5217) );
  OA22X1_LVT U6606 ( .A1(n5262), .A2(n5218), .A3(n5217), .A4(n5261), .Y(n5204)
         );
  AND3X1_LVT U6607 ( .A1(n5205), .A2(n3794), .A3(n5204), .Y(N805) );
  AO21X1_LVT U6608 ( .A1(n5305), .A2(n5275), .A3(n_T_1298[25]), .Y(n5207) );
  OA22X1_LVT U6609 ( .A1(n5271), .A2(n5218), .A3(n5217), .A4(n5270), .Y(n5206)
         );
  AND3X1_LVT U6610 ( .A1(n5207), .A2(n3794), .A3(n5206), .Y(N804) );
  AO21X1_LVT U6611 ( .A1(n5305), .A2(n5285), .A3(n_T_1298[27]), .Y(n5209) );
  OA22X1_LVT U6612 ( .A1(n5295), .A2(n5218), .A3(n5217), .A4(n5292), .Y(n5208)
         );
  AND3X1_LVT U6613 ( .A1(n5209), .A2(n3794), .A3(n5208), .Y(N806) );
  AO21X1_LVT U6614 ( .A1(n5317), .A2(n5248), .A3(n_T_1298[30]), .Y(n5214) );
  INVX1_LVT U6615 ( .A(n5211), .Y(n5224) );
  INVX1_LVT U6616 ( .A(n5212), .Y(n5223) );
  OA22X1_LVT U6617 ( .A1(n5251), .A2(n5224), .A3(n5223), .A4(n5250), .Y(n5213)
         );
  AND3X1_LVT U6618 ( .A1(n5214), .A2(n3794), .A3(n5213), .Y(N809) );
  AO21X1_LVT U6619 ( .A1(n5317), .A2(n5275), .A3(n_T_1298[29]), .Y(n5216) );
  OA22X1_LVT U6620 ( .A1(n5277), .A2(n5224), .A3(n5223), .A4(n5276), .Y(n5215)
         );
  AND3X1_LVT U6621 ( .A1(n5216), .A2(n3794), .A3(n5215), .Y(N808) );
  AO21X1_LVT U6622 ( .A1(n5305), .A2(n5265), .A3(n_T_1298[24]), .Y(n5220) );
  OA22X1_LVT U6623 ( .A1(n5281), .A2(n5218), .A3(n5217), .A4(n5280), .Y(n5219)
         );
  AND3X1_LVT U6624 ( .A1(n5220), .A2(n3794), .A3(n5219), .Y(N803) );
  AO21X1_LVT U6625 ( .A1(n5317), .A2(n5265), .A3(n_T_1298[28]), .Y(n5222) );
  OA22X1_LVT U6626 ( .A1(n5267), .A2(n5224), .A3(n5223), .A4(n5266), .Y(n5221)
         );
  AND3X1_LVT U6627 ( .A1(n5222), .A2(n3794), .A3(n5221), .Y(N807) );
  AO21X1_LVT U6628 ( .A1(n5317), .A2(n5285), .A3(n_T_1298[31]), .Y(n5226) );
  OA22X1_LVT U6629 ( .A1(n5288), .A2(n5224), .A3(n5223), .A4(n5286), .Y(n5225)
         );
  AND3X1_LVT U6630 ( .A1(n5226), .A2(n3794), .A3(n5225), .Y(N810) );
  AO21X1_LVT U6631 ( .A1(n5382), .A2(n5285), .A3(n_T_1298[15]), .Y(n5230) );
  NAND2X0_LVT U6632 ( .A1(n5228), .A2(io_fpu_dmem_resp_tag[3]), .Y(n5244) );
  OA22X1_LVT U6633 ( .A1(n5245), .A2(n5288), .A3(n5244), .A4(n5286), .Y(n5229)
         );
  AND3X1_LVT U6634 ( .A1(n5230), .A2(n3794), .A3(n5229), .Y(N794) );
  AO21X1_LVT U6635 ( .A1(n5382), .A2(n5248), .A3(n_T_1298[14]), .Y(n5232) );
  OA22X1_LVT U6636 ( .A1(n5245), .A2(n5251), .A3(n5244), .A4(n5250), .Y(n5231)
         );
  AND3X1_LVT U6637 ( .A1(n5232), .A2(n3794), .A3(n5231), .Y(N793) );
  OR2X1_LVT U6638 ( .A1(io_fpu_sboard_clra[2]), .A2(n5245), .Y(n5238) );
  NAND3X0_LVT U6639 ( .A1(n3198), .A2(n3102), .A3(wb_waddr[3]), .Y(n5359) );
  NOR3X0_LVT U6640 ( .A1(reset), .A2(n5359), .A3(n5254), .Y(n5239) );
  OA22X1_LVT U6641 ( .A1(n5238), .A2(n5262), .A3(n5237), .A4(n5261), .Y(n5234)
         );
  AO22X1_LVT U6642 ( .A1(n5239), .A2(n5303), .A3(n_T_1298[10]), .A4(n3793), 
        .Y(n5233) );
  AND2X1_LVT U6643 ( .A1(n5234), .A2(n5233), .Y(N789) );
  OA22X1_LVT U6644 ( .A1(n5238), .A2(n5281), .A3(n5237), .A4(n5280), .Y(n5236)
         );
  AO22X1_LVT U6645 ( .A1(n5239), .A2(n5282), .A3(n_T_1298[8]), .A4(n3793), .Y(
        n5235) );
  AND2X1_LVT U6646 ( .A1(n5236), .A2(n5235), .Y(N787) );
  OA22X1_LVT U6647 ( .A1(n5238), .A2(n5271), .A3(n5237), .A4(n5270), .Y(n5241)
         );
  AO22X1_LVT U6648 ( .A1(n5239), .A2(n5272), .A3(n_T_1298[9]), .A4(n3793), .Y(
        n5240) );
  AND2X1_LVT U6649 ( .A1(n5241), .A2(n5240), .Y(N788) );
  AO21X1_LVT U6650 ( .A1(n5382), .A2(n5265), .A3(n_T_1298[12]), .Y(n5243) );
  OA22X1_LVT U6651 ( .A1(n5245), .A2(n5267), .A3(n5244), .A4(n5266), .Y(n5242)
         );
  AND3X1_LVT U6652 ( .A1(n5243), .A2(n5296), .A3(n5242), .Y(N791) );
  AO21X1_LVT U6653 ( .A1(n5382), .A2(n5275), .A3(n_T_1298[13]), .Y(n5247) );
  OA22X1_LVT U6654 ( .A1(n5245), .A2(n5277), .A3(n5244), .A4(n5276), .Y(n5246)
         );
  AND3X1_LVT U6655 ( .A1(n5247), .A2(n5296), .A3(n5246), .Y(N792) );
  AND3X1_LVT U6656 ( .A1(n3199), .A2(n3043), .A3(wb_waddr[4]), .Y(n5325) );
  AO21X1_LVT U6657 ( .A1(n5325), .A2(n5248), .A3(n_T_1298[22]), .Y(n5253) );
  INVX1_LVT U6658 ( .A(n5258), .Y(n5289) );
  AND2X1_LVT U6659 ( .A1(n5249), .A2(io_fpu_dmem_resp_tag[4]), .Y(n5260) );
  OA22X1_LVT U6660 ( .A1(n5289), .A2(n5251), .A3(n5287), .A4(n5250), .Y(n5252)
         );
  AND3X1_LVT U6661 ( .A1(n5253), .A2(n5296), .A3(n5252), .Y(N801) );
  AND2X1_LVT U6662 ( .A1(n5255), .A2(wb_waddr[4]), .Y(n5326) );
  AND3X1_LVT U6663 ( .A1(n5256), .A2(n5326), .A3(n4498), .Y(n5297) );
  AO22X1_LVT U6664 ( .A1(n5303), .A2(n5297), .A3(n3793), .A4(n_T_1298[18]), 
        .Y(n5264) );
  NAND2X0_LVT U6665 ( .A1(n5258), .A2(n5257), .Y(n5294) );
  NAND2X0_LVT U6666 ( .A1(n5260), .A2(n5259), .Y(n5293) );
  OA22X1_LVT U6667 ( .A1(n5262), .A2(n5294), .A3(n5293), .A4(n5261), .Y(n5263)
         );
  AND2X1_LVT U6668 ( .A1(n5264), .A2(n5263), .Y(N797) );
  AO21X1_LVT U6669 ( .A1(n5325), .A2(n5265), .A3(n_T_1298[20]), .Y(n5269) );
  OA22X1_LVT U6670 ( .A1(n5289), .A2(n5267), .A3(n5287), .A4(n5266), .Y(n5268)
         );
  AND3X1_LVT U6671 ( .A1(n5269), .A2(n5296), .A3(n5268), .Y(N799) );
  OA22X1_LVT U6672 ( .A1(n5271), .A2(n5294), .A3(n5293), .A4(n5270), .Y(n5274)
         );
  AO22X1_LVT U6673 ( .A1(n5272), .A2(n5297), .A3(n3793), .A4(n_T_1298[17]), 
        .Y(n5273) );
  AND2X1_LVT U6674 ( .A1(n5274), .A2(n5273), .Y(N796) );
  AO21X1_LVT U6675 ( .A1(n5325), .A2(n5275), .A3(n_T_1298[21]), .Y(n5279) );
  OA22X1_LVT U6676 ( .A1(n5289), .A2(n5277), .A3(n5287), .A4(n5276), .Y(n5278)
         );
  AND3X1_LVT U6677 ( .A1(n5279), .A2(n5296), .A3(n5278), .Y(N800) );
  OA22X1_LVT U6678 ( .A1(n5281), .A2(n5294), .A3(n5293), .A4(n5280), .Y(n5284)
         );
  AO22X1_LVT U6679 ( .A1(n5282), .A2(n5297), .A3(n3793), .A4(n_T_1298[16]), 
        .Y(n5283) );
  AND2X1_LVT U6680 ( .A1(n5284), .A2(n5283), .Y(N795) );
  AO21X1_LVT U6681 ( .A1(n5325), .A2(n5285), .A3(n_T_1298[23]), .Y(n5291) );
  OA22X1_LVT U6682 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .Y(n5290)
         );
  AND3X1_LVT U6683 ( .A1(n5291), .A2(n3793), .A3(n5290), .Y(N802) );
  OA22X1_LVT U6684 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .Y(n5300)
         );
  AO22X1_LVT U6685 ( .A1(n5298), .A2(n5297), .A3(n3793), .A4(n_T_1298[19]), 
        .Y(n5299) );
  AND2X1_LVT U6686 ( .A1(n5300), .A2(n5299), .Y(N798) );
  AND2X1_LVT U6687 ( .A1(n5301), .A2(csr_io_retire), .Y(n9380) );
  NAND2X0_LVT U6688 ( .A1(n3046), .A2(n4498), .Y(n5302) );
  AND2X1_LVT U6689 ( .A1(n5304), .A2(n5303), .Y(n5374) );
  NAND2X0_LVT U6690 ( .A1(n5378), .A2(n5305), .Y(n5310) );
  NAND2X0_LVT U6691 ( .A1(n5307), .A2(n5335), .Y(n5308) );
  NAND3X0_LVT U6692 ( .A1(n5308), .A2(n2572), .A3(n_T_1187[27]), .Y(n5309) );
  AND2X1_LVT U6693 ( .A1(n5379), .A2(n5313), .Y(n5367) );
  AND2X1_LVT U6694 ( .A1(n5339), .A2(n3046), .Y(n5363) );
  AND2X1_LVT U6695 ( .A1(n5313), .A2(n5363), .Y(n5385) );
  AND2X1_LVT U6696 ( .A1(n_T_1187[30]), .A2(n2572), .Y(n5312) );
  AND2X1_LVT U6697 ( .A1(n5356), .A2(n3046), .Y(n5390) );
  AND2X1_LVT U6698 ( .A1(n5313), .A2(n5390), .Y(n5371) );
  NAND2X0_LVT U6699 ( .A1(n5371), .A2(n5314), .Y(n5311) );
  AO22X1_LVT U6700 ( .A1(n5317), .A2(n5374), .A3(n5312), .A4(n5311), .Y(N776)
         );
  AND2X1_LVT U6701 ( .A1(n_T_1187[31]), .A2(n2572), .Y(n5316) );
  AND2X1_LVT U6702 ( .A1(n5335), .A2(n3046), .Y(n5360) );
  AND2X1_LVT U6703 ( .A1(n5360), .A2(n5313), .Y(n5375) );
  NAND2X0_LVT U6704 ( .A1(n5375), .A2(n5314), .Y(n5315) );
  AO22X1_LVT U6705 ( .A1(n5378), .A2(n5317), .A3(n5316), .A4(n5315), .Y(N777)
         );
  NAND2X0_LVT U6706 ( .A1(n5366), .A2(n5325), .Y(n5320) );
  NAND2X0_LVT U6707 ( .A1(n5367), .A2(n5328), .Y(n5318) );
  NAND3X0_LVT U6708 ( .A1(n5318), .A2(n_T_1187[20]), .A3(n2572), .Y(n5319) );
  NAND2X0_LVT U6709 ( .A1(n5320), .A2(n5319), .Y(N766) );
  AND2X1_LVT U6710 ( .A1(n_T_1187[22]), .A2(n2572), .Y(n5322) );
  NAND2X0_LVT U6711 ( .A1(n5371), .A2(n5328), .Y(n5321) );
  AO22X1_LVT U6712 ( .A1(n5325), .A2(n5374), .A3(n5322), .A4(n5321), .Y(N768)
         );
  AND2X1_LVT U6713 ( .A1(n_T_1187[23]), .A2(n2572), .Y(n5324) );
  NAND2X0_LVT U6714 ( .A1(n5375), .A2(n5328), .Y(n5323) );
  AO22X1_LVT U6715 ( .A1(n5378), .A2(n5325), .A3(n5324), .A4(n5323), .Y(N769)
         );
  AND2X1_LVT U6716 ( .A1(n5328), .A2(n2575), .Y(n5332) );
  AO21X1_LVT U6717 ( .A1(n5360), .A2(n5332), .A3(n3258), .Y(n5329) );
  OAI22X1_LVT U6718 ( .A1(n5334), .A2(n5362), .A3(n5329), .A4(n3185), .Y(N765)
         );
  AO21X1_LVT U6719 ( .A1(n5363), .A2(n5332), .A3(n3113), .Y(n5330) );
  OAI22X1_LVT U6720 ( .A1(n5334), .A2(n5365), .A3(n5330), .A4(n3185), .Y(N763)
         );
  AO21X1_LVT U6721 ( .A1(n5379), .A2(n5332), .A3(n3261), .Y(n5331) );
  OAI22X1_LVT U6722 ( .A1(n5381), .A2(n5334), .A3(n5331), .A4(n3185), .Y(N762)
         );
  AO21X1_LVT U6723 ( .A1(n5390), .A2(n5332), .A3(n3263), .Y(n5333) );
  OAI22X1_LVT U6724 ( .A1(n5334), .A2(n5392), .A3(n5333), .A4(n3185), .Y(N764)
         );
  NAND2X0_LVT U6725 ( .A1(n5378), .A2(n5355), .Y(n5338) );
  AND2X1_LVT U6726 ( .A1(n5426), .A2(n5428), .Y(n5351) );
  NAND2X0_LVT U6727 ( .A1(n5357), .A2(n5335), .Y(n5336) );
  NAND3X0_LVT U6728 ( .A1(n2572), .A2(n_T_1187[3]), .A3(n5336), .Y(n5337) );
  NAND2X0_LVT U6729 ( .A1(n5338), .A2(n5337), .Y(N749) );
  NAND2X0_LVT U6730 ( .A1(n5383), .A2(n5355), .Y(n5342) );
  NAND2X0_LVT U6731 ( .A1(n5357), .A2(n5339), .Y(n5340) );
  NAND3X0_LVT U6732 ( .A1(n2572), .A2(n_T_1187[1]), .A3(n5340), .Y(n5341) );
  NAND2X0_LVT U6733 ( .A1(n5342), .A2(n5341), .Y(N747) );
  NAND2X0_LVT U6734 ( .A1(n5383), .A2(n5354), .Y(n5345) );
  NAND2X0_LVT U6735 ( .A1(n5385), .A2(n5351), .Y(n5343) );
  NAND3X0_LVT U6736 ( .A1(n5343), .A2(n_T_1187[5]), .A3(n2572), .Y(n5344) );
  NAND2X0_LVT U6737 ( .A1(n5345), .A2(n5344), .Y(N751) );
  AND2X1_LVT U6738 ( .A1(n_T_1187[6]), .A2(n2572), .Y(n5347) );
  NAND2X0_LVT U6739 ( .A1(n5371), .A2(n5351), .Y(n5346) );
  AO22X1_LVT U6740 ( .A1(n5354), .A2(n5374), .A3(n5347), .A4(n5346), .Y(N752)
         );
  NAND2X0_LVT U6741 ( .A1(n5366), .A2(n5354), .Y(n5350) );
  NAND2X0_LVT U6742 ( .A1(n5367), .A2(n5351), .Y(n5348) );
  NAND3X0_LVT U6743 ( .A1(n5348), .A2(n_T_1187[4]), .A3(n2572), .Y(n5349) );
  NAND2X0_LVT U6744 ( .A1(n5350), .A2(n5349), .Y(N750) );
  AND2X1_LVT U6745 ( .A1(n_T_1187[7]), .A2(n2572), .Y(n5353) );
  NAND2X0_LVT U6746 ( .A1(n5375), .A2(n5351), .Y(n5352) );
  AO22X1_LVT U6747 ( .A1(n5378), .A2(n5354), .A3(n5353), .A4(n5352), .Y(N753)
         );
  AND2X1_LVT U6748 ( .A1(n5384), .A2(n2575), .Y(n5389) );
  AO21X1_LVT U6749 ( .A1(n5360), .A2(n5389), .A3(n3259), .Y(n5361) );
  OAI22X1_LVT U6750 ( .A1(n5393), .A2(n5362), .A3(n5361), .A4(n3185), .Y(N757)
         );
  AO21X1_LVT U6751 ( .A1(n5363), .A2(n5389), .A3(n3133), .Y(n5364) );
  OAI22X1_LVT U6752 ( .A1(n5393), .A2(n5365), .A3(n5364), .A4(n3185), .Y(N755)
         );
  NAND2X0_LVT U6753 ( .A1(n5366), .A2(n5382), .Y(n5370) );
  NAND2X0_LVT U6754 ( .A1(n5367), .A2(n5384), .Y(n5368) );
  NAND3X0_LVT U6755 ( .A1(n5368), .A2(n_T_1187[12]), .A3(n2572), .Y(n5369) );
  NAND2X0_LVT U6756 ( .A1(n5370), .A2(n5369), .Y(N758) );
  AND2X1_LVT U6757 ( .A1(n_T_1187[14]), .A2(n2572), .Y(n5373) );
  NAND2X0_LVT U6758 ( .A1(n5371), .A2(n5384), .Y(n5372) );
  AO22X1_LVT U6759 ( .A1(n5382), .A2(n5374), .A3(n5373), .A4(n5372), .Y(N760)
         );
  AND2X1_LVT U6760 ( .A1(n_T_1187[15]), .A2(n2572), .Y(n5377) );
  NAND2X0_LVT U6761 ( .A1(n5375), .A2(n5384), .Y(n5376) );
  AO22X1_LVT U6762 ( .A1(n5378), .A2(n5382), .A3(n5377), .A4(n5376), .Y(N761)
         );
  AO21X1_LVT U6763 ( .A1(n5379), .A2(n5389), .A3(n3134), .Y(n5380) );
  OAI22X1_LVT U6764 ( .A1(n5381), .A2(n5393), .A3(n5380), .A4(n3185), .Y(N754)
         );
  NAND2X0_LVT U6765 ( .A1(n5383), .A2(n5382), .Y(n5388) );
  NAND2X0_LVT U6766 ( .A1(n5385), .A2(n5384), .Y(n5386) );
  NAND3X0_LVT U6767 ( .A1(n5386), .A2(n_T_1187[13]), .A3(n2572), .Y(n5387) );
  NAND2X0_LVT U6768 ( .A1(n5388), .A2(n5387), .Y(N759) );
  AO21X1_LVT U6769 ( .A1(n5390), .A2(n5389), .A3(n3129), .Y(n5391) );
  OAI22X1_LVT U6770 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n3185), .Y(N756)
         );
  NOR3X0_LVT U6771 ( .A1(io_fpu_inst[23]), .A2(n5394), .A3(io_fpu_inst[22]), 
        .Y(n5395) );
  INVX1_LVT U6772 ( .A(io_dmem_perf_release), .Y(n5399) );
  OR3X1_LVT U6773 ( .A1(csr_io_time[0]), .A2(csr_io_time[4]), .A3(
        csr_io_time[3]), .Y(n5397) );
  OR3X1_LVT U6774 ( .A1(csr_io_time[1]), .A2(csr_io_time[2]), .A3(n5397), .Y(
        n5398) );
  AND3X1_LVT U6775 ( .A1(n9418), .A2(n5399), .A3(n5398), .Y(n5400) );
  OA21X1_LVT U6776 ( .A1(id_reg_pause), .A2(n5401), .A3(n5400), .Y(n1820) );
  NAND3X0_LVT U6777 ( .A1(io_imem_bht_update_valid), .A2(n3251), .A3(n5404), 
        .Y(io_fpu_killm) );
  AND2X1_LVT U6778 ( .A1(io_fpu_killm), .A2(n_T_1057), .Y(div_io_kill) );
  NAND2X0_LVT U6779 ( .A1(n5419), .A2(n5421), .Y(n5480) );
  OR2X1_LVT U6780 ( .A1(n5420), .A2(n5480), .Y(do_bypass_1) );
  INVX1_LVT U6781 ( .A(n5409), .Y(n5407) );
  AND2X1_LVT U6782 ( .A1(mem_ctrl_wxd), .A2(n2492), .Y(n5408) );
  AO222X1_LVT U6783 ( .A1(n6249), .A2(mem_br_target[0]), .A3(n6855), .A4(
        n_T_918[0]), .A5(io_fpu_toint_data[0]), .A6(n6856), .Y(N598) );
  AND2X1_LVT U6784 ( .A1(n5414), .A2(n5413), .Y(n5416) );
  AO22X1_LVT U6785 ( .A1(n6860), .A2(io_dmem_resp_bits_data[0]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[0]), .Y(n5417) );
  AO21X1_LVT U6786 ( .A1(n3854), .A2(div_io_resp_bits_data[0]), .A3(n5417), 
        .Y(n5418) );
  AO21X1_LVT U6787 ( .A1(n3841), .A2(csr_io_rw_rdata[0]), .A3(n5418), .Y(
        n_T_427__T_1136_data[0]) );
  NAND3X0_LVT U6788 ( .A1(n5420), .A2(n572), .A3(n5419), .Y(n5422) );
  AND2X1_LVT U6789 ( .A1(n5422), .A2(n5421), .Y(n5468) );
  AND2X1_LVT U6790 ( .A1(n5425), .A2(n5424), .Y(n5433) );
  NAND2X0_LVT U6791 ( .A1(n9398), .A2(n9403), .Y(n9386) );
  AND2X1_LVT U6792 ( .A1(n5429), .A2(n9388), .Y(n5430) );
  AND2X1_LVT U6793 ( .A1(n5451), .A2(n2878), .Y(n6795) );
  AND2X1_LVT U6794 ( .A1(n5456), .A2(n2878), .Y(n6869) );
  AND2X1_LVT U6795 ( .A1(n5454), .A2(n2878), .Y(n6715) );
  AO22X1_LVT U6796 ( .A1(n3811), .A2(n_T_427[895]), .A3(n_T_427[640]), .A4(
        n3861), .Y(n5442) );
  AO22X1_LVT U6797 ( .A1(n_T_427[704]), .A2(n3804), .A3(n3860), .A4(
        n_T_427[192]), .Y(n5441) );
  AO22X1_LVT U6798 ( .A1(n_T_427[831]), .A2(n6871), .A3(n3872), .A4(
        n_T_427[256]), .Y(n5440) );
  AO22X1_LVT U6799 ( .A1(n3815), .A2(n_T_427[128]), .A3(n3839), .A4(n_T_427[0]), .Y(n5439) );
  NOR4X1_LVT U6800 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .Y(n5443)
         );
  NAND2X0_LVT U6801 ( .A1(n4318), .A2(n3959), .Y(n5444) );
  AND2X1_LVT U6802 ( .A1(n5446), .A2(n5456), .Y(n6880) );
  AND2X1_LVT U6803 ( .A1(n5446), .A2(n5455), .Y(n6891) );
  INVX1_LVT U6804 ( .A(n5447), .Y(n5448) );
  AND2X1_LVT U6805 ( .A1(n5457), .A2(n5450), .Y(n6893) );
  AO22X1_LVT U6806 ( .A1(n3934), .A2(n_T_427[1407]), .A3(n_T_427[1279]), .A4(
        n3929), .Y(n5461) );
  AND2X1_LVT U6807 ( .A1(n5457), .A2(n5452), .Y(n6895) );
  AO22X1_LVT U6808 ( .A1(n3944), .A2(n_T_427[1151]), .A3(n_T_427[1215]), .A4(
        n3939), .Y(n5460) );
  AND2X1_LVT U6809 ( .A1(n5457), .A2(n5454), .Y(n6897) );
  AO22X1_LVT U6810 ( .A1(n3954), .A2(n_T_427[1087]), .A3(n_T_427[959]), .A4(
        n3949), .Y(n5459) );
  AND2X1_LVT U6811 ( .A1(n5457), .A2(n5456), .Y(n6883) );
  AO22X1_LVT U6812 ( .A1(n3900), .A2(n_T_427[1023]), .A3(n_T_427[64]), .A4(
        n3831), .Y(n5458) );
  NOR4X1_LVT U6813 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .Y(n5462)
         );
  NAND3X0_LVT U6814 ( .A1(n5462), .A2(n5463), .A3(n5464), .Y(n5467) );
  INVX1_LVT U6815 ( .A(do_bypass_1), .Y(n5465) );
  AND2X1_LVT U6816 ( .A1(n5466), .A2(n5465), .Y(n9382) );
  MUX21X1_LVT U6817 ( .A1(n5468), .A2(n5467), .S0(n9382), .Y(N678) );
  AO222X1_LVT U6818 ( .A1(mem_br_target[1]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[1]), .A5(n_T_918[1]), .A6(n6855), .Y(N599) );
  NAND2X0_LVT U6819 ( .A1(csr_io_rw_rdata[1]), .A2(n3844), .Y(n5471) );
  AOI22X1_LVT U6820 ( .A1(n3852), .A2(io_dmem_resp_bits_data[1]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[1]), .Y(n5470) );
  NAND2X0_LVT U6821 ( .A1(div_io_resp_bits_data[1]), .A2(n3857), .Y(n5469) );
  NAND3X0_LVT U6822 ( .A1(n5471), .A2(n5470), .A3(n5469), .Y(
        n_T_427__T_1136_data[1]) );
  AO22X1_LVT U6823 ( .A1(n_T_427[896]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[449]), .Y(n5478) );
  AO22X1_LVT U6824 ( .A1(n3815), .A2(n_T_427[129]), .A3(n3871), .A4(
        n_T_427[257]), .Y(n5477) );
  AOI22X1_LVT U6825 ( .A1(n3797), .A2(n_T_427[577]), .A3(n3867), .A4(
        n_T_427[321]), .Y(n5475) );
  AOI22X1_LVT U6826 ( .A1(n6765), .A2(n_T_427[705]), .A3(n3859), .A4(
        n_T_427[193]), .Y(n5474) );
  AOI22X1_LVT U6827 ( .A1(n_T_427[641]), .A2(n3861), .A3(n3868), .A4(
        n_T_427[513]), .Y(n5473) );
  NAND2X0_LVT U6828 ( .A1(n3840), .A2(n_T_427[1]), .Y(n5472) );
  NAND4X0_LVT U6829 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .Y(n5476) );
  OR3X1_LVT U6830 ( .A1(n5478), .A2(n5477), .A3(n5476), .Y(n5479) );
  NAND2X0_LVT U6831 ( .A1(n_T_918[0]), .A2(n6899), .Y(n9125) );
  AND2X1_LVT U6832 ( .A1(n594), .A2(n_T_635[1]), .Y(n5484) );
  NAND2X0_LVT U6833 ( .A1(io_imem_sfence_bits_addr[0]), .A2(n6900), .Y(n9124)
         );
  OR2X1_LVT U6834 ( .A1(ex_reg_rs_bypass_1), .A2(n594), .Y(n9123) );
  INVX1_LVT U6835 ( .A(n5483), .Y(n9120) );
  NAND2X0_LVT U6836 ( .A1(n9120), .A2(io_fpu_dmem_resp_data[0]), .Y(n5482) );
  NAND4X0_LVT U6837 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n5482), .Y(
        n_T_702[0]) );
  NAND2X0_LVT U6838 ( .A1(n_T_918[1]), .A2(n6899), .Y(n9137) );
  NAND2X0_LVT U6839 ( .A1(n_T_635[1]), .A2(n3243), .Y(n9135) );
  NAND2X0_LVT U6840 ( .A1(io_imem_sfence_bits_addr[1]), .A2(n5484), .Y(n9136)
         );
  AO222X1_LVT U6841 ( .A1(mem_br_target[2]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[2]), .A5(n_T_918[2]), .A6(n6855), .Y(N600) );
  AO22X1_LVT U6842 ( .A1(n6860), .A2(io_dmem_resp_bits_data[2]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[2]), .Y(n5485) );
  AO21X1_LVT U6843 ( .A1(n3854), .A2(div_io_resp_bits_data[2]), .A3(n5485), 
        .Y(n5486) );
  NAND2X0_LVT U6844 ( .A1(n4324), .A2(n3958), .Y(n5503) );
  AO22X1_LVT U6845 ( .A1(n3899), .A2(n_T_427[1025]), .A3(n_T_427[194]), .A4(
        n2830), .Y(n5490) );
  AO22X1_LVT U6846 ( .A1(n3832), .A2(n_T_427[66]), .A3(n_T_427[897]), .A4(
        n3896), .Y(n5489) );
  AO22X1_LVT U6847 ( .A1(n2864), .A2(n_T_427[386]), .A3(n_T_427[706]), .A4(
        n3904), .Y(n5488) );
  AO22X1_LVT U6848 ( .A1(n2833), .A2(n_T_427[833]), .A3(n_T_427[2]), .A4(n3913), .Y(n5487) );
  NOR4X1_LVT U6849 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .Y(n5502)
         );
  AOI22X1_LVT U6850 ( .A1(n3838), .A2(n_T_427[450]), .A3(n3871), .A4(
        n_T_427[258]), .Y(n5494) );
  AOI22X1_LVT U6851 ( .A1(n3870), .A2(n_T_427[514]), .A3(n_T_427[578]), .A4(
        n3795), .Y(n5493) );
  OA22X1_LVT U6852 ( .A1(n3519), .A2(n6766), .A3(n3173), .A4(n3083), .Y(n5492)
         );
  AOI22X1_LVT U6853 ( .A1(n3816), .A2(n_T_427[130]), .A3(n_T_427[769]), .A4(
        n3812), .Y(n5491) );
  NAND4X0_LVT U6854 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .Y(n5495) );
  AO22X1_LVT U6855 ( .A1(n3923), .A2(n_T_427[1473]), .A3(n_T_427[1345]), .A4(
        n3917), .Y(n5499) );
  AO22X1_LVT U6856 ( .A1(n3933), .A2(n_T_427[1409]), .A3(n_T_427[1281]), .A4(
        n3927), .Y(n5498) );
  AO22X1_LVT U6857 ( .A1(n3943), .A2(n_T_427[1153]), .A3(n_T_427[1217]), .A4(
        n3937), .Y(n5497) );
  AO22X1_LVT U6858 ( .A1(n3953), .A2(n_T_427[1089]), .A3(n_T_427[961]), .A4(
        n3947), .Y(n5496) );
  NOR4X1_LVT U6859 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .Y(n5500)
         );
  NAND4X0_LVT U6860 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .Y(
        id_rs_1[2]) );
  NAND2X0_LVT U6861 ( .A1(n_T_918[2]), .A2(n6899), .Y(n9150) );
  NAND2X0_LVT U6862 ( .A1(n_T_635[2]), .A2(n6901), .Y(n9149) );
  NAND2X0_LVT U6863 ( .A1(io_imem_sfence_bits_addr[2]), .A2(n6900), .Y(n9148)
         );
  AO222X1_LVT U6864 ( .A1(mem_br_target[3]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[3]), .A5(n_T_918[3]), .A6(n6855), .Y(N601) );
  AO22X1_LVT U6865 ( .A1(n6860), .A2(io_dmem_resp_bits_data[3]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[3]), .Y(n5504) );
  AO21X1_LVT U6866 ( .A1(n3854), .A2(div_io_resp_bits_data[3]), .A3(n5504), 
        .Y(n5505) );
  AO22X1_LVT U6867 ( .A1(n3830), .A2(n_T_427[1793]), .A3(n_T_427[1666]), .A4(
        n3826), .Y(n5509) );
  AO22X1_LVT U6868 ( .A1(n3891), .A2(n_T_427[1538]), .A3(n_T_427[1602]), .A4(
        n3885), .Y(n5508) );
  AO22X1_LVT U6869 ( .A1(n3923), .A2(n_T_427[1474]), .A3(n_T_427[1346]), .A4(
        n3917), .Y(n5507) );
  AO22X1_LVT U6870 ( .A1(n3933), .A2(n_T_427[1410]), .A3(n_T_427[1282]), .A4(
        n3927), .Y(n5506) );
  NOR4X1_LVT U6871 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .Y(n5527)
         );
  AO22X1_LVT U6872 ( .A1(n3943), .A2(n_T_427[1154]), .A3(n_T_427[1218]), .A4(
        n3937), .Y(n5513) );
  AO22X1_LVT U6873 ( .A1(n3953), .A2(n_T_427[1090]), .A3(n_T_427[962]), .A4(
        n3947), .Y(n5512) );
  AO22X1_LVT U6874 ( .A1(n3899), .A2(n_T_427[1026]), .A3(n_T_427[898]), .A4(
        n2831), .Y(n5511) );
  AO22X1_LVT U6875 ( .A1(n3834), .A2(n_T_427[387]), .A3(n_T_427[67]), .A4(
        n3831), .Y(n5510) );
  NOR4X1_LVT U6876 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .Y(n5526)
         );
  AO22X1_LVT U6877 ( .A1(n3907), .A2(n_T_427[770]), .A3(n_T_427[451]), .A4(
        n2824), .Y(n5515) );
  AO22X1_LVT U6878 ( .A1(n2826), .A2(n_T_427[3]), .A3(n_T_427[643]), .A4(n3821), .Y(n5514) );
  AO22X1_LVT U6879 ( .A1(n6796), .A2(n_T_427[131]), .A3(n_T_427[834]), .A4(
        n3875), .Y(n5519) );
  AO22X1_LVT U6880 ( .A1(n6765), .A2(n_T_427[707]), .A3(n3859), .A4(
        n_T_427[195]), .Y(n5518) );
  AO22X1_LVT U6881 ( .A1(n_T_427[515]), .A2(n3868), .A3(n6868), .A4(
        n_T_427[323]), .Y(n5517) );
  AO22X1_LVT U6882 ( .A1(n_T_427[579]), .A2(n3796), .A3(n3871), .A4(
        n_T_427[259]), .Y(n5516) );
  NOR4X1_LVT U6883 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .Y(n5520)
         );
  AOI22X1_LVT U6884 ( .A1(n6764), .A2(n_T_427[1849]), .A3(n_T_427[1730]), .A4(
        n2866), .Y(n5522) );
  NAND2X0_LVT U6885 ( .A1(n4327), .A2(n3957), .Y(n5521) );
  AND3X1_LVT U6886 ( .A1(n5523), .A2(n5522), .A3(n5521), .Y(n5524) );
  NAND4X0_LVT U6887 ( .A1(n5527), .A2(n5524), .A3(n5525), .A4(n5526), .Y(
        id_rs_1[3]) );
  NAND2X0_LVT U6888 ( .A1(n_T_918[3]), .A2(n6899), .Y(n9157) );
  NAND2X0_LVT U6889 ( .A1(n_T_635[3]), .A2(n3243), .Y(n9156) );
  NAND2X0_LVT U6890 ( .A1(io_imem_sfence_bits_addr[3]), .A2(n6900), .Y(n9155)
         );
  AO222X1_LVT U6891 ( .A1(mem_br_target[4]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[4]), .A5(n_T_918[4]), .A6(n6855), .Y(N602) );
  AO22X1_LVT U6892 ( .A1(n6860), .A2(io_dmem_resp_bits_data[4]), .A3(n3847), 
        .A4(io_imem_sfence_bits_addr[4]), .Y(n5528) );
  AO21X1_LVT U6893 ( .A1(n3854), .A2(div_io_resp_bits_data[4]), .A3(n5528), 
        .Y(n5529) );
  AOI22X1_LVT U6894 ( .A1(n6765), .A2(n_T_427[708]), .A3(n3859), .A4(
        n_T_427[196]), .Y(n5533) );
  AOI22X1_LVT U6895 ( .A1(n6871), .A2(n_T_427[835]), .A3(n3871), .A4(
        n_T_427[260]), .Y(n5532) );
  OA22X1_LVT U6896 ( .A1(n3520), .A2(n6766), .A3(n3174), .A4(n3083), .Y(n5531)
         );
  AOI22X1_LVT U6897 ( .A1(n_T_427[899]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[580]), .Y(n5530) );
  NAND4X0_LVT U6898 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .Y(n5534) );
  NAND2X0_LVT U6899 ( .A1(n_T_918[4]), .A2(n6899), .Y(n9161) );
  NAND2X0_LVT U6900 ( .A1(n_T_635[4]), .A2(n6901), .Y(n9160) );
  NAND2X0_LVT U6901 ( .A1(io_imem_sfence_bits_addr[4]), .A2(n6900), .Y(n9159)
         );
  AO222X1_LVT U6902 ( .A1(mem_br_target[5]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[5]), .A5(n_T_918[5]), .A6(n6855), .Y(N603) );
  AO22X1_LVT U6903 ( .A1(n6860), .A2(io_dmem_resp_bits_data[5]), .A3(n3847), 
        .A4(io_imem_sfence_bits_addr[5]), .Y(n5535) );
  AO21X1_LVT U6904 ( .A1(n3854), .A2(div_io_resp_bits_data[5]), .A3(n5535), 
        .Y(n5536) );
  NAND2X0_LVT U6905 ( .A1(n4333), .A2(n3958), .Y(n5554) );
  AO22X1_LVT U6906 ( .A1(n3923), .A2(n_T_427[1476]), .A3(n_T_427[1348]), .A4(
        n3917), .Y(n5540) );
  AO22X1_LVT U6907 ( .A1(n3933), .A2(n_T_427[1412]), .A3(n_T_427[1284]), .A4(
        n3927), .Y(n5539) );
  AO22X1_LVT U6908 ( .A1(n3943), .A2(n_T_427[1156]), .A3(n_T_427[1220]), .A4(
        n3937), .Y(n5538) );
  AO22X1_LVT U6909 ( .A1(n3953), .A2(n_T_427[1092]), .A3(n_T_427[964]), .A4(
        n3947), .Y(n5537) );
  NOR4X1_LVT U6910 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .Y(n5553)
         );
  AOI22X1_LVT U6911 ( .A1(n3797), .A2(n_T_427[581]), .A3(n3867), .A4(
        n_T_427[325]), .Y(n5544) );
  AOI22X1_LVT U6912 ( .A1(n6765), .A2(n_T_427[709]), .A3(n3864), .A4(
        n_T_427[69]), .Y(n5543) );
  AOI22X1_LVT U6913 ( .A1(n3838), .A2(n_T_427[453]), .A3(n_T_427[836]), .A4(
        n3875), .Y(n5542) );
  AOI22X1_LVT U6914 ( .A1(n3863), .A2(n_T_427[645]), .A3(n3865), .A4(
        n_T_427[389]), .Y(n5541) );
  NAND4X0_LVT U6915 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .Y(n5545) );
  AO22X1_LVT U6916 ( .A1(n3899), .A2(n_T_427[1028]), .A3(n_T_427[197]), .A4(
        n2830), .Y(n5550) );
  AO22X1_LVT U6917 ( .A1(n2861), .A2(n_T_427[772]), .A3(n_T_427[900]), .A4(
        n3896), .Y(n5549) );
  AO22X1_LVT U6918 ( .A1(n2826), .A2(n_T_427[5]), .A3(n_T_427[133]), .A4(n3908), .Y(n5548) );
  AO22X1_LVT U6919 ( .A1(n3819), .A2(n_T_427[517]), .A3(n_T_427[261]), .A4(
        n2828), .Y(n5547) );
  NOR4X1_LVT U6920 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .Y(n5551)
         );
  NAND4X0_LVT U6921 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .Y(
        id_rs_1[5]) );
  NAND2X0_LVT U6922 ( .A1(io_fpu_dmem_resp_data[5]), .A2(n9165), .Y(n5558) );
  NAND2X0_LVT U6923 ( .A1(n_T_918[5]), .A2(n6899), .Y(n5557) );
  NAND2X0_LVT U6924 ( .A1(io_imem_sfence_bits_addr[5]), .A2(n6900), .Y(n5556)
         );
  NAND2X0_LVT U6925 ( .A1(n_T_635[5]), .A2(n3243), .Y(n5555) );
  NAND4X0_LVT U6926 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .Y(
        n_T_702[5]) );
  AO222X1_LVT U6927 ( .A1(mem_br_target[6]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[6]), .A5(n6855), .A6(n_T_918[6]), .Y(N604) );
  AO22X1_LVT U6928 ( .A1(n6860), .A2(io_dmem_resp_bits_data[6]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[6]), .Y(n5559) );
  AO21X1_LVT U6929 ( .A1(n3854), .A2(div_io_resp_bits_data[6]), .A3(n5559), 
        .Y(n5560) );
  AO22X1_LVT U6930 ( .A1(n3933), .A2(n_T_427[1413]), .A3(n_T_427[1285]), .A4(
        n3927), .Y(n5564) );
  AO22X1_LVT U6931 ( .A1(n3943), .A2(n_T_427[1157]), .A3(n_T_427[1221]), .A4(
        n3937), .Y(n5563) );
  AO22X1_LVT U6932 ( .A1(n3953), .A2(n_T_427[1093]), .A3(n_T_427[965]), .A4(
        n3947), .Y(n5562) );
  AO22X1_LVT U6933 ( .A1(n3900), .A2(n_T_427[1029]), .A3(n_T_427[70]), .A4(
        n3832), .Y(n5561) );
  NOR4X1_LVT U6934 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .Y(n5577)
         );
  AO22X1_LVT U6935 ( .A1(n3906), .A2(n_T_427[773]), .A3(n_T_427[710]), .A4(
        n2827), .Y(n5566) );
  AO22X1_LVT U6936 ( .A1(n1919), .A2(n_T_427[326]), .A3(n_T_427[6]), .A4(n3914), .Y(n5565) );
  AO22X1_LVT U6937 ( .A1(n6867), .A2(n_T_427[390]), .A3(n3859), .A4(
        n_T_427[198]), .Y(n5570) );
  AO22X1_LVT U6938 ( .A1(n3870), .A2(n_T_427[518]), .A3(n_T_427[454]), .A4(
        n3836), .Y(n5569) );
  AO22X1_LVT U6939 ( .A1(n_T_427[901]), .A2(n3811), .A3(n3871), .A4(
        n_T_427[262]), .Y(n5568) );
  AO22X1_LVT U6940 ( .A1(n3816), .A2(n_T_427[134]), .A3(n_T_427[837]), .A4(
        n3874), .Y(n5567) );
  NOR4X1_LVT U6941 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .Y(n5571)
         );
  AOI22X1_LVT U6942 ( .A1(n3915), .A2(n_T_427[582]), .A3(n_T_427[646]), .A4(
        n6812), .Y(n5573) );
  NAND2X0_LVT U6943 ( .A1(n4336), .A2(n3958), .Y(n5572) );
  AND3X1_LVT U6944 ( .A1(n5574), .A2(n5573), .A3(n5572), .Y(n5575) );
  NAND4X0_LVT U6945 ( .A1(n5577), .A2(n5578), .A3(n5576), .A4(n5575), .Y(
        id_rs_1[6]) );
  NAND2X0_LVT U6946 ( .A1(io_fpu_dmem_resp_data[6]), .A2(n9165), .Y(n5582) );
  NAND2X0_LVT U6947 ( .A1(n_T_918[6]), .A2(n6899), .Y(n5581) );
  NAND2X0_LVT U6948 ( .A1(io_imem_sfence_bits_addr[6]), .A2(n6900), .Y(n5580)
         );
  NAND2X0_LVT U6949 ( .A1(n_T_635[6]), .A2(n3243), .Y(n5579) );
  NAND4X0_LVT U6950 ( .A1(n5582), .A2(n5581), .A3(n5580), .A4(n5579), .Y(
        n_T_702[6]) );
  AO222X1_LVT U6951 ( .A1(mem_br_target[7]), .A2(n6249), .A3(n6856), .A4(
        io_fpu_toint_data[7]), .A5(n6855), .A6(n_T_918[7]), .Y(N605) );
  AO22X1_LVT U6952 ( .A1(n6860), .A2(io_dmem_resp_bits_data[7]), .A3(n3847), 
        .A4(io_imem_sfence_bits_addr[7]), .Y(n5583) );
  AO21X1_LVT U6953 ( .A1(n3854), .A2(div_io_resp_bits_data[7]), .A3(n5583), 
        .Y(n5584) );
  AO22X1_LVT U6954 ( .A1(n3829), .A2(n_T_427[1797]), .A3(n_T_427[1670]), .A4(
        n3825), .Y(n5588) );
  AO22X1_LVT U6955 ( .A1(n3891), .A2(n_T_427[1542]), .A3(n_T_427[1606]), .A4(
        n3885), .Y(n5587) );
  AO22X1_LVT U6956 ( .A1(n3923), .A2(n_T_427[1478]), .A3(n_T_427[1350]), .A4(
        n3917), .Y(n5586) );
  AO22X1_LVT U6957 ( .A1(n3933), .A2(n_T_427[1414]), .A3(n_T_427[1286]), .A4(
        n3927), .Y(n5585) );
  NOR4X1_LVT U6958 ( .A1(n5588), .A2(n5587), .A3(n5586), .A4(n5585), .Y(n5602)
         );
  AO22X1_LVT U6959 ( .A1(n2860), .A2(n_T_427[774]), .A3(n_T_427[391]), .A4(
        n2865), .Y(n5590) );
  AO22X1_LVT U6960 ( .A1(n1918), .A2(n_T_427[327]), .A3(n_T_427[583]), .A4(
        n2870), .Y(n5589) );
  NOR2X0_LVT U6961 ( .A1(n5590), .A2(n5589), .Y(n5600) );
  AO22X1_LVT U6962 ( .A1(n_T_427[647]), .A2(n3863), .A3(n3804), .A4(
        n_T_427[711]), .Y(n5594) );
  AO22X1_LVT U6963 ( .A1(n3870), .A2(n_T_427[519]), .A3(n_T_427[455]), .A4(
        n3836), .Y(n5593) );
  AO22X1_LVT U6964 ( .A1(n_T_427[838]), .A2(n6871), .A3(n3871), .A4(
        n_T_427[263]), .Y(n5592) );
  AO22X1_LVT U6965 ( .A1(n3816), .A2(n_T_427[135]), .A3(n6838), .A4(n_T_427[7]), .Y(n5591) );
  NOR4X1_LVT U6966 ( .A1(n5594), .A2(n5593), .A3(n5592), .A4(n5591), .Y(n5595)
         );
  AOI22X1_LVT U6967 ( .A1(n3801), .A2(n_T_427[1853]), .A3(n_T_427[1734]), .A4(
        n2866), .Y(n5597) );
  NAND2X0_LVT U6968 ( .A1(n4339), .A2(n3958), .Y(n5596) );
  AND3X1_LVT U6969 ( .A1(n5598), .A2(n5597), .A3(n5596), .Y(n5599) );
  NAND4X0_LVT U6970 ( .A1(n5602), .A2(n5601), .A3(n5600), .A4(n5599), .Y(
        id_rs_1[7]) );
  AO22X1_LVT U6971 ( .A1(n6860), .A2(io_dmem_resp_bits_data[8]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[8]), .Y(n5603) );
  AO21X1_LVT U6972 ( .A1(n3854), .A2(div_io_resp_bits_data[8]), .A3(n5603), 
        .Y(n5604) );
  AO22X1_LVT U6973 ( .A1(n3933), .A2(n_T_427[1415]), .A3(n_T_427[1287]), .A4(
        n3927), .Y(n5608) );
  AO22X1_LVT U6974 ( .A1(n3943), .A2(n_T_427[1159]), .A3(n_T_427[1223]), .A4(
        n3937), .Y(n5607) );
  AO22X1_LVT U6975 ( .A1(n3953), .A2(n_T_427[1095]), .A3(n_T_427[967]), .A4(
        n3947), .Y(n5606) );
  AO22X1_LVT U6976 ( .A1(n3900), .A2(n_T_427[1031]), .A3(n_T_427[903]), .A4(
        n2831), .Y(n5605) );
  NOR4X1_LVT U6977 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .Y(n5621)
         );
  AO22X1_LVT U6978 ( .A1(n3907), .A2(n_T_427[775]), .A3(n_T_427[72]), .A4(
        n2871), .Y(n5610) );
  AO22X1_LVT U6979 ( .A1(n3911), .A2(n_T_427[456]), .A3(n_T_427[8]), .A4(n3913), .Y(n5609) );
  NOR2X0_LVT U6980 ( .A1(n5610), .A2(n5609), .Y(n5620) );
  AO22X1_LVT U6981 ( .A1(n6765), .A2(n_T_427[712]), .A3(n3865), .A4(
        n_T_427[392]), .Y(n5614) );
  AO22X1_LVT U6982 ( .A1(n_T_427[648]), .A2(n3863), .A3(n3859), .A4(
        n_T_427[200]), .Y(n5613) );
  AO22X1_LVT U6983 ( .A1(n3870), .A2(n_T_427[520]), .A3(n_T_427[584]), .A4(
        n3795), .Y(n5612) );
  AO22X1_LVT U6984 ( .A1(n6796), .A2(n_T_427[136]), .A3(n_T_427[839]), .A4(
        n3875), .Y(n5611) );
  NOR4X1_LVT U6985 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .Y(n5615)
         );
  AOI22X1_LVT U6986 ( .A1(n3817), .A2(n_T_427[328]), .A3(n_T_427[264]), .A4(
        n3810), .Y(n5617) );
  NAND2X0_LVT U6987 ( .A1(n4342), .A2(n3959), .Y(n5616) );
  AND3X1_LVT U6988 ( .A1(n5618), .A2(n5617), .A3(n5616), .Y(n5619) );
  NAND4X0_LVT U6989 ( .A1(n5621), .A2(n5622), .A3(n5620), .A4(n5619), .Y(
        id_rs_1[8]) );
  NAND2X0_LVT U6990 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[8]), .Y(n5626) );
  NAND2X0_LVT U6991 ( .A1(n6899), .A2(n_T_918[8]), .Y(n5625) );
  NAND2X0_LVT U6992 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[8]), .Y(n5624)
         );
  NAND2X0_LVT U6993 ( .A1(n6901), .A2(n_T_635[8]), .Y(n5623) );
  NAND4X0_LVT U6994 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .Y(
        n_T_702[8]) );
  AO22X1_LVT U6995 ( .A1(n6860), .A2(io_dmem_resp_bits_data[9]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[9]), .Y(n5627) );
  AO21X1_LVT U6996 ( .A1(n3854), .A2(div_io_resp_bits_data[9]), .A3(n5627), 
        .Y(n5628) );
  AO22X1_LVT U6997 ( .A1(n3934), .A2(n_T_427[1416]), .A3(n_T_427[1288]), .A4(
        n3927), .Y(n5632) );
  AO22X1_LVT U6998 ( .A1(n3944), .A2(n_T_427[1160]), .A3(n_T_427[1224]), .A4(
        n3937), .Y(n5631) );
  AO22X1_LVT U6999 ( .A1(n3954), .A2(n_T_427[1096]), .A3(n_T_427[968]), .A4(
        n3947), .Y(n5630) );
  AO22X1_LVT U7000 ( .A1(n3899), .A2(n_T_427[1032]), .A3(n_T_427[201]), .A4(
        n3806), .Y(n5629) );
  NOR4X1_LVT U7001 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .Y(n5645)
         );
  AO22X1_LVT U7002 ( .A1(n3834), .A2(n_T_427[393]), .A3(n_T_427[73]), .A4(
        n3833), .Y(n5634) );
  AO22X1_LVT U7003 ( .A1(n3817), .A2(n_T_427[329]), .A3(n_T_427[713]), .A4(
        n3903), .Y(n5633) );
  NOR2X0_LVT U7004 ( .A1(n5634), .A2(n5633), .Y(n5644) );
  AO22X1_LVT U7005 ( .A1(n3797), .A2(n_T_427[585]), .A3(n_T_427[457]), .A4(
        n3836), .Y(n5638) );
  AO22X1_LVT U7006 ( .A1(n_T_427[904]), .A2(n3811), .A3(n3871), .A4(
        n_T_427[265]), .Y(n5637) );
  AO22X1_LVT U7007 ( .A1(n3814), .A2(n_T_427[776]), .A3(n_T_427[840]), .A4(
        n3874), .Y(n5636) );
  AO22X1_LVT U7008 ( .A1(n3816), .A2(n_T_427[137]), .A3(n6838), .A4(n_T_427[9]), .Y(n5635) );
  NOR4X1_LVT U7009 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .Y(n5639)
         );
  AOI22X1_LVT U7010 ( .A1(n2851), .A2(n_T_427[521]), .A3(n_T_427[649]), .A4(
        n3821), .Y(n5641) );
  NAND2X0_LVT U7011 ( .A1(n4345), .A2(n3958), .Y(n5640) );
  AND3X1_LVT U7012 ( .A1(n5642), .A2(n5641), .A3(n5640), .Y(n5643) );
  NAND4X0_LVT U7013 ( .A1(n5645), .A2(n5646), .A3(n5644), .A4(n5643), .Y(
        id_rs_1[9]) );
  NAND2X0_LVT U7014 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[9]), .Y(n5650) );
  NAND2X0_LVT U7015 ( .A1(n6899), .A2(n_T_918[9]), .Y(n5649) );
  NAND2X0_LVT U7016 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[9]), .Y(n5648)
         );
  NAND2X0_LVT U7017 ( .A1(n3243), .A2(n_T_635[9]), .Y(n5647) );
  NAND4X0_LVT U7018 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .Y(
        n_T_702[9]) );
  AO22X1_LVT U7019 ( .A1(n3851), .A2(io_dmem_resp_bits_data[10]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[10]), .Y(n5651) );
  AO21X1_LVT U7020 ( .A1(n3854), .A2(div_io_resp_bits_data[10]), .A3(n5651), 
        .Y(n5652) );
  AO22X1_LVT U7021 ( .A1(n3933), .A2(n_T_427[1417]), .A3(n_T_427[1289]), .A4(
        n3927), .Y(n5656) );
  AO22X1_LVT U7022 ( .A1(n3943), .A2(n_T_427[1161]), .A3(n_T_427[1225]), .A4(
        n3937), .Y(n5655) );
  AO22X1_LVT U7023 ( .A1(n3953), .A2(n_T_427[1097]), .A3(n_T_427[969]), .A4(
        n3947), .Y(n5654) );
  AO22X1_LVT U7024 ( .A1(n3900), .A2(n_T_427[1033]), .A3(n3806), .A4(
        n_T_427[202]), .Y(n5653) );
  NOR4X1_LVT U7025 ( .A1(n5656), .A2(n5655), .A3(n5654), .A4(n5653), .Y(n5669)
         );
  AO22X1_LVT U7026 ( .A1(n2864), .A2(n_T_427[394]), .A3(n_T_427[458]), .A4(
        n3912), .Y(n5658) );
  AO22X1_LVT U7027 ( .A1(n3833), .A2(n_T_427[74]), .A3(n_T_427[905]), .A4(
        n3897), .Y(n5657) );
  AO22X1_LVT U7028 ( .A1(n_T_427[650]), .A2(n3863), .A3(n3804), .A4(
        n_T_427[714]), .Y(n5662) );
  AO22X1_LVT U7029 ( .A1(n3814), .A2(n_T_427[777]), .A3(n_T_427[841]), .A4(
        n3874), .Y(n5661) );
  AO22X1_LVT U7030 ( .A1(n_T_427[522]), .A2(n3868), .A3(n3872), .A4(
        n_T_427[266]), .Y(n5660) );
  AO22X1_LVT U7031 ( .A1(n6796), .A2(n_T_427[138]), .A3(n3839), .A4(
        n_T_427[10]), .Y(n5659) );
  NOR4X1_LVT U7032 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .Y(n5663)
         );
  AOI22X1_LVT U7033 ( .A1(n2857), .A2(n_T_427[330]), .A3(n_T_427[586]), .A4(
        n2869), .Y(n5665) );
  NAND2X0_LVT U7034 ( .A1(n4348), .A2(n3958), .Y(n5664) );
  AND3X1_LVT U7035 ( .A1(n5666), .A2(n5665), .A3(n5664), .Y(n5667) );
  NAND4X0_LVT U7036 ( .A1(n5669), .A2(n5670), .A3(n5668), .A4(n5667), .Y(
        id_rs_1[10]) );
  NAND2X0_LVT U7037 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[10]), .Y(n5674) );
  NAND2X0_LVT U7038 ( .A1(n6899), .A2(n_T_918[10]), .Y(n5673) );
  NAND2X0_LVT U7039 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[10]), .Y(n5672)
         );
  NAND2X0_LVT U7040 ( .A1(n3243), .A2(n_T_635[10]), .Y(n5671) );
  NAND4X0_LVT U7041 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .Y(
        n_T_702[10]) );
  AO22X1_LVT U7042 ( .A1(n2861), .A2(n_T_427[778]), .A3(n_T_427[587]), .A4(
        n3915), .Y(n5676) );
  AO22X1_LVT U7043 ( .A1(n3896), .A2(n_T_427[906]), .A3(n_T_427[139]), .A4(
        n3908), .Y(n5675) );
  AO22X1_LVT U7044 ( .A1(n6867), .A2(n_T_427[395]), .A3(n3859), .A4(
        n_T_427[203]), .Y(n5680) );
  AO22X1_LVT U7045 ( .A1(n_T_427[715]), .A2(n3804), .A3(n3864), .A4(
        n_T_427[75]), .Y(n5679) );
  AO22X1_LVT U7046 ( .A1(n_T_427[651]), .A2(n3863), .A3(n3867), .A4(
        n_T_427[331]), .Y(n5678) );
  AO22X1_LVT U7047 ( .A1(n3837), .A2(n_T_427[459]), .A3(n3872), .A4(
        n_T_427[267]), .Y(n5677) );
  NOR4X1_LVT U7048 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .Y(n5681)
         );
  AO22X1_LVT U7049 ( .A1(n3851), .A2(io_dmem_resp_bits_data[12]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[12]), .Y(n5682) );
  AO21X1_LVT U7050 ( .A1(n3854), .A2(div_io_resp_bits_data[12]), .A3(n5682), 
        .Y(n5683) );
  AO22X1_LVT U7051 ( .A1(n3933), .A2(n_T_427[1419]), .A3(n_T_427[1291]), .A4(
        n3927), .Y(n5687) );
  AO22X1_LVT U7052 ( .A1(n3943), .A2(n_T_427[1163]), .A3(n_T_427[1227]), .A4(
        n3937), .Y(n5686) );
  AO22X1_LVT U7053 ( .A1(n3953), .A2(n_T_427[1099]), .A3(n_T_427[971]), .A4(
        n3947), .Y(n5685) );
  AO22X1_LVT U7054 ( .A1(n3900), .A2(n_T_427[1035]), .A3(n_T_427[76]), .A4(
        n2871), .Y(n5684) );
  NOR4X1_LVT U7055 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .Y(n5700)
         );
  AO22X1_LVT U7056 ( .A1(n2856), .A2(n_T_427[332]), .A3(n_T_427[588]), .A4(
        n3916), .Y(n5689) );
  AO22X1_LVT U7057 ( .A1(n3907), .A2(n_T_427[779]), .A3(n_T_427[716]), .A4(
        n3903), .Y(n5688) );
  AO22X1_LVT U7058 ( .A1(n6867), .A2(n_T_427[396]), .A3(n3859), .A4(
        n_T_427[204]), .Y(n5693) );
  AO22X1_LVT U7059 ( .A1(n3870), .A2(n_T_427[524]), .A3(n_T_427[460]), .A4(
        n3836), .Y(n5692) );
  AO22X1_LVT U7060 ( .A1(n_T_427[907]), .A2(n3811), .A3(n3872), .A4(
        n_T_427[268]), .Y(n5691) );
  AO22X1_LVT U7061 ( .A1(n3816), .A2(n_T_427[140]), .A3(n6838), .A4(
        n_T_427[12]), .Y(n5690) );
  NOR4X1_LVT U7062 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .Y(n5694)
         );
  AOI22X1_LVT U7063 ( .A1(n2833), .A2(n_T_427[843]), .A3(n_T_427[652]), .A4(
        n2829), .Y(n5696) );
  NAND2X0_LVT U7064 ( .A1(n4354), .A2(n3958), .Y(n5695) );
  AND3X1_LVT U7065 ( .A1(n5697), .A2(n5696), .A3(n5695), .Y(n5698) );
  NAND4X0_LVT U7066 ( .A1(n5700), .A2(n5701), .A3(n5699), .A4(n5698), .Y(
        id_rs_1[12]) );
  NAND2X0_LVT U7067 ( .A1(io_fpu_dmem_resp_data[12]), .A2(n9165), .Y(n5705) );
  NAND2X0_LVT U7068 ( .A1(n_T_918[12]), .A2(n6899), .Y(n5704) );
  NAND2X0_LVT U7069 ( .A1(io_imem_sfence_bits_addr[12]), .A2(n6900), .Y(n5703)
         );
  NAND2X0_LVT U7070 ( .A1(n_T_635[12]), .A2(n6901), .Y(n5702) );
  NAND4X0_LVT U7071 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .Y(
        n_T_702[12]) );
  AO22X1_LVT U7072 ( .A1(n3851), .A2(io_dmem_resp_bits_data[13]), .A3(n3850), 
        .A4(io_imem_sfence_bits_addr[13]), .Y(n5706) );
  AO21X1_LVT U7073 ( .A1(n3855), .A2(div_io_resp_bits_data[13]), .A3(n5706), 
        .Y(n5707) );
  AO22X1_LVT U7074 ( .A1(n3832), .A2(n_T_427[77]), .A3(n_T_427[717]), .A4(
        n3905), .Y(n5718) );
  AO22X1_LVT U7075 ( .A1(n2826), .A2(n_T_427[13]), .A3(n_T_427[141]), .A4(
        n3908), .Y(n5717) );
  AO22X1_LVT U7076 ( .A1(n2857), .A2(n_T_427[333]), .A3(n_T_427[525]), .A4(
        n3818), .Y(n5716) );
  AO22X1_LVT U7077 ( .A1(n_T_427[653]), .A2(n3863), .A3(n3796), .A4(
        n_T_427[589]), .Y(n5711) );
  AO22X1_LVT U7078 ( .A1(n6867), .A2(n_T_427[397]), .A3(n3859), .A4(
        n_T_427[205]), .Y(n5710) );
  AO22X1_LVT U7079 ( .A1(n_T_427[461]), .A2(n3837), .A3(n3872), .A4(
        n_T_427[269]), .Y(n5709) );
  AO22X1_LVT U7080 ( .A1(n3814), .A2(n_T_427[780]), .A3(n_T_427[844]), .A4(
        n3875), .Y(n5708) );
  NOR4X1_LVT U7081 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .Y(n5712)
         );
  NAND2X0_LVT U7082 ( .A1(n4356), .A2(n3958), .Y(n5713) );
  NAND2X0_LVT U7083 ( .A1(n5714), .A2(n5713), .Y(n5715) );
  NOR4X1_LVT U7084 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), .Y(n5725)
         );
  AO22X1_LVT U7085 ( .A1(n3933), .A2(n_T_427[1420]), .A3(n_T_427[1292]), .A4(
        n3927), .Y(n5722) );
  AO22X1_LVT U7086 ( .A1(n3943), .A2(n_T_427[1164]), .A3(n_T_427[1228]), .A4(
        n3938), .Y(n5721) );
  AO22X1_LVT U7087 ( .A1(n3953), .A2(n_T_427[1100]), .A3(n_T_427[972]), .A4(
        n3948), .Y(n5720) );
  AO22X1_LVT U7088 ( .A1(n3899), .A2(n_T_427[1036]), .A3(n_T_427[908]), .A4(
        n3897), .Y(n5719) );
  NOR4X1_LVT U7089 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .Y(n5723)
         );
  NAND3X0_LVT U7090 ( .A1(n5725), .A2(n5724), .A3(n5723), .Y(id_rs_1[13]) );
  NAND2X0_LVT U7091 ( .A1(io_fpu_dmem_resp_data[13]), .A2(n9165), .Y(n5729) );
  NAND2X0_LVT U7092 ( .A1(n_T_918[13]), .A2(n6899), .Y(n5728) );
  NAND2X0_LVT U7093 ( .A1(io_imem_sfence_bits_addr[13]), .A2(n6900), .Y(n5727)
         );
  NAND2X0_LVT U7094 ( .A1(n_T_635[13]), .A2(n6901), .Y(n5726) );
  NAND4X0_LVT U7095 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .Y(
        n_T_702[13]) );
  AO22X1_LVT U7096 ( .A1(n3851), .A2(io_dmem_resp_bits_data[14]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[14]), .Y(n5730) );
  AO21X1_LVT U7097 ( .A1(n3855), .A2(div_io_resp_bits_data[14]), .A3(n5730), 
        .Y(n5731) );
  AO22X1_LVT U7098 ( .A1(n_T_427[909]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[462]), .Y(n5735) );
  AO22X1_LVT U7099 ( .A1(n_T_427[654]), .A2(n3863), .A3(n3859), .A4(
        n_T_427[206]), .Y(n5734) );
  AO22X1_LVT U7100 ( .A1(n_T_427[718]), .A2(n3804), .A3(n3864), .A4(
        n_T_427[78]), .Y(n5733) );
  AO22X1_LVT U7101 ( .A1(n3816), .A2(n_T_427[142]), .A3(n3872), .A4(
        n_T_427[270]), .Y(n5732) );
  OR4X1_LVT U7102 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .Y(n5736)
         );
  AO22X1_LVT U7103 ( .A1(n3835), .A2(n_T_427[398]), .A3(n_T_427[1037]), .A4(
        n3898), .Y(n5740) );
  AO22X1_LVT U7104 ( .A1(n3906), .A2(n_T_427[781]), .A3(n_T_427[14]), .A4(
        n2826), .Y(n5739) );
  AO22X1_LVT U7105 ( .A1(n2856), .A2(n_T_427[334]), .A3(n_T_427[590]), .A4(
        n2870), .Y(n5738) );
  AO22X1_LVT U7106 ( .A1(n2850), .A2(n_T_427[526]), .A3(n_T_427[845]), .A4(
        n6813), .Y(n5737) );
  NAND2X0_LVT U7107 ( .A1(io_fpu_dmem_resp_data[14]), .A2(n9165), .Y(n5744) );
  NAND2X0_LVT U7108 ( .A1(n_T_918[14]), .A2(n6899), .Y(n5743) );
  NAND2X0_LVT U7109 ( .A1(io_imem_sfence_bits_addr[14]), .A2(n6900), .Y(n5742)
         );
  NAND2X0_LVT U7110 ( .A1(n_T_635[14]), .A2(n6901), .Y(n5741) );
  NAND4X0_LVT U7111 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .Y(
        n_T_702[14]) );
  AO22X1_LVT U7112 ( .A1(n3851), .A2(io_dmem_resp_bits_data[15]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[15]), .Y(n5745) );
  AO21X1_LVT U7113 ( .A1(n3855), .A2(div_io_resp_bits_data[15]), .A3(n5745), 
        .Y(n5746) );
  AO22X1_LVT U7114 ( .A1(n3835), .A2(n_T_427[399]), .A3(n_T_427[79]), .A4(
        n3833), .Y(n5757) );
  AO22X1_LVT U7115 ( .A1(n2860), .A2(n_T_427[782]), .A3(n_T_427[463]), .A4(
        n3911), .Y(n5756) );
  AO22X1_LVT U7116 ( .A1(n1919), .A2(n_T_427[335]), .A3(n_T_427[591]), .A4(
        n3916), .Y(n5755) );
  AO22X1_LVT U7117 ( .A1(n_T_427[655]), .A2(n3863), .A3(n3804), .A4(
        n_T_427[719]), .Y(n5750) );
  AO22X1_LVT U7118 ( .A1(n_T_427[910]), .A2(n3811), .A3(n3868), .A4(
        n_T_427[527]), .Y(n5749) );
  AO22X1_LVT U7119 ( .A1(n_T_427[846]), .A2(n3874), .A3(n3872), .A4(
        n_T_427[271]), .Y(n5748) );
  AO22X1_LVT U7120 ( .A1(n3816), .A2(n_T_427[143]), .A3(n3840), .A4(
        n_T_427[15]), .Y(n5747) );
  NOR4X1_LVT U7121 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .Y(n5751)
         );
  NAND2X0_LVT U7122 ( .A1(n4361), .A2(n3958), .Y(n5752) );
  NAND2X0_LVT U7123 ( .A1(n5753), .A2(n5752), .Y(n5754) );
  NOR4X1_LVT U7124 ( .A1(n5757), .A2(n5756), .A3(n5755), .A4(n5754), .Y(n5764)
         );
  AO22X1_LVT U7125 ( .A1(n3934), .A2(n_T_427[1422]), .A3(n_T_427[1294]), .A4(
        n3928), .Y(n5761) );
  AO22X1_LVT U7126 ( .A1(n3944), .A2(n_T_427[1166]), .A3(n_T_427[1230]), .A4(
        n3938), .Y(n5760) );
  AO22X1_LVT U7127 ( .A1(n3954), .A2(n_T_427[1102]), .A3(n_T_427[974]), .A4(
        n3948), .Y(n5759) );
  AO22X1_LVT U7128 ( .A1(n3899), .A2(n_T_427[1038]), .A3(n_T_427[207]), .A4(
        n3806), .Y(n5758) );
  NOR4X1_LVT U7129 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .Y(n5762)
         );
  NAND3X0_LVT U7130 ( .A1(n5764), .A2(n5763), .A3(n5762), .Y(id_rs_1[15]) );
  NAND2X0_LVT U7131 ( .A1(io_fpu_dmem_resp_data[15]), .A2(n9165), .Y(n5768) );
  NAND2X0_LVT U7132 ( .A1(n_T_918[15]), .A2(n6899), .Y(n5767) );
  NAND2X0_LVT U7133 ( .A1(io_imem_sfence_bits_addr[15]), .A2(n6900), .Y(n5766)
         );
  NAND2X0_LVT U7134 ( .A1(n_T_635[15]), .A2(n6901), .Y(n5765) );
  NAND4X0_LVT U7135 ( .A1(n5768), .A2(n5767), .A3(n5766), .A4(n5765), .Y(
        n_T_702[15]) );
  NAND2X0_LVT U7136 ( .A1(csr_io_rw_rdata[16]), .A2(n3844), .Y(n5771) );
  AOI22X1_LVT U7137 ( .A1(n3852), .A2(io_dmem_resp_bits_data[16]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[16]), .Y(n5770) );
  NAND2X0_LVT U7138 ( .A1(div_io_resp_bits_data[16]), .A2(n3856), .Y(n5769) );
  NAND3X0_LVT U7139 ( .A1(n5771), .A2(n5770), .A3(n5769), .Y(
        n_T_427__T_1136_data[16]) );
  AOI22X1_LVT U7140 ( .A1(n3870), .A2(n_T_427[528]), .A3(n3867), .A4(
        n_T_427[336]), .Y(n5775) );
  AOI22X1_LVT U7141 ( .A1(n3874), .A2(n_T_427[847]), .A3(n3840), .A4(
        n_T_427[16]), .Y(n5774) );
  OA22X1_LVT U7142 ( .A1(n3521), .A2(n6423), .A3(n3175), .A4(n6422), .Y(n5773)
         );
  AOI22X1_LVT U7143 ( .A1(n_T_427[911]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[592]), .Y(n5772) );
  NAND4X0_LVT U7144 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .Y(n5776) );
  NAND2X0_LVT U7145 ( .A1(csr_io_rw_rdata[17]), .A2(n3844), .Y(n5779) );
  AOI22X1_LVT U7146 ( .A1(n3852), .A2(io_dmem_resp_bits_data[17]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[17]), .Y(n5778) );
  NAND2X0_LVT U7147 ( .A1(div_io_resp_bits_data[17]), .A2(n3858), .Y(n5777) );
  NAND3X0_LVT U7148 ( .A1(n5779), .A2(n5778), .A3(n5777), .Y(
        n_T_427__T_1136_data[17]) );
  AO22X1_LVT U7149 ( .A1(n3816), .A2(n_T_427[145]), .A3(n_T_427[784]), .A4(
        n3812), .Y(n5783) );
  AO22X1_LVT U7150 ( .A1(n3797), .A2(n_T_427[593]), .A3(n_T_427[465]), .A4(
        n3836), .Y(n5782) );
  AO22X1_LVT U7151 ( .A1(n_T_427[912]), .A2(n3811), .A3(n3872), .A4(
        n_T_427[273]), .Y(n5781) );
  AO22X1_LVT U7152 ( .A1(n3859), .A2(n_T_427[209]), .A3(n3864), .A4(
        n_T_427[81]), .Y(n5780) );
  NOR4X1_LVT U7153 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .Y(n5784)
         );
  OA22X1_LVT U7154 ( .A1(n3541), .A2(n3799), .A3(n3139), .A4(n3803), .Y(n5787)
         );
  OA22X1_LVT U7155 ( .A1(n3142), .A2(n3081), .A3(n3494), .A4(n3082), .Y(n5786)
         );
  AOI22X1_LVT U7156 ( .A1(n3894), .A2(n_T_427[1552]), .A3(n_T_427[1616]), .A4(
        n3889), .Y(n5785) );
  AND4X1_LVT U7157 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .Y(n5796)
         );
  AO22X1_LVT U7158 ( .A1(n3924), .A2(n_T_427[1488]), .A3(n_T_427[1360]), .A4(
        n3918), .Y(n5792) );
  AO22X1_LVT U7159 ( .A1(n3934), .A2(n_T_427[1424]), .A3(n_T_427[1296]), .A4(
        n3928), .Y(n5791) );
  AO22X1_LVT U7160 ( .A1(n3944), .A2(n_T_427[1168]), .A3(n_T_427[1232]), .A4(
        n3938), .Y(n5790) );
  AO22X1_LVT U7161 ( .A1(n3954), .A2(n_T_427[1104]), .A3(n_T_427[976]), .A4(
        n3948), .Y(n5789) );
  NOR4X1_LVT U7162 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .Y(n5795)
         );
  NAND2X0_LVT U7163 ( .A1(n3958), .A2(n4367), .Y(n5793) );
  NAND4X0_LVT U7164 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .Y(
        id_rs_1[17]) );
  NAND2X0_LVT U7165 ( .A1(io_fpu_dmem_resp_data[17]), .A2(n9165), .Y(n5800) );
  NAND2X0_LVT U7166 ( .A1(n_T_918[17]), .A2(n6899), .Y(n5799) );
  NAND2X0_LVT U7167 ( .A1(io_imem_sfence_bits_addr[17]), .A2(n6900), .Y(n5798)
         );
  NAND2X0_LVT U7168 ( .A1(n_T_635[17]), .A2(n3243), .Y(n5797) );
  NAND4X0_LVT U7169 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .Y(
        n_T_702[17]) );
  AO22X1_LVT U7170 ( .A1(n3852), .A2(io_dmem_resp_bits_data[18]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[18]), .Y(n5801) );
  AO21X1_LVT U7171 ( .A1(n3855), .A2(div_io_resp_bits_data[18]), .A3(n5801), 
        .Y(n5802) );
  AO21X1_LVT U7172 ( .A1(n3843), .A2(csr_io_rw_rdata[18]), .A3(n5802), .Y(
        n_T_427__T_1136_data[18]) );
  AO22X1_LVT U7173 ( .A1(n3934), .A2(n_T_427[1425]), .A3(n_T_427[1297]), .A4(
        n3928), .Y(n5806) );
  AO22X1_LVT U7174 ( .A1(n3944), .A2(n_T_427[1169]), .A3(n_T_427[1233]), .A4(
        n3938), .Y(n5805) );
  AO22X1_LVT U7175 ( .A1(n3954), .A2(n_T_427[1105]), .A3(n_T_427[977]), .A4(
        n3948), .Y(n5804) );
  AO22X1_LVT U7176 ( .A1(n3900), .A2(n_T_427[1041]), .A3(n_T_427[913]), .A4(
        n2832), .Y(n5803) );
  NOR4X1_LVT U7177 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .Y(n5819)
         );
  AO22X1_LVT U7178 ( .A1(n2824), .A2(n_T_427[466]), .A3(n_T_427[722]), .A4(
        n3904), .Y(n5808) );
  AO22X1_LVT U7179 ( .A1(n2826), .A2(n_T_427[18]), .A3(n_T_427[146]), .A4(
        n3909), .Y(n5807) );
  NOR2X0_LVT U7180 ( .A1(n5808), .A2(n5807), .Y(n5818) );
  AOI22X1_LVT U7181 ( .A1(n2833), .A2(n_T_427[849]), .A3(n_T_427[274]), .A4(
        n2828), .Y(n5816) );
  NAND2X0_LVT U7182 ( .A1(n4370), .A2(n3959), .Y(n5815) );
  AO22X1_LVT U7183 ( .A1(n_T_427[658]), .A2(n3862), .A3(n3859), .A4(
        n_T_427[210]), .Y(n5812) );
  AO22X1_LVT U7184 ( .A1(n3813), .A2(n_T_427[785]), .A3(n_T_427[594]), .A4(
        n3795), .Y(n5811) );
  AO22X1_LVT U7185 ( .A1(n6867), .A2(n_T_427[402]), .A3(n3864), .A4(
        n_T_427[82]), .Y(n5810) );
  AO22X1_LVT U7186 ( .A1(n_T_427[530]), .A2(n3868), .A3(n6868), .A4(
        n_T_427[338]), .Y(n5809) );
  NOR4X1_LVT U7187 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .Y(n5813)
         );
  AND3X1_LVT U7188 ( .A1(n5816), .A2(n5815), .A3(n5814), .Y(n5817) );
  NAND4X0_LVT U7189 ( .A1(n5819), .A2(n5820), .A3(n5818), .A4(n5817), .Y(
        id_rs_1[18]) );
  NAND2X0_LVT U7190 ( .A1(io_fpu_dmem_resp_data[18]), .A2(n9165), .Y(n5824) );
  NAND2X0_LVT U7191 ( .A1(n_T_918[18]), .A2(n6899), .Y(n5823) );
  NAND2X0_LVT U7192 ( .A1(io_imem_sfence_bits_addr[18]), .A2(n6900), .Y(n5822)
         );
  NAND2X0_LVT U7193 ( .A1(n_T_635[18]), .A2(n3243), .Y(n5821) );
  NAND4X0_LVT U7194 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .Y(
        n_T_702[18]) );
  AO22X1_LVT U7195 ( .A1(n3852), .A2(io_dmem_resp_bits_data[19]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[19]), .Y(n5825) );
  AO21X1_LVT U7196 ( .A1(n3855), .A2(div_io_resp_bits_data[19]), .A3(n5825), 
        .Y(n5826) );
  AO21X1_LVT U7197 ( .A1(n3843), .A2(csr_io_rw_rdata[19]), .A3(n5826), .Y(
        n_T_427__T_1136_data[19]) );
  AO22X1_LVT U7198 ( .A1(n_T_427[659]), .A2(n3862), .A3(n3804), .A4(
        n_T_427[723]), .Y(n5830) );
  AO22X1_LVT U7199 ( .A1(n_T_427[914]), .A2(n3811), .A3(n3875), .A4(
        n_T_427[850]), .Y(n5829) );
  AO22X1_LVT U7200 ( .A1(n3869), .A2(n_T_427[531]), .A3(n_T_427[595]), .A4(
        n3795), .Y(n5828) );
  AO22X1_LVT U7201 ( .A1(n3815), .A2(n_T_427[147]), .A3(n3840), .A4(
        n_T_427[19]), .Y(n5827) );
  NOR4X1_LVT U7202 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .Y(n5831)
         );
  OA22X1_LVT U7203 ( .A1(n3543), .A2(n3881), .A3(n3878), .A4(n5831), .Y(n5833)
         );
  NAND2X0_LVT U7204 ( .A1(n4373), .A2(n3959), .Y(n5832) );
  NAND2X0_LVT U7205 ( .A1(io_fpu_dmem_resp_data[19]), .A2(n9165), .Y(n5837) );
  NAND2X0_LVT U7206 ( .A1(n_T_918[19]), .A2(n6899), .Y(n5836) );
  NAND2X0_LVT U7207 ( .A1(io_imem_sfence_bits_addr[19]), .A2(n6900), .Y(n5835)
         );
  NAND2X0_LVT U7208 ( .A1(n_T_635[19]), .A2(n3243), .Y(n5834) );
  NAND4X0_LVT U7209 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .Y(
        n_T_702[19]) );
  AO22X1_LVT U7210 ( .A1(n3852), .A2(io_dmem_resp_bits_data[20]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[20]), .Y(n5838) );
  AO21X1_LVT U7211 ( .A1(n3855), .A2(div_io_resp_bits_data[20]), .A3(n5838), 
        .Y(n5839) );
  AO21X1_LVT U7212 ( .A1(n3844), .A2(csr_io_rw_rdata[20]), .A3(n5839), .Y(
        n_T_427__T_1136_data[20]) );
  AO22X1_LVT U7213 ( .A1(n3933), .A2(n_T_427[1427]), .A3(n_T_427[1299]), .A4(
        n3928), .Y(n5843) );
  AO22X1_LVT U7214 ( .A1(n3943), .A2(n_T_427[1171]), .A3(n_T_427[1235]), .A4(
        n3938), .Y(n5842) );
  AO22X1_LVT U7215 ( .A1(n3953), .A2(n_T_427[1107]), .A3(n_T_427[979]), .A4(
        n3948), .Y(n5841) );
  AO22X1_LVT U7216 ( .A1(n3900), .A2(n_T_427[1043]), .A3(n_T_427[915]), .A4(
        n3896), .Y(n5840) );
  NOR4X1_LVT U7217 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .Y(n5856)
         );
  AO22X1_LVT U7218 ( .A1(n3835), .A2(n_T_427[404]), .A3(n_T_427[724]), .A4(
        n2827), .Y(n5845) );
  AO22X1_LVT U7219 ( .A1(n3913), .A2(n_T_427[20]), .A3(n_T_427[148]), .A4(
        n2863), .Y(n5844) );
  AO22X1_LVT U7220 ( .A1(n3869), .A2(n_T_427[532]), .A3(n_T_427[596]), .A4(
        n3795), .Y(n5849) );
  AO22X1_LVT U7221 ( .A1(n_T_427[660]), .A2(n3862), .A3(n3866), .A4(
        n_T_427[340]), .Y(n5848) );
  AO22X1_LVT U7222 ( .A1(n3813), .A2(n_T_427[787]), .A3(n_T_427[468]), .A4(
        n3836), .Y(n5847) );
  AO22X1_LVT U7223 ( .A1(n3860), .A2(n_T_427[212]), .A3(n6866), .A4(
        n_T_427[84]), .Y(n5846) );
  NOR4X1_LVT U7224 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .Y(n5850)
         );
  OA22X1_LVT U7225 ( .A1(n3544), .A2(n3881), .A3(n3878), .A4(n5850), .Y(n5853)
         );
  AOI22X1_LVT U7226 ( .A1(n3823), .A2(n_T_427[851]), .A3(n_T_427[276]), .A4(
        n3809), .Y(n5852) );
  NAND2X0_LVT U7227 ( .A1(n4376), .A2(n3959), .Y(n5851) );
  AND3X1_LVT U7228 ( .A1(n5853), .A2(n5852), .A3(n5851), .Y(n5854) );
  NAND4X0_LVT U7229 ( .A1(n5856), .A2(n5857), .A3(n5855), .A4(n5854), .Y(
        id_rs_1[20]) );
  NAND2X0_LVT U7230 ( .A1(io_fpu_dmem_resp_data[20]), .A2(n9165), .Y(n5861) );
  NAND2X0_LVT U7231 ( .A1(n_T_918[20]), .A2(n6899), .Y(n5860) );
  NAND2X0_LVT U7232 ( .A1(io_imem_sfence_bits_addr[20]), .A2(n6900), .Y(n5859)
         );
  NAND2X0_LVT U7233 ( .A1(n_T_635[20]), .A2(n6901), .Y(n5858) );
  NAND4X0_LVT U7234 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .Y(
        n_T_702[20]) );
  AO22X1_LVT U7235 ( .A1(n3852), .A2(io_dmem_resp_bits_data[21]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[21]), .Y(n5862) );
  AO21X1_LVT U7236 ( .A1(n3855), .A2(div_io_resp_bits_data[21]), .A3(n5862), 
        .Y(n5863) );
  AO22X1_LVT U7237 ( .A1(n_T_427[916]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[597]), .Y(n5867) );
  AO22X1_LVT U7238 ( .A1(n_T_427[661]), .A2(n3862), .A3(n3859), .A4(
        n_T_427[213]), .Y(n5866) );
  AO22X1_LVT U7239 ( .A1(n_T_427[725]), .A2(n6765), .A3(n3864), .A4(
        n_T_427[85]), .Y(n5865) );
  AO22X1_LVT U7240 ( .A1(n_T_427[852]), .A2(n3875), .A3(n3839), .A4(
        n_T_427[21]), .Y(n5864) );
  NOR4X1_LVT U7241 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .Y(n5868)
         );
  OA22X1_LVT U7242 ( .A1(n3095), .A2(n3596), .A3(n3878), .A4(n5868), .Y(n5870)
         );
  NAND2X0_LVT U7243 ( .A1(n_T_427[533]), .A2(n3819), .Y(n5869) );
  AO22X1_LVT U7244 ( .A1(n3921), .A2(n_T_427[1364]), .A3(n_T_427[1428]), .A4(
        n3932), .Y(n5874) );
  AO22X1_LVT U7245 ( .A1(n3928), .A2(n_T_427[1300]), .A3(n_T_427[1172]), .A4(
        n3942), .Y(n5873) );
  AO22X1_LVT U7246 ( .A1(n3941), .A2(n_T_427[1236]), .A3(n_T_427[1108]), .A4(
        n3952), .Y(n5872) );
  AO22X1_LVT U7247 ( .A1(n3951), .A2(n_T_427[980]), .A3(n_T_427[1044]), .A4(
        n3898), .Y(n5871) );
  NOR4X1_LVT U7248 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .Y(n5875)
         );
  NAND3X0_LVT U7249 ( .A1(n5877), .A2(n5876), .A3(n5875), .Y(id_rs_1[21]) );
  NAND2X0_LVT U7250 ( .A1(io_fpu_dmem_resp_data[21]), .A2(n9165), .Y(n5881) );
  NAND2X0_LVT U7251 ( .A1(n_T_918[21]), .A2(n6899), .Y(n5880) );
  NAND2X0_LVT U7252 ( .A1(io_imem_sfence_bits_addr[21]), .A2(n6900), .Y(n5879)
         );
  NAND2X0_LVT U7253 ( .A1(n_T_635[21]), .A2(n6901), .Y(n5878) );
  NAND4X0_LVT U7254 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .Y(
        n_T_702[21]) );
  AO22X1_LVT U7255 ( .A1(n3921), .A2(n_T_427[1365]), .A3(n_T_427[1429]), .A4(
        n3932), .Y(n5885) );
  AO22X1_LVT U7256 ( .A1(n3931), .A2(n_T_427[1301]), .A3(n_T_427[1173]), .A4(
        n3942), .Y(n5884) );
  AO22X1_LVT U7257 ( .A1(n3941), .A2(n_T_427[1237]), .A3(n_T_427[1109]), .A4(
        n3952), .Y(n5883) );
  AO22X1_LVT U7258 ( .A1(n3951), .A2(n_T_427[981]), .A3(n_T_427[1045]), .A4(
        n3899), .Y(n5882) );
  NOR4X1_LVT U7259 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .Y(n5896)
         );
  AO22X1_LVT U7260 ( .A1(n6765), .A2(n_T_427[726]), .A3(n3865), .A4(
        n_T_427[406]), .Y(n5889) );
  AO22X1_LVT U7261 ( .A1(n_T_427[662]), .A2(n3862), .A3(n3860), .A4(
        n_T_427[214]), .Y(n5888) );
  AO22X1_LVT U7262 ( .A1(n_T_427[853]), .A2(n6871), .A3(n3872), .A4(
        n_T_427[278]), .Y(n5887) );
  AO22X1_LVT U7263 ( .A1(n3815), .A2(n_T_427[150]), .A3(n_T_427[789]), .A4(
        n3812), .Y(n5886) );
  NOR4X1_LVT U7264 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .Y(n5890)
         );
  OA22X1_LVT U7265 ( .A1(n3094), .A2(n3596), .A3(n3878), .A4(n5890), .Y(n5893)
         );
  AOI22X1_LVT U7266 ( .A1(n2850), .A2(n_T_427[534]), .A3(n_T_427[22]), .A4(
        n3913), .Y(n5892) );
  NAND2X0_LVT U7267 ( .A1(n_T_427[598]), .A2(n2870), .Y(n5891) );
  AND3X1_LVT U7268 ( .A1(n5893), .A2(n5892), .A3(n5891), .Y(n5894) );
  NAND4X0_LVT U7269 ( .A1(n5897), .A2(n5895), .A3(n5896), .A4(n5894), .Y(
        id_rs_1[22]) );
  NAND2X0_LVT U7270 ( .A1(io_fpu_dmem_resp_data[22]), .A2(n9165), .Y(n5901) );
  NAND2X0_LVT U7271 ( .A1(n_T_918[22]), .A2(n6899), .Y(n5900) );
  NAND2X0_LVT U7272 ( .A1(io_imem_sfence_bits_addr[22]), .A2(n6900), .Y(n5899)
         );
  NAND2X0_LVT U7273 ( .A1(n_T_635[22]), .A2(n3243), .Y(n5898) );
  NAND4X0_LVT U7274 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .Y(
        n_T_702[22]) );
  NAND2X0_LVT U7275 ( .A1(csr_io_rw_rdata[23]), .A2(n3844), .Y(n5904) );
  AOI22X1_LVT U7276 ( .A1(n3852), .A2(io_dmem_resp_bits_data[23]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[23]), .Y(n5903) );
  NAND2X0_LVT U7277 ( .A1(div_io_resp_bits_data[23]), .A2(n3858), .Y(n5902) );
  NAND3X0_LVT U7278 ( .A1(n5904), .A2(n5903), .A3(n5902), .Y(
        n_T_427__T_1136_data[23]) );
  AOI22X1_LVT U7279 ( .A1(n3870), .A2(n_T_427[535]), .A3(n_T_427[599]), .A4(
        n3795), .Y(n5910) );
  AOI22X1_LVT U7280 ( .A1(n3814), .A2(n_T_427[790]), .A3(n3871), .A4(
        n_T_427[279]), .Y(n5909) );
  AOI22X1_LVT U7281 ( .A1(n6765), .A2(n_T_427[727]), .A3(n6868), .A4(
        n_T_427[343]), .Y(n5908) );
  OA22X1_LVT U7282 ( .A1(n5906), .A2(n3526), .A3(n3177), .A4(n5905), .Y(n5907)
         );
  NAND4X0_LVT U7283 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .Y(n5911) );
  AO22X1_LVT U7284 ( .A1(n3924), .A2(n_T_427[1494]), .A3(n_T_427[1366]), .A4(
        n3918), .Y(n5915) );
  AO22X1_LVT U7285 ( .A1(n3934), .A2(n_T_427[1430]), .A3(n_T_427[1302]), .A4(
        n3928), .Y(n5914) );
  AO22X1_LVT U7286 ( .A1(n3944), .A2(n_T_427[1174]), .A3(n_T_427[1238]), .A4(
        n3938), .Y(n5913) );
  AO22X1_LVT U7287 ( .A1(n3954), .A2(n_T_427[1110]), .A3(n_T_427[982]), .A4(
        n3948), .Y(n5912) );
  NOR4X1_LVT U7288 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .Y(n5922)
         );
  AO22X1_LVT U7289 ( .A1(n2865), .A2(n_T_427[407]), .A3(n_T_427[471]), .A4(
        n3911), .Y(n5919) );
  AO22X1_LVT U7290 ( .A1(n3900), .A2(n_T_427[1046]), .A3(n_T_427[215]), .A4(
        n3808), .Y(n5918) );
  AO22X1_LVT U7291 ( .A1(n2871), .A2(n_T_427[87]), .A3(n_T_427[918]), .A4(
        n3897), .Y(n5917) );
  AO22X1_LVT U7292 ( .A1(n2833), .A2(n_T_427[854]), .A3(n_T_427[663]), .A4(
        n3820), .Y(n5916) );
  NOR4X1_LVT U7293 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .Y(n5921)
         );
  NAND2X0_LVT U7294 ( .A1(n3957), .A2(n4383), .Y(n5920) );
  NAND4X0_LVT U7295 ( .A1(n5922), .A2(n5923), .A3(n5921), .A4(n5920), .Y(
        id_rs_1[23]) );
  NAND2X0_LVT U7296 ( .A1(io_fpu_dmem_resp_data[23]), .A2(n9165), .Y(n5927) );
  NAND2X0_LVT U7297 ( .A1(n_T_918[23]), .A2(n6899), .Y(n5926) );
  NAND2X0_LVT U7298 ( .A1(io_imem_sfence_bits_addr[23]), .A2(n6900), .Y(n5925)
         );
  NAND2X0_LVT U7299 ( .A1(n_T_635[23]), .A2(n3243), .Y(n5924) );
  NAND4X0_LVT U7300 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .Y(
        n_T_702[23]) );
  AO22X1_LVT U7301 ( .A1(n3852), .A2(io_dmem_resp_bits_data[24]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[24]), .Y(n5928) );
  AO21X1_LVT U7302 ( .A1(n3855), .A2(div_io_resp_bits_data[24]), .A3(n5928), 
        .Y(n5929) );
  AO21X1_LVT U7303 ( .A1(n3844), .A2(csr_io_rw_rdata[24]), .A3(n5929), .Y(
        n_T_427__T_1136_data[24]) );
  AO22X1_LVT U7304 ( .A1(n3944), .A2(n_T_427[1175]), .A3(n_T_427[1239]), .A4(
        n3938), .Y(n5933) );
  AO22X1_LVT U7305 ( .A1(n3954), .A2(n_T_427[1111]), .A3(n_T_427[983]), .A4(
        n3948), .Y(n5932) );
  AO22X1_LVT U7306 ( .A1(n3900), .A2(n_T_427[1047]), .A3(n_T_427[216]), .A4(
        n2830), .Y(n5931) );
  AO22X1_LVT U7307 ( .A1(n3907), .A2(n_T_427[791]), .A3(n_T_427[408]), .A4(
        n3834), .Y(n5930) );
  NOR4X1_LVT U7308 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .Y(n5946)
         );
  AO22X1_LVT U7309 ( .A1(n3817), .A2(n_T_427[344]), .A3(n_T_427[600]), .A4(
        n2869), .Y(n5935) );
  AO22X1_LVT U7310 ( .A1(n3912), .A2(n_T_427[472]), .A3(n_T_427[24]), .A4(
        n2879), .Y(n5934) );
  NAND2X0_LVT U7311 ( .A1(n4386), .A2(n3959), .Y(n5943) );
  AO22X1_LVT U7312 ( .A1(n_T_427[664]), .A2(n3862), .A3(n3868), .A4(
        n_T_427[536]), .Y(n5939) );
  AO22X1_LVT U7313 ( .A1(n3815), .A2(n_T_427[152]), .A3(n_T_427[855]), .A4(
        n3874), .Y(n5938) );
  AO22X1_LVT U7314 ( .A1(n_T_427[728]), .A2(n6765), .A3(n3864), .A4(
        n_T_427[88]), .Y(n5937) );
  AO22X1_LVT U7315 ( .A1(n_T_427[919]), .A2(n3811), .A3(n3872), .A4(
        n_T_427[280]), .Y(n5936) );
  NOR4X1_LVT U7316 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .Y(n5940)
         );
  OA22X1_LVT U7317 ( .A1(n3545), .A2(n3881), .A3(n3878), .A4(n5940), .Y(n5942)
         );
  OA22X1_LVT U7318 ( .A1(n3546), .A2(n3799), .A3(n3137), .A4(n3803), .Y(n5941)
         );
  AND3X1_LVT U7319 ( .A1(n5943), .A2(n5942), .A3(n5941), .Y(n5944) );
  NAND4X0_LVT U7320 ( .A1(n5946), .A2(n5947), .A3(n5945), .A4(n5944), .Y(
        id_rs_1[24]) );
  NAND2X0_LVT U7321 ( .A1(io_fpu_dmem_resp_data[24]), .A2(n9165), .Y(n5951) );
  NAND2X0_LVT U7322 ( .A1(n_T_918[24]), .A2(n6899), .Y(n5950) );
  NAND2X0_LVT U7323 ( .A1(io_imem_sfence_bits_addr[24]), .A2(n6900), .Y(n5949)
         );
  NAND2X0_LVT U7324 ( .A1(n_T_635[24]), .A2(n6901), .Y(n5948) );
  NAND4X0_LVT U7325 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .Y(
        n_T_702[24]) );
  AO22X1_LVT U7326 ( .A1(n3852), .A2(io_dmem_resp_bits_data[25]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[25]), .Y(n5952) );
  AO21X1_LVT U7327 ( .A1(n3855), .A2(div_io_resp_bits_data[25]), .A3(n5952), 
        .Y(n5953) );
  AO22X1_LVT U7328 ( .A1(n3907), .A2(n_T_427[792]), .A3(n_T_427[217]), .A4(
        n3807), .Y(n5964) );
  AO22X1_LVT U7329 ( .A1(n2872), .A2(n_T_427[89]), .A3(n_T_427[153]), .A4(
        n3909), .Y(n5963) );
  AO22X1_LVT U7330 ( .A1(n2824), .A2(n_T_427[473]), .A3(n_T_427[537]), .A4(
        n2851), .Y(n5962) );
  AO22X1_LVT U7331 ( .A1(n_T_427[920]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[601]), .Y(n5957) );
  AO22X1_LVT U7332 ( .A1(n3804), .A2(n_T_427[729]), .A3(n3865), .A4(
        n_T_427[409]), .Y(n5956) );
  AO22X1_LVT U7333 ( .A1(n_T_427[665]), .A2(n3862), .A3(n3867), .A4(
        n_T_427[345]), .Y(n5955) );
  AO22X1_LVT U7334 ( .A1(n_T_427[856]), .A2(n3875), .A3(n3872), .A4(
        n_T_427[281]), .Y(n5954) );
  NOR4X1_LVT U7335 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .Y(n5958)
         );
  OA22X1_LVT U7336 ( .A1(n3097), .A2(n3596), .A3(n3878), .A4(n5958), .Y(n5960)
         );
  NAND2X0_LVT U7337 ( .A1(n_T_427[25]), .A2(n3914), .Y(n5959) );
  NAND2X0_LVT U7338 ( .A1(n5960), .A2(n5959), .Y(n5961) );
  AO22X1_LVT U7339 ( .A1(n2866), .A2(n_T_427[1752]), .A3(n_T_427[1814]), .A4(
        n3829), .Y(n5967) );
  AO22X1_LVT U7340 ( .A1(n_T_427[1868]), .A2(n3802), .A3(n3884), .A4(
        n_T_427[1906]), .Y(n5966) );
  AO22X1_LVT U7341 ( .A1(n3826), .A2(n_T_427[1688]), .A3(n_T_427[1560]), .A4(
        n3890), .Y(n5965) );
  NAND2X0_LVT U7342 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[25]), .Y(n5971) );
  NAND2X0_LVT U7343 ( .A1(n_T_918[25]), .A2(n6899), .Y(n5970) );
  NAND2X0_LVT U7344 ( .A1(io_imem_sfence_bits_addr[25]), .A2(n6900), .Y(n5969)
         );
  NAND2X0_LVT U7345 ( .A1(n_T_635[25]), .A2(n6901), .Y(n5968) );
  NAND4X0_LVT U7346 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .Y(
        n_T_702[25]) );
  AO22X1_LVT U7347 ( .A1(n3852), .A2(io_dmem_resp_bits_data[26]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[26]), .Y(n5972) );
  AO21X1_LVT U7348 ( .A1(n3855), .A2(div_io_resp_bits_data[26]), .A3(n5972), 
        .Y(n5973) );
  AO22X1_LVT U7349 ( .A1(n3921), .A2(n_T_427[1369]), .A3(n_T_427[1433]), .A4(
        n3932), .Y(n5977) );
  AO22X1_LVT U7350 ( .A1(n3931), .A2(n_T_427[1305]), .A3(n_T_427[1177]), .A4(
        n3942), .Y(n5976) );
  AO22X1_LVT U7351 ( .A1(n3941), .A2(n_T_427[1241]), .A3(n_T_427[1113]), .A4(
        n3952), .Y(n5975) );
  AO22X1_LVT U7352 ( .A1(n3951), .A2(n_T_427[985]), .A3(n_T_427[1049]), .A4(
        n3898), .Y(n5974) );
  NOR4X1_LVT U7353 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .Y(n5990)
         );
  AO22X1_LVT U7354 ( .A1(n3831), .A2(n_T_427[90]), .A3(n_T_427[218]), .A4(
        n2830), .Y(n5979) );
  AO22X1_LVT U7355 ( .A1(n2857), .A2(n_T_427[346]), .A3(n_T_427[921]), .A4(
        n3895), .Y(n5978) );
  AO22X1_LVT U7356 ( .A1(n6765), .A2(n_T_427[730]), .A3(n_T_427[602]), .A4(
        n3795), .Y(n5983) );
  AO22X1_LVT U7357 ( .A1(n3813), .A2(n_T_427[793]), .A3(n_T_427[857]), .A4(
        n3874), .Y(n5982) );
  AO22X1_LVT U7358 ( .A1(n3837), .A2(n_T_427[474]), .A3(n3872), .A4(
        n_T_427[282]), .Y(n5981) );
  AO22X1_LVT U7359 ( .A1(n3815), .A2(n_T_427[154]), .A3(n6838), .A4(
        n_T_427[26]), .Y(n5980) );
  NOR4X1_LVT U7360 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .Y(n5984)
         );
  OA22X1_LVT U7361 ( .A1(n3096), .A2(n3596), .A3(n3878), .A4(n5984), .Y(n5987)
         );
  AOI22X1_LVT U7362 ( .A1(n3835), .A2(n_T_427[410]), .A3(n_T_427[666]), .A4(
        n3820), .Y(n5986) );
  NAND2X0_LVT U7363 ( .A1(n_T_427[538]), .A2(n3818), .Y(n5985) );
  AND3X1_LVT U7364 ( .A1(n5987), .A2(n5986), .A3(n5985), .Y(n5988) );
  NAND4X0_LVT U7365 ( .A1(n5990), .A2(n5991), .A3(n5989), .A4(n5988), .Y(
        id_rs_1[26]) );
  NAND2X0_LVT U7366 ( .A1(io_fpu_dmem_resp_data[26]), .A2(n9165), .Y(n5995) );
  NAND2X0_LVT U7367 ( .A1(n_T_918[26]), .A2(n6899), .Y(n5994) );
  NAND2X0_LVT U7368 ( .A1(io_imem_sfence_bits_addr[26]), .A2(n6900), .Y(n5993)
         );
  NAND2X0_LVT U7369 ( .A1(n_T_635[26]), .A2(n3243), .Y(n5992) );
  NAND4X0_LVT U7370 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .Y(
        n_T_702[26]) );
  AO22X1_LVT U7371 ( .A1(n3852), .A2(io_dmem_resp_bits_data[27]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[27]), .Y(n5996) );
  AO21X1_LVT U7372 ( .A1(n3856), .A2(div_io_resp_bits_data[27]), .A3(n5996), 
        .Y(n5997) );
  AO21X1_LVT U7373 ( .A1(n3843), .A2(csr_io_rw_rdata[27]), .A3(n5997), .Y(
        n_T_427__T_1136_data[27]) );
  AOI22X1_LVT U7374 ( .A1(n3797), .A2(n_T_427[603]), .A3(n3871), .A4(
        n_T_427[283]), .Y(n6001) );
  AOI22X1_LVT U7375 ( .A1(n3814), .A2(n_T_427[794]), .A3(n_T_427[858]), .A4(
        n3875), .Y(n6000) );
  AOI22X1_LVT U7376 ( .A1(n6765), .A2(n_T_427[731]), .A3(n3864), .A4(
        n_T_427[91]), .Y(n5999) );
  AOI22X1_LVT U7377 ( .A1(n3863), .A2(n_T_427[667]), .A3(n3865), .A4(
        n_T_427[411]), .Y(n5998) );
  NAND4X0_LVT U7378 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .Y(n6002) );
  NAND2X0_LVT U7379 ( .A1(n6877), .A2(n6002), .Y(n6005) );
  NAND2X0_LVT U7380 ( .A1(n3957), .A2(n4393), .Y(n6004) );
  NAND2X0_LVT U7381 ( .A1(n_T_427[1908]), .A2(n3884), .Y(n6003) );
  AO22X1_LVT U7382 ( .A1(n3934), .A2(n_T_427[1434]), .A3(n_T_427[1306]), .A4(
        n3928), .Y(n6009) );
  AO22X1_LVT U7383 ( .A1(n3944), .A2(n_T_427[1178]), .A3(n_T_427[1242]), .A4(
        n3938), .Y(n6008) );
  AO22X1_LVT U7384 ( .A1(n3954), .A2(n_T_427[1114]), .A3(n_T_427[986]), .A4(
        n3948), .Y(n6007) );
  AO22X1_LVT U7385 ( .A1(n3900), .A2(n_T_427[1050]), .A3(n_T_427[219]), .A4(
        n2830), .Y(n6006) );
  NOR4X1_LVT U7386 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .Y(n6010)
         );
  NAND3X0_LVT U7387 ( .A1(n6012), .A2(n6011), .A3(n6010), .Y(id_rs_1[27]) );
  AO22X1_LVT U7388 ( .A1(n3851), .A2(io_dmem_resp_bits_data[28]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[28]), .Y(n6013) );
  AO21X1_LVT U7389 ( .A1(n3855), .A2(div_io_resp_bits_data[28]), .A3(n6013), 
        .Y(n6014) );
  AO22X1_LVT U7390 ( .A1(n2864), .A2(n_T_427[412]), .A3(n_T_427[220]), .A4(
        n3807), .Y(n6025) );
  AO22X1_LVT U7391 ( .A1(n2871), .A2(n_T_427[92]), .A3(n_T_427[28]), .A4(n3914), .Y(n6024) );
  AO22X1_LVT U7392 ( .A1(n3910), .A2(n_T_427[476]), .A3(n3810), .A4(
        n_T_427[284]), .Y(n6023) );
  AO22X1_LVT U7393 ( .A1(n_T_427[668]), .A2(n3862), .A3(n3804), .A4(
        n_T_427[732]), .Y(n6018) );
  AO22X1_LVT U7394 ( .A1(n_T_427[923]), .A2(n3811), .A3(n3875), .A4(
        n_T_427[859]), .Y(n6017) );
  AO22X1_LVT U7395 ( .A1(n3815), .A2(n_T_427[156]), .A3(n_T_427[795]), .A4(
        n3812), .Y(n6016) );
  AO22X1_LVT U7396 ( .A1(n_T_427[540]), .A2(n3869), .A3(n3866), .A4(
        n_T_427[348]), .Y(n6015) );
  NOR4X1_LVT U7397 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .Y(n6019)
         );
  OA22X1_LVT U7398 ( .A1(n3596), .A2(n3090), .A3(n3878), .A4(n6019), .Y(n6021)
         );
  NAND2X0_LVT U7399 ( .A1(n_T_427[604]), .A2(n3915), .Y(n6020) );
  NAND2X0_LVT U7400 ( .A1(n6021), .A2(n6020), .Y(n6022) );
  NAND2X0_LVT U7401 ( .A1(io_fpu_dmem_resp_data[28]), .A2(n9165), .Y(n6029) );
  NAND2X0_LVT U7402 ( .A1(n_T_918[28]), .A2(n6899), .Y(n6028) );
  NAND2X0_LVT U7403 ( .A1(io_imem_sfence_bits_addr[28]), .A2(n6900), .Y(n6027)
         );
  NAND2X0_LVT U7404 ( .A1(n_T_635[28]), .A2(n3243), .Y(n6026) );
  NAND4X0_LVT U7405 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .Y(
        n_T_702[28]) );
  AO22X1_LVT U7406 ( .A1(n3851), .A2(io_dmem_resp_bits_data[29]), .A3(n3849), 
        .A4(io_imem_sfence_bits_addr[29]), .Y(n6030) );
  AO21X1_LVT U7407 ( .A1(n3856), .A2(div_io_resp_bits_data[29]), .A3(n6030), 
        .Y(n6031) );
  AO21X1_LVT U7408 ( .A1(n3843), .A2(csr_io_rw_rdata[29]), .A3(n6031), .Y(
        n_T_427__T_1136_data[29]) );
  AO22X1_LVT U7409 ( .A1(n3831), .A2(n_T_427[93]), .A3(n_T_427[221]), .A4(
        n3808), .Y(n6041) );
  AO22X1_LVT U7410 ( .A1(n2832), .A2(n_T_427[924]), .A3(n_T_427[29]), .A4(
        n2879), .Y(n6040) );
  AO22X1_LVT U7411 ( .A1(n2865), .A2(n_T_427[413]), .A3(n_T_427[860]), .A4(
        n3823), .Y(n6039) );
  AOI22X1_LVT U7412 ( .A1(n3797), .A2(n_T_427[605]), .A3(n3867), .A4(
        n_T_427[349]), .Y(n6035) );
  AOI22X1_LVT U7413 ( .A1(n_T_427[477]), .A2(n3837), .A3(n3871), .A4(
        n_T_427[285]), .Y(n6034) );
  AOI22X1_LVT U7414 ( .A1(n3816), .A2(n_T_427[157]), .A3(n_T_427[796]), .A4(
        n3812), .Y(n6033) );
  AOI22X1_LVT U7415 ( .A1(n3863), .A2(n_T_427[669]), .A3(n3804), .A4(
        n_T_427[733]), .Y(n6032) );
  NAND4X0_LVT U7416 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .Y(n6036) );
  AO22X1_LVT U7417 ( .A1(n3957), .A2(n4398), .A3(n6036), .A4(n6877), .Y(n6037)
         );
  AO21X1_LVT U7418 ( .A1(n_T_427[541]), .A2(n3819), .A3(n6037), .Y(n6038) );
  NOR4X1_LVT U7419 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .Y(n6048)
         );
  AO22X1_LVT U7420 ( .A1(n3921), .A2(n_T_427[1372]), .A3(n_T_427[1436]), .A4(
        n3932), .Y(n6045) );
  AO22X1_LVT U7421 ( .A1(n3931), .A2(n_T_427[1308]), .A3(n_T_427[1180]), .A4(
        n3942), .Y(n6044) );
  AO22X1_LVT U7422 ( .A1(n3941), .A2(n_T_427[1244]), .A3(n_T_427[1116]), .A4(
        n3952), .Y(n6043) );
  AO22X1_LVT U7423 ( .A1(n3951), .A2(n_T_427[988]), .A3(n_T_427[1052]), .A4(
        n3899), .Y(n6042) );
  NOR4X1_LVT U7424 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .Y(n6046)
         );
  NAND3X0_LVT U7425 ( .A1(n6048), .A2(n6047), .A3(n6046), .Y(id_rs_1[29]) );
  NAND2X0_LVT U7426 ( .A1(io_fpu_dmem_resp_data[29]), .A2(n9165), .Y(n6052) );
  NAND2X0_LVT U7427 ( .A1(n_T_918[29]), .A2(n6899), .Y(n6051) );
  NAND2X0_LVT U7428 ( .A1(io_imem_sfence_bits_addr[29]), .A2(n6900), .Y(n6050)
         );
  NAND2X0_LVT U7429 ( .A1(n_T_635[29]), .A2(n3243), .Y(n6049) );
  NAND4X0_LVT U7430 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .Y(
        n_T_702[29]) );
  AO22X1_LVT U7431 ( .A1(n3851), .A2(io_dmem_resp_bits_data[30]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[30]), .Y(n6053) );
  AO21X1_LVT U7432 ( .A1(n3856), .A2(div_io_resp_bits_data[30]), .A3(n6053), 
        .Y(n6054) );
  AO21X1_LVT U7433 ( .A1(n3843), .A2(csr_io_rw_rdata[30]), .A3(n6054), .Y(
        n_T_427__T_1136_data[30]) );
  AO22X1_LVT U7434 ( .A1(n3830), .A2(n_T_427[1819]), .A3(n_T_427[1693]), .A4(
        n3827), .Y(n6058) );
  AO22X1_LVT U7435 ( .A1(n3892), .A2(n_T_427[1565]), .A3(n_T_427[1629]), .A4(
        n3886), .Y(n6057) );
  AO22X1_LVT U7436 ( .A1(n3924), .A2(n_T_427[1501]), .A3(n_T_427[1373]), .A4(
        n3918), .Y(n6056) );
  AO22X1_LVT U7437 ( .A1(n3934), .A2(n_T_427[1437]), .A3(n_T_427[1309]), .A4(
        n3928), .Y(n6055) );
  NOR4X1_LVT U7438 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .Y(n6076)
         );
  AO22X1_LVT U7439 ( .A1(n3944), .A2(n_T_427[1181]), .A3(n_T_427[1245]), .A4(
        n3938), .Y(n6062) );
  AO22X1_LVT U7440 ( .A1(n3954), .A2(n_T_427[1117]), .A3(n_T_427[989]), .A4(
        n3948), .Y(n6061) );
  AO22X1_LVT U7441 ( .A1(n3900), .A2(n_T_427[1053]), .A3(n_T_427[222]), .A4(
        n3806), .Y(n6060) );
  AO22X1_LVT U7442 ( .A1(n2865), .A2(n_T_427[414]), .A3(n_T_427[734]), .A4(
        n3904), .Y(n6059) );
  NOR4X1_LVT U7443 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .Y(n6075)
         );
  AO22X1_LVT U7444 ( .A1(n1918), .A2(n_T_427[350]), .A3(n_T_427[478]), .A4(
        n3910), .Y(n6064) );
  AO22X1_LVT U7445 ( .A1(n2851), .A2(n_T_427[542]), .A3(n_T_427[861]), .A4(
        n3822), .Y(n6063) );
  NOR2X0_LVT U7446 ( .A1(n6064), .A2(n6063), .Y(n6074) );
  AO22X1_LVT U7447 ( .A1(n_T_427[925]), .A2(n3811), .A3(n3796), .A4(
        n_T_427[606]), .Y(n6068) );
  AO22X1_LVT U7448 ( .A1(n_T_427[670]), .A2(n3862), .A3(n3864), .A4(
        n_T_427[94]), .Y(n6067) );
  AO22X1_LVT U7449 ( .A1(n_T_427[797]), .A2(n3812), .A3(n3872), .A4(
        n_T_427[286]), .Y(n6066) );
  AO22X1_LVT U7450 ( .A1(n3815), .A2(n_T_427[158]), .A3(n3840), .A4(
        n_T_427[30]), .Y(n6065) );
  NOR4X1_LVT U7451 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .Y(n6069)
         );
  OA22X1_LVT U7452 ( .A1(n3547), .A2(n3881), .A3(n3878), .A4(n6069), .Y(n6072)
         );
  OA22X1_LVT U7453 ( .A1(n3548), .A2(n3799), .A3(n3140), .A4(n3803), .Y(n6071)
         );
  NAND2X0_LVT U7454 ( .A1(n4401), .A2(n3959), .Y(n6070) );
  AND3X1_LVT U7455 ( .A1(n6072), .A2(n6071), .A3(n6070), .Y(n6073) );
  NAND4X0_LVT U7456 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .Y(
        id_rs_1[30]) );
  NAND2X0_LVT U7457 ( .A1(io_fpu_dmem_resp_data[30]), .A2(n9165), .Y(n6080) );
  NAND2X0_LVT U7458 ( .A1(n_T_918[30]), .A2(n6899), .Y(n6079) );
  NAND2X0_LVT U7459 ( .A1(io_imem_sfence_bits_addr[30]), .A2(n6900), .Y(n6078)
         );
  NAND2X0_LVT U7460 ( .A1(n_T_635[30]), .A2(n6901), .Y(n6077) );
  NAND4X0_LVT U7461 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .Y(
        n_T_702[30]) );
  AO22X1_LVT U7462 ( .A1(n6856), .A2(io_fpu_toint_data[31]), .A3(n6855), .A4(
        n_T_918[31]), .Y(n6081) );
  AO21X1_LVT U7463 ( .A1(mem_br_target[31]), .A2(n6249), .A3(n6081), .Y(N629)
         );
  AO22X1_LVT U7464 ( .A1(n3851), .A2(io_dmem_resp_bits_data[31]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[31]), .Y(n6082) );
  AO21X1_LVT U7465 ( .A1(n3856), .A2(div_io_resp_bits_data[31]), .A3(n6082), 
        .Y(n6083) );
  AO22X1_LVT U7466 ( .A1(n_T_427[671]), .A2(n3862), .A3(n3868), .A4(
        n_T_427[543]), .Y(n6087) );
  AO22X1_LVT U7467 ( .A1(n6867), .A2(n_T_427[415]), .A3(n3860), .A4(
        n_T_427[223]), .Y(n6086) );
  AO22X1_LVT U7468 ( .A1(n3837), .A2(n_T_427[479]), .A3(n3873), .A4(
        n_T_427[287]), .Y(n6085) );
  AO22X1_LVT U7469 ( .A1(n_T_427[798]), .A2(n3812), .A3(n3839), .A4(
        n_T_427[31]), .Y(n6084) );
  NOR4X1_LVT U7470 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .Y(n6088)
         );
  OA22X1_LVT U7471 ( .A1(n3099), .A2(n3596), .A3(n3878), .A4(n6088), .Y(n6090)
         );
  NAND2X0_LVT U7472 ( .A1(n_T_427[607]), .A2(n2869), .Y(n6089) );
  AO22X1_LVT U7473 ( .A1(n3921), .A2(n_T_427[1374]), .A3(n_T_427[1438]), .A4(
        n3932), .Y(n6094) );
  AO22X1_LVT U7474 ( .A1(n3931), .A2(n_T_427[1310]), .A3(n_T_427[1182]), .A4(
        n3942), .Y(n6093) );
  AO22X1_LVT U7475 ( .A1(n3941), .A2(n_T_427[1246]), .A3(n_T_427[1118]), .A4(
        n3952), .Y(n6092) );
  AO22X1_LVT U7476 ( .A1(n3951), .A2(n_T_427[990]), .A3(n_T_427[1054]), .A4(
        n3899), .Y(n6091) );
  NOR4X1_LVT U7477 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .Y(n6095)
         );
  NAND3X0_LVT U7478 ( .A1(n6097), .A2(n6096), .A3(n6095), .Y(id_rs_1[31]) );
  NAND2X0_LVT U7479 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[31]), .Y(n6101) );
  NAND2X0_LVT U7480 ( .A1(n_T_918[31]), .A2(n6899), .Y(n6100) );
  NAND2X0_LVT U7481 ( .A1(io_imem_sfence_bits_addr[31]), .A2(n6900), .Y(n6099)
         );
  NAND2X0_LVT U7482 ( .A1(n_T_635[31]), .A2(n6901), .Y(n6098) );
  NAND4X0_LVT U7483 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .Y(
        n_T_702[31]) );
  AO22X1_LVT U7484 ( .A1(n6856), .A2(io_fpu_toint_data[32]), .A3(n6855), .A4(
        n_T_918[32]), .Y(n6102) );
  AO21X1_LVT U7485 ( .A1(mem_br_target[32]), .A2(n6249), .A3(n6102), .Y(N630)
         );
  NAND2X0_LVT U7486 ( .A1(csr_io_rw_rdata[32]), .A2(n3844), .Y(n6105) );
  AOI22X1_LVT U7487 ( .A1(n3852), .A2(io_dmem_resp_bits_data[32]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[32]), .Y(n6104) );
  NAND2X0_LVT U7488 ( .A1(div_io_resp_bits_data[32]), .A2(n3858), .Y(n6103) );
  NAND3X0_LVT U7489 ( .A1(n6105), .A2(n6104), .A3(n6103), .Y(
        n_T_427__T_1136_data[32]) );
  AO22X1_LVT U7490 ( .A1(n_T_427[672]), .A2(n3862), .A3(n3865), .A4(
        n_T_427[416]), .Y(n6109) );
  AO22X1_LVT U7491 ( .A1(n3815), .A2(n_T_427[160]), .A3(n_T_427[799]), .A4(
        n3812), .Y(n6108) );
  AO22X1_LVT U7492 ( .A1(n3837), .A2(n_T_427[480]), .A3(n3866), .A4(
        n_T_427[352]), .Y(n6107) );
  AO22X1_LVT U7493 ( .A1(n_T_427[927]), .A2(n3811), .A3(n3873), .A4(
        n_T_427[288]), .Y(n6106) );
  NOR4X1_LVT U7494 ( .A1(n6109), .A2(n6108), .A3(n6107), .A4(n6106), .Y(n6110)
         );
  NAND2X0_LVT U7495 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[32]), .Y(n6114) );
  NAND2X0_LVT U7496 ( .A1(n6899), .A2(n_T_918[32]), .Y(n6113) );
  NAND2X0_LVT U7497 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[32]), .Y(n6112)
         );
  NAND2X0_LVT U7498 ( .A1(n3243), .A2(n_T_635[32]), .Y(n6111) );
  NAND4X0_LVT U7499 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .Y(
        n_T_702[32]) );
  AO22X1_LVT U7500 ( .A1(n6856), .A2(io_fpu_toint_data[33]), .A3(n6855), .A4(
        n_T_918[33]), .Y(n6115) );
  AO21X1_LVT U7501 ( .A1(mem_br_target[33]), .A2(n6249), .A3(n6115), .Y(N631)
         );
  NAND2X0_LVT U7502 ( .A1(csr_io_rw_rdata[33]), .A2(n3844), .Y(n6118) );
  AOI22X1_LVT U7503 ( .A1(n3853), .A2(io_dmem_resp_bits_data[33]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[33]), .Y(n6117) );
  NAND2X0_LVT U7504 ( .A1(div_io_resp_bits_data[33]), .A2(n3858), .Y(n6116) );
  AO22X1_LVT U7505 ( .A1(n3918), .A2(n_T_427[1376]), .A3(n_T_427[1440]), .A4(
        n3932), .Y(n6122) );
  AO22X1_LVT U7506 ( .A1(n3930), .A2(n_T_427[1312]), .A3(n_T_427[1184]), .A4(
        n3942), .Y(n6121) );
  AO22X1_LVT U7507 ( .A1(n3940), .A2(n_T_427[1248]), .A3(n_T_427[1120]), .A4(
        n3952), .Y(n6120) );
  AO22X1_LVT U7508 ( .A1(n3950), .A2(n_T_427[992]), .A3(n_T_427[1056]), .A4(
        n3899), .Y(n6119) );
  NOR4X1_LVT U7509 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .Y(n6133)
         );
  AO22X1_LVT U7510 ( .A1(n6765), .A2(n_T_427[737]), .A3(n3865), .A4(
        n_T_427[417]), .Y(n6126) );
  AO22X1_LVT U7511 ( .A1(n3869), .A2(n_T_427[545]), .A3(n_T_427[609]), .A4(
        n3795), .Y(n6125) );
  AO22X1_LVT U7512 ( .A1(n_T_427[673]), .A2(n3862), .A3(n3866), .A4(
        n_T_427[353]), .Y(n6124) );
  AO22X1_LVT U7513 ( .A1(n3813), .A2(n_T_427[800]), .A3(n_T_427[864]), .A4(
        n3874), .Y(n6123) );
  NOR4X1_LVT U7514 ( .A1(n6126), .A2(n6125), .A3(n6124), .A4(n6123), .Y(n6127)
         );
  OA22X1_LVT U7515 ( .A1(n3091), .A2(n3596), .A3(n3878), .A4(n6127), .Y(n6130)
         );
  AOI22X1_LVT U7516 ( .A1(n3911), .A2(n_T_427[481]), .A3(n_T_427[289]), .A4(
        n6774), .Y(n6129) );
  NAND2X0_LVT U7517 ( .A1(n_T_427[33]), .A2(n2879), .Y(n6128) );
  AND3X1_LVT U7518 ( .A1(n6130), .A2(n6129), .A3(n6128), .Y(n6131) );
  NAND4X0_LVT U7519 ( .A1(n6133), .A2(n6134), .A3(n6132), .A4(n6131), .Y(
        id_rs_1[33]) );
  NAND2X0_LVT U7520 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[33]), .Y(n6138) );
  NAND2X0_LVT U7521 ( .A1(n6899), .A2(n_T_918[33]), .Y(n6137) );
  NAND2X0_LVT U7522 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[33]), .Y(n6136)
         );
  NAND2X0_LVT U7523 ( .A1(n6901), .A2(n_T_635[33]), .Y(n6135) );
  NAND4X0_LVT U7524 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .Y(
        n_T_702[33]) );
  NAND2X0_LVT U7525 ( .A1(csr_io_rw_rdata[34]), .A2(n3844), .Y(n6141) );
  AOI22X1_LVT U7526 ( .A1(n3853), .A2(io_dmem_resp_bits_data[34]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[34]), .Y(n6140) );
  NAND2X0_LVT U7527 ( .A1(div_io_resp_bits_data[34]), .A2(n3858), .Y(n6139) );
  NAND3X0_LVT U7528 ( .A1(n6141), .A2(n6140), .A3(n6139), .Y(
        n_T_427__T_1136_data[34]) );
  AOI22X1_LVT U7529 ( .A1(n3816), .A2(n_T_427[162]), .A3(n_T_427[801]), .A4(
        n3812), .Y(n6145) );
  OA22X1_LVT U7530 ( .A1(n6767), .A2(n3527), .A3(n3141), .A4(n3805), .Y(n6144)
         );
  AOI22X1_LVT U7531 ( .A1(n_T_427[674]), .A2(n3861), .A3(n3868), .A4(
        n_T_427[546]), .Y(n6143) );
  AOI22X1_LVT U7532 ( .A1(n_T_427[929]), .A2(n6794), .A3(n3875), .A4(
        n_T_427[865]), .Y(n6142) );
  NAND4X0_LVT U7533 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .Y(n6146) );
  AO22X1_LVT U7534 ( .A1(n3924), .A2(n_T_427[1505]), .A3(n_T_427[1377]), .A4(
        n3919), .Y(n6150) );
  AO22X1_LVT U7535 ( .A1(n3934), .A2(n_T_427[1441]), .A3(n_T_427[1313]), .A4(
        n3929), .Y(n6149) );
  AO22X1_LVT U7536 ( .A1(n3944), .A2(n_T_427[1185]), .A3(n_T_427[1249]), .A4(
        n3939), .Y(n6148) );
  AO22X1_LVT U7537 ( .A1(n3954), .A2(n_T_427[1121]), .A3(n_T_427[993]), .A4(
        n3949), .Y(n6147) );
  NOR4X1_LVT U7538 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .Y(n6157)
         );
  AO22X1_LVT U7539 ( .A1(n2824), .A2(n_T_427[482]), .A3(n_T_427[98]), .A4(
        n2871), .Y(n6154) );
  AO22X1_LVT U7540 ( .A1(n3901), .A2(n_T_427[1057]), .A3(n_T_427[226]), .A4(
        n3807), .Y(n6153) );
  AO22X1_LVT U7541 ( .A1(n1919), .A2(n_T_427[354]), .A3(n_T_427[34]), .A4(
        n3913), .Y(n6152) );
  AO22X1_LVT U7542 ( .A1(n3916), .A2(n_T_427[610]), .A3(n_T_427[290]), .A4(
        n3810), .Y(n6151) );
  NOR4X1_LVT U7543 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .Y(n6156)
         );
  NAND2X0_LVT U7544 ( .A1(n3957), .A2(n4411), .Y(n6155) );
  NAND4X0_LVT U7545 ( .A1(n6157), .A2(n6158), .A3(n6156), .A4(n6155), .Y(
        id_rs_1[34]) );
  NAND2X0_LVT U7546 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[34]), .Y(n6162) );
  NAND2X0_LVT U7547 ( .A1(n6899), .A2(n_T_918[34]), .Y(n6161) );
  NAND2X0_LVT U7548 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[34]), .Y(n6160)
         );
  NAND2X0_LVT U7549 ( .A1(n3243), .A2(n_T_635[34]), .Y(n6159) );
  NAND4X0_LVT U7550 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .Y(
        n_T_702[34]) );
  AO22X1_LVT U7551 ( .A1(n6856), .A2(io_fpu_toint_data[35]), .A3(n6855), .A4(
        n_T_918[35]), .Y(n6163) );
  AO21X1_LVT U7552 ( .A1(mem_br_target[35]), .A2(n6249), .A3(n6163), .Y(N633)
         );
  NAND2X0_LVT U7553 ( .A1(csr_io_rw_rdata[35]), .A2(n3845), .Y(n6166) );
  AOI22X1_LVT U7554 ( .A1(n3853), .A2(io_dmem_resp_bits_data[35]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[35]), .Y(n6165) );
  NAND2X0_LVT U7555 ( .A1(div_io_resp_bits_data[35]), .A2(n3858), .Y(n6164) );
  AO22X1_LVT U7556 ( .A1(n3920), .A2(n_T_427[1378]), .A3(n_T_427[1442]), .A4(
        n3932), .Y(n6170) );
  AO22X1_LVT U7557 ( .A1(n3931), .A2(n_T_427[1314]), .A3(n_T_427[1186]), .A4(
        n3942), .Y(n6169) );
  AO22X1_LVT U7558 ( .A1(n3938), .A2(n_T_427[1250]), .A3(n_T_427[1122]), .A4(
        n3952), .Y(n6168) );
  AO22X1_LVT U7559 ( .A1(n3948), .A2(n_T_427[994]), .A3(n_T_427[1058]), .A4(
        n3899), .Y(n6167) );
  NOR4X1_LVT U7560 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .Y(n6183)
         );
  AO22X1_LVT U7561 ( .A1(n3835), .A2(n_T_427[419]), .A3(n_T_427[611]), .A4(
        n2870), .Y(n6172) );
  AO22X1_LVT U7562 ( .A1(n3806), .A2(n_T_427[227]), .A3(n_T_427[738]), .A4(
        n3903), .Y(n6171) );
  AOI22X1_LVT U7563 ( .A1(n6886), .A2(n_T_427[163]), .A3(n_T_427[675]), .A4(
        n2829), .Y(n6180) );
  NAND2X0_LVT U7564 ( .A1(n_T_427[291]), .A2(n3809), .Y(n6179) );
  AO22X1_LVT U7565 ( .A1(n_T_427[930]), .A2(n3811), .A3(n3875), .A4(
        n_T_427[866]), .Y(n6176) );
  AO22X1_LVT U7566 ( .A1(n3870), .A2(n_T_427[547]), .A3(n_T_427[483]), .A4(
        n3836), .Y(n6175) );
  AO22X1_LVT U7567 ( .A1(n_T_427[802]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[35]), .Y(n6174) );
  AO22X1_LVT U7568 ( .A1(n6866), .A2(n_T_427[99]), .A3(n3866), .A4(
        n_T_427[355]), .Y(n6173) );
  NOR4X1_LVT U7569 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .Y(n6177)
         );
  OA22X1_LVT U7570 ( .A1(n3183), .A2(n3596), .A3(n3878), .A4(n6177), .Y(n6178)
         );
  AND3X1_LVT U7571 ( .A1(n6180), .A2(n6179), .A3(n6178), .Y(n6181) );
  NAND4X0_LVT U7572 ( .A1(n6183), .A2(n6184), .A3(n6182), .A4(n6181), .Y(
        id_rs_1[35]) );
  NAND2X0_LVT U7573 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[35]), .Y(n6188) );
  NAND2X0_LVT U7574 ( .A1(n6899), .A2(n_T_918[35]), .Y(n6187) );
  NAND2X0_LVT U7575 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[35]), .Y(n6186)
         );
  NAND2X0_LVT U7576 ( .A1(n3243), .A2(n_T_635[35]), .Y(n6185) );
  NAND4X0_LVT U7577 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .Y(
        n_T_702[35]) );
  AO22X1_LVT U7578 ( .A1(n3851), .A2(io_dmem_resp_bits_data[36]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[36]), .Y(n6189) );
  AO21X1_LVT U7579 ( .A1(n3856), .A2(div_io_resp_bits_data[36]), .A3(n6189), 
        .Y(n6190) );
  AO21X1_LVT U7580 ( .A1(n3843), .A2(csr_io_rw_rdata[36]), .A3(n6190), .Y(
        n_T_427__T_1136_data[36]) );
  AO22X1_LVT U7581 ( .A1(n3916), .A2(n_T_427[612]), .A3(n_T_427[164]), .A4(
        n3909), .Y(n6192) );
  AO22X1_LVT U7582 ( .A1(n2828), .A2(n_T_427[292]), .A3(n_T_427[676]), .A4(
        n6812), .Y(n6191) );
  NOR2X0_LVT U7583 ( .A1(n6192), .A2(n6191), .Y(n6202) );
  AO22X1_LVT U7584 ( .A1(n3869), .A2(n_T_427[548]), .A3(n_T_427[867]), .A4(
        n3874), .Y(n6196) );
  AO22X1_LVT U7585 ( .A1(n6867), .A2(n_T_427[420]), .A3(n6866), .A4(
        n_T_427[100]), .Y(n6195) );
  AO22X1_LVT U7586 ( .A1(n3860), .A2(n_T_427[228]), .A3(n3866), .A4(
        n_T_427[356]), .Y(n6194) );
  AO22X1_LVT U7587 ( .A1(n_T_427[803]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[36]), .Y(n6193) );
  NOR4X1_LVT U7588 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .Y(n6197)
         );
  OA22X1_LVT U7589 ( .A1(n3549), .A2(n3881), .A3(n3878), .A4(n6197), .Y(n6200)
         );
  OA22X1_LVT U7590 ( .A1(n3145), .A2(n3803), .A3(n3497), .A4(n3800), .Y(n6199)
         );
  NAND2X0_LVT U7591 ( .A1(n4416), .A2(n3959), .Y(n6198) );
  AND3X1_LVT U7592 ( .A1(n6200), .A2(n6199), .A3(n6198), .Y(n6201) );
  NAND4X0_LVT U7593 ( .A1(n6203), .A2(n6204), .A3(n6202), .A4(n6201), .Y(
        id_rs_1[36]) );
  NAND2X0_LVT U7594 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[36]), .Y(n6208) );
  NAND2X0_LVT U7595 ( .A1(n6899), .A2(n_T_918[36]), .Y(n6207) );
  NAND2X0_LVT U7596 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[36]), .Y(n6206)
         );
  NAND2X0_LVT U7597 ( .A1(n3243), .A2(n_T_635[36]), .Y(n6205) );
  NAND4X0_LVT U7598 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .Y(
        n_T_702[36]) );
  NAND2X0_LVT U7599 ( .A1(csr_io_rw_rdata[37]), .A2(n3845), .Y(n6211) );
  AOI22X1_LVT U7600 ( .A1(n3853), .A2(io_dmem_resp_bits_data[37]), .A3(n3846), 
        .A4(io_imem_sfence_bits_addr[37]), .Y(n6210) );
  NAND2X0_LVT U7601 ( .A1(div_io_resp_bits_data[37]), .A2(n3858), .Y(n6209) );
  NAND3X0_LVT U7602 ( .A1(n6211), .A2(n6210), .A3(n6209), .Y(
        n_T_427__T_1136_data[37]) );
  AO22X1_LVT U7603 ( .A1(n3910), .A2(n_T_427[485]), .A3(n_T_427[165]), .A4(
        n2862), .Y(n6213) );
  AO22X1_LVT U7604 ( .A1(n3818), .A2(n_T_427[549]), .A3(n_T_427[868]), .A4(
        n3823), .Y(n6212) );
  NOR2X0_LVT U7605 ( .A1(n6213), .A2(n6212), .Y(n6223) );
  AO22X1_LVT U7606 ( .A1(n_T_427[677]), .A2(n3861), .A3(n3865), .A4(
        n_T_427[421]), .Y(n6217) );
  AO22X1_LVT U7607 ( .A1(n_T_427[613]), .A2(n3797), .A3(n3866), .A4(
        n_T_427[357]), .Y(n6216) );
  AO22X1_LVT U7608 ( .A1(n_T_427[932]), .A2(n3811), .A3(n3873), .A4(
        n_T_427[293]), .Y(n6215) );
  AO22X1_LVT U7609 ( .A1(n_T_427[804]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[37]), .Y(n6214) );
  NOR4X1_LVT U7610 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .Y(n6218)
         );
  OA22X1_LVT U7611 ( .A1(n3550), .A2(n3881), .A3(n3878), .A4(n6218), .Y(n6221)
         );
  OA22X1_LVT U7612 ( .A1(n3146), .A2(n3803), .A3(n3498), .A4(n3800), .Y(n6220)
         );
  NAND2X0_LVT U7613 ( .A1(n3957), .A2(n4419), .Y(n6219) );
  AND3X1_LVT U7614 ( .A1(n6221), .A2(n6220), .A3(n6219), .Y(n6222) );
  NAND4X0_LVT U7615 ( .A1(n6224), .A2(n6225), .A3(n6223), .A4(n6222), .Y(
        id_rs_1[37]) );
  NAND2X0_LVT U7616 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[37]), .Y(n6229) );
  NAND2X0_LVT U7617 ( .A1(n6899), .A2(n_T_918[37]), .Y(n6228) );
  NAND2X0_LVT U7618 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[37]), .Y(n6227)
         );
  NAND2X0_LVT U7619 ( .A1(n6901), .A2(n_T_635[37]), .Y(n6226) );
  NAND4X0_LVT U7620 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .Y(
        n_T_702[37]) );
  AO22X1_LVT U7621 ( .A1(n6856), .A2(io_fpu_toint_data[38]), .A3(n6855), .A4(
        n_T_918[38]), .Y(n6230) );
  AO21X1_LVT U7622 ( .A1(mem_br_target[38]), .A2(n6249), .A3(n6230), .Y(N636)
         );
  AO22X1_LVT U7623 ( .A1(n3851), .A2(io_dmem_resp_bits_data[38]), .A3(n3848), 
        .A4(io_imem_sfence_bits_addr[38]), .Y(n6231) );
  AO21X1_LVT U7624 ( .A1(n3856), .A2(div_io_resp_bits_data[38]), .A3(n6231), 
        .Y(n6232) );
  AO22X1_LVT U7625 ( .A1(n3806), .A2(n_T_427[230]), .A3(n_T_427[166]), .A4(
        n2862), .Y(n6244) );
  AO22X1_LVT U7626 ( .A1(n2869), .A2(n_T_427[614]), .A3(n_T_427[102]), .A4(
        n3832), .Y(n6243) );
  AO22X1_LVT U7627 ( .A1(n3913), .A2(n_T_427[38]), .A3(n_T_427[294]), .A4(
        n3809), .Y(n6242) );
  AO22X1_LVT U7628 ( .A1(n_T_427[933]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[486]), .Y(n6236) );
  AO22X1_LVT U7629 ( .A1(n6765), .A2(n_T_427[741]), .A3(n3865), .A4(
        n_T_427[422]), .Y(n6235) );
  AO22X1_LVT U7630 ( .A1(n_T_427[678]), .A2(n3861), .A3(n3866), .A4(
        n_T_427[358]), .Y(n6234) );
  AO22X1_LVT U7631 ( .A1(n3813), .A2(n_T_427[805]), .A3(n_T_427[869]), .A4(
        n3874), .Y(n6233) );
  NOR4X1_LVT U7632 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .Y(n6237)
         );
  OA22X1_LVT U7633 ( .A1(n3098), .A2(n3596), .A3(n3877), .A4(n6237), .Y(n6240)
         );
  NAND2X0_LVT U7634 ( .A1(n_T_427[550]), .A2(n2850), .Y(n6239) );
  NAND2X0_LVT U7635 ( .A1(n6240), .A2(n6239), .Y(n6241) );
  NAND2X0_LVT U7636 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[38]), .Y(n6248) );
  NAND2X0_LVT U7637 ( .A1(n6899), .A2(n_T_918[38]), .Y(n6247) );
  NAND2X0_LVT U7638 ( .A1(n6900), .A2(io_imem_sfence_bits_addr[38]), .Y(n6246)
         );
  NAND2X0_LVT U7639 ( .A1(n3243), .A2(n_T_635[38]), .Y(n6245) );
  NAND4X0_LVT U7640 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .Y(
        n_T_702[38]) );
  AOI22X1_LVT U7641 ( .A1(n6856), .A2(io_fpu_toint_data[39]), .A3(n6855), .A4(
        n_T_918[39]), .Y(n6250) );
  NAND2X0_LVT U7642 ( .A1(n6857), .A2(n6250), .Y(N637) );
  NAND2X0_LVT U7643 ( .A1(csr_io_rw_rdata[39]), .A2(n3845), .Y(n6253) );
  AOI22X1_LVT U7644 ( .A1(n3853), .A2(io_dmem_resp_bits_data[39]), .A3(n3846), 
        .A4(n_T_1165[39]), .Y(n6252) );
  NAND2X0_LVT U7645 ( .A1(div_io_resp_bits_data[39]), .A2(n3858), .Y(n6251) );
  NAND3X0_LVT U7646 ( .A1(n6253), .A2(n6252), .A3(n6251), .Y(
        n_T_427__T_1136_data[39]) );
  AOI22X1_LVT U7647 ( .A1(n3870), .A2(n_T_427[551]), .A3(n_T_427[615]), .A4(
        n3795), .Y(n6257) );
  AOI22X1_LVT U7648 ( .A1(n6871), .A2(n_T_427[870]), .A3(n6838), .A4(
        n_T_427[39]), .Y(n6256) );
  AOI22X1_LVT U7649 ( .A1(n3865), .A2(n_T_427[423]), .A3(n_T_427[742]), .A4(
        n3804), .Y(n6255) );
  OA22X1_LVT U7650 ( .A1(n3523), .A2(n6423), .A3(n3179), .A4(n3083), .Y(n6254)
         );
  NAND4X0_LVT U7651 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .Y(n6258) );
  AO22X1_LVT U7652 ( .A1(n3925), .A2(n_T_427[1510]), .A3(n_T_427[1382]), .A4(
        n3919), .Y(n6262) );
  AO22X1_LVT U7653 ( .A1(n3935), .A2(n_T_427[1446]), .A3(n_T_427[1318]), .A4(
        n3929), .Y(n6261) );
  AO22X1_LVT U7654 ( .A1(n3945), .A2(n_T_427[1190]), .A3(n_T_427[1254]), .A4(
        n3939), .Y(n6260) );
  AO22X1_LVT U7655 ( .A1(n3955), .A2(n_T_427[1126]), .A3(n_T_427[998]), .A4(
        n3949), .Y(n6259) );
  NOR4X1_LVT U7656 ( .A1(n6262), .A2(n6261), .A3(n6260), .A4(n6259), .Y(n6269)
         );
  AO22X1_LVT U7657 ( .A1(n2860), .A2(n_T_427[806]), .A3(n_T_427[103]), .A4(
        n3832), .Y(n6266) );
  AO22X1_LVT U7658 ( .A1(n3901), .A2(n_T_427[1062]), .A3(n_T_427[934]), .A4(
        n3895), .Y(n6265) );
  AO22X1_LVT U7659 ( .A1(n3910), .A2(n_T_427[487]), .A3(n_T_427[167]), .A4(
        n2863), .Y(n6264) );
  AO22X1_LVT U7660 ( .A1(n2857), .A2(n_T_427[359]), .A3(n_T_427[295]), .A4(
        n3809), .Y(n6263) );
  NOR4X1_LVT U7661 ( .A1(n6266), .A2(n6265), .A3(n6264), .A4(n6263), .Y(n6268)
         );
  NAND2X0_LVT U7662 ( .A1(n3957), .A2(n4424), .Y(n6267) );
  NAND4X0_LVT U7663 ( .A1(n6269), .A2(n6270), .A3(n6268), .A4(n6267), .Y(
        id_rs_1[39]) );
  NAND2X0_LVT U7664 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[39]), .Y(n6274) );
  NAND2X0_LVT U7665 ( .A1(n6899), .A2(n_T_918[39]), .Y(n6273) );
  NAND2X0_LVT U7666 ( .A1(n6900), .A2(n_T_1165[39]), .Y(n6272) );
  NAND2X0_LVT U7667 ( .A1(n6901), .A2(n_T_635[39]), .Y(n6271) );
  NAND4X0_LVT U7668 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6271), .Y(
        n_T_702[39]) );
  AOI22X1_LVT U7669 ( .A1(n6856), .A2(io_fpu_toint_data[40]), .A3(n6855), .A4(
        n_T_918[40]), .Y(n6275) );
  NAND2X0_LVT U7670 ( .A1(n6857), .A2(n6275), .Y(N638) );
  NAND2X0_LVT U7671 ( .A1(csr_io_rw_rdata[40]), .A2(n3845), .Y(n6278) );
  AOI22X1_LVT U7672 ( .A1(n3853), .A2(io_dmem_resp_bits_data[40]), .A3(n3846), 
        .A4(n_T_1165[40]), .Y(n6277) );
  NAND2X0_LVT U7673 ( .A1(div_io_resp_bits_data[40]), .A2(n3858), .Y(n6276) );
  NAND3X0_LVT U7674 ( .A1(n6278), .A2(n6277), .A3(n6276), .Y(
        n_T_427__T_1136_data[40]) );
  AO22X1_LVT U7675 ( .A1(n2861), .A2(n_T_427[807]), .A3(n_T_427[168]), .A4(
        n2863), .Y(n6280) );
  AO22X1_LVT U7676 ( .A1(n3817), .A2(n_T_427[360]), .A3(n_T_427[680]), .A4(
        n6812), .Y(n6279) );
  AO22X1_LVT U7677 ( .A1(n6765), .A2(n_T_427[743]), .A3(n3865), .A4(
        n_T_427[424]), .Y(n6284) );
  AO22X1_LVT U7678 ( .A1(n3869), .A2(n_T_427[552]), .A3(n_T_427[616]), .A4(
        n3795), .Y(n6283) );
  AO22X1_LVT U7679 ( .A1(n3837), .A2(n_T_427[488]), .A3(n3873), .A4(
        n_T_427[296]), .Y(n6282) );
  AO22X1_LVT U7680 ( .A1(n_T_427[871]), .A2(n6871), .A3(n3839), .A4(
        n_T_427[40]), .Y(n6281) );
  NOR4X1_LVT U7681 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .Y(n6285)
         );
  OA22X1_LVT U7682 ( .A1(n3551), .A2(n3881), .A3(n3877), .A4(n6285), .Y(n6288)
         );
  NAND2X0_LVT U7683 ( .A1(n3958), .A2(n4427), .Y(n6287) );
  OA22X1_LVT U7684 ( .A1(n3147), .A2(n3803), .A3(n3499), .A4(n3800), .Y(n6286)
         );
  AND3X1_LVT U7685 ( .A1(n6288), .A2(n6287), .A3(n6286), .Y(n6289) );
  NAND4X0_LVT U7686 ( .A1(n6291), .A2(n6292), .A3(n6290), .A4(n6289), .Y(
        id_rs_1[40]) );
  NAND2X0_LVT U7687 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[40]), .Y(n6296) );
  NAND2X0_LVT U7688 ( .A1(n6899), .A2(n_T_918[40]), .Y(n6295) );
  NAND2X0_LVT U7689 ( .A1(n6900), .A2(n_T_1165[40]), .Y(n6294) );
  NAND2X0_LVT U7690 ( .A1(n3243), .A2(n_T_635[40]), .Y(n6293) );
  NAND4X0_LVT U7691 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .Y(
        n_T_702[40]) );
  AOI22X1_LVT U7692 ( .A1(n6856), .A2(io_fpu_toint_data[41]), .A3(n6855), .A4(
        n_T_918[41]), .Y(n6297) );
  NAND2X0_LVT U7693 ( .A1(n6857), .A2(n6297), .Y(N639) );
  AO22X1_LVT U7694 ( .A1(n3851), .A2(io_dmem_resp_bits_data[41]), .A3(n3848), 
        .A4(n_T_1165[41]), .Y(n6298) );
  AO21X1_LVT U7695 ( .A1(n3856), .A2(div_io_resp_bits_data[41]), .A3(n6298), 
        .Y(n6299) );
  AO21X1_LVT U7696 ( .A1(n3842), .A2(csr_io_rw_rdata[41]), .A3(n6299), .Y(
        n_T_427__T_1136_data[41]) );
  AO22X1_LVT U7697 ( .A1(n3945), .A2(n_T_427[1192]), .A3(n_T_427[1256]), .A4(
        n3939), .Y(n6303) );
  AO22X1_LVT U7698 ( .A1(n3955), .A2(n_T_427[1128]), .A3(n_T_427[1000]), .A4(
        n3949), .Y(n6302) );
  AO22X1_LVT U7699 ( .A1(n3901), .A2(n_T_427[1064]), .A3(n_T_427[233]), .A4(
        n6773), .Y(n6301) );
  AO22X1_LVT U7700 ( .A1(n2861), .A2(n_T_427[808]), .A3(n_T_427[489]), .A4(
        n3911), .Y(n6300) );
  NOR4X1_LVT U7701 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .Y(n6316)
         );
  AO22X1_LVT U7702 ( .A1(n2833), .A2(n_T_427[872]), .A3(n_T_427[169]), .A4(
        n2862), .Y(n6305) );
  AO22X1_LVT U7703 ( .A1(n3809), .A2(n_T_427[297]), .A3(n_T_427[681]), .A4(
        n3821), .Y(n6304) );
  NOR2X0_LVT U7704 ( .A1(n6305), .A2(n6304), .Y(n6315) );
  AO22X1_LVT U7705 ( .A1(n3869), .A2(n_T_427[553]), .A3(n_T_427[617]), .A4(
        n3795), .Y(n6309) );
  AO22X1_LVT U7706 ( .A1(n_T_427[744]), .A2(n3804), .A3(n6866), .A4(
        n_T_427[105]), .Y(n6308) );
  AO22X1_LVT U7707 ( .A1(n6867), .A2(n_T_427[425]), .A3(n3866), .A4(
        n_T_427[361]), .Y(n6307) );
  AO22X1_LVT U7708 ( .A1(n_T_427[936]), .A2(n6794), .A3(n3839), .A4(
        n_T_427[41]), .Y(n6306) );
  NOR4X1_LVT U7709 ( .A1(n6309), .A2(n6308), .A3(n6307), .A4(n6306), .Y(n6310)
         );
  OA22X1_LVT U7710 ( .A1(n3552), .A2(n3881), .A3(n1993), .A4(n6310), .Y(n6313)
         );
  OA22X1_LVT U7711 ( .A1(n3148), .A2(n3803), .A3(n3500), .A4(n3799), .Y(n6312)
         );
  NAND2X0_LVT U7712 ( .A1(n4430), .A2(n3959), .Y(n6311) );
  AND3X1_LVT U7713 ( .A1(n6313), .A2(n6312), .A3(n6311), .Y(n6314) );
  NAND4X0_LVT U7714 ( .A1(n6316), .A2(n6317), .A3(n6315), .A4(n6314), .Y(
        id_rs_1[41]) );
  NAND2X0_LVT U7715 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[41]), .Y(n6321) );
  NAND2X0_LVT U7716 ( .A1(n6899), .A2(n_T_918[41]), .Y(n6320) );
  NAND2X0_LVT U7717 ( .A1(n6900), .A2(n_T_1165[41]), .Y(n6319) );
  NAND2X0_LVT U7718 ( .A1(n6901), .A2(n_T_635[41]), .Y(n6318) );
  NAND4X0_LVT U7719 ( .A1(n6321), .A2(n6320), .A3(n6319), .A4(n6318), .Y(
        n_T_702[41]) );
  AOI22X1_LVT U7720 ( .A1(n6856), .A2(io_fpu_toint_data[42]), .A3(n6855), .A4(
        n_T_918[42]), .Y(n6322) );
  NAND2X0_LVT U7721 ( .A1(n6857), .A2(n6322), .Y(N640) );
  AO22X1_LVT U7722 ( .A1(n3851), .A2(io_dmem_resp_bits_data[42]), .A3(n3848), 
        .A4(n_T_1165[42]), .Y(n6323) );
  AO21X1_LVT U7723 ( .A1(n3857), .A2(div_io_resp_bits_data[42]), .A3(n6323), 
        .Y(n6324) );
  AO21X1_LVT U7724 ( .A1(n3842), .A2(csr_io_rw_rdata[42]), .A3(n6324), .Y(
        n_T_427__T_1136_data[42]) );
  AO22X1_LVT U7725 ( .A1(n3945), .A2(n_T_427[1193]), .A3(n_T_427[1257]), .A4(
        n3940), .Y(n6328) );
  AO22X1_LVT U7726 ( .A1(n3955), .A2(n_T_427[1129]), .A3(n_T_427[1001]), .A4(
        n3950), .Y(n6327) );
  AO22X1_LVT U7727 ( .A1(n3901), .A2(n_T_427[1065]), .A3(n_T_427[234]), .A4(
        n6773), .Y(n6326) );
  AO22X1_LVT U7728 ( .A1(n2865), .A2(n_T_427[426]), .A3(n_T_427[745]), .A4(
        n3904), .Y(n6325) );
  NOR4X1_LVT U7729 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .Y(n6341)
         );
  AO22X1_LVT U7730 ( .A1(n3912), .A2(n_T_427[490]), .A3(n_T_427[170]), .A4(
        n3908), .Y(n6330) );
  AO22X1_LVT U7731 ( .A1(n2833), .A2(n_T_427[873]), .A3(n_T_427[298]), .A4(
        n3809), .Y(n6329) );
  AO22X1_LVT U7732 ( .A1(n_T_427[937]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[618]), .Y(n6334) );
  AO22X1_LVT U7733 ( .A1(n_T_427[682]), .A2(n3861), .A3(n6866), .A4(
        n_T_427[106]), .Y(n6333) );
  AO22X1_LVT U7734 ( .A1(n_T_427[554]), .A2(n3869), .A3(n3866), .A4(
        n_T_427[362]), .Y(n6332) );
  AO22X1_LVT U7735 ( .A1(n_T_427[809]), .A2(n3813), .A3(n3839), .A4(
        n_T_427[42]), .Y(n6331) );
  NOR4X1_LVT U7736 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .Y(n6335)
         );
  OA22X1_LVT U7737 ( .A1(n3553), .A2(n3881), .A3(n1993), .A4(n6335), .Y(n6338)
         );
  OA22X1_LVT U7738 ( .A1(n3149), .A2(n3803), .A3(n3501), .A4(n3799), .Y(n6337)
         );
  NAND2X0_LVT U7739 ( .A1(n4433), .A2(n3959), .Y(n6336) );
  AND3X1_LVT U7740 ( .A1(n6338), .A2(n6337), .A3(n6336), .Y(n6339) );
  NAND4X0_LVT U7741 ( .A1(n6341), .A2(n6342), .A3(n6340), .A4(n6339), .Y(
        id_rs_1[42]) );
  NAND2X0_LVT U7742 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[42]), .Y(n6346) );
  NAND2X0_LVT U7743 ( .A1(n6899), .A2(n_T_918[42]), .Y(n6345) );
  NAND2X0_LVT U7744 ( .A1(n6900), .A2(n_T_1165[42]), .Y(n6344) );
  NAND2X0_LVT U7745 ( .A1(n3243), .A2(n_T_635[42]), .Y(n6343) );
  NAND4X0_LVT U7746 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .Y(
        n_T_702[42]) );
  AOI22X1_LVT U7747 ( .A1(n6856), .A2(io_fpu_toint_data[43]), .A3(n6855), .A4(
        n_T_918[43]), .Y(n6347) );
  NAND2X0_LVT U7748 ( .A1(n6857), .A2(n6347), .Y(N641) );
  AO22X1_LVT U7749 ( .A1(n3851), .A2(io_dmem_resp_bits_data[43]), .A3(n3848), 
        .A4(n_T_1165[43]), .Y(n6348) );
  AO21X1_LVT U7750 ( .A1(n3857), .A2(div_io_resp_bits_data[43]), .A3(n6348), 
        .Y(n6349) );
  AO21X1_LVT U7751 ( .A1(n3842), .A2(csr_io_rw_rdata[43]), .A3(n6349), .Y(
        n_T_427__T_1136_data[43]) );
  AO22X1_LVT U7752 ( .A1(n3915), .A2(n_T_427[619]), .A3(n_T_427[171]), .A4(
        n3909), .Y(n6351) );
  AO22X1_LVT U7753 ( .A1(n3810), .A2(n_T_427[299]), .A3(n_T_427[683]), .A4(
        n2829), .Y(n6350) );
  NOR2X0_LVT U7754 ( .A1(n6351), .A2(n6350), .Y(n6361) );
  AO22X1_LVT U7755 ( .A1(n3869), .A2(n_T_427[555]), .A3(n_T_427[491]), .A4(
        n3836), .Y(n6355) );
  AO22X1_LVT U7756 ( .A1(n6867), .A2(n_T_427[427]), .A3(n6866), .A4(
        n_T_427[107]), .Y(n6354) );
  AO22X1_LVT U7757 ( .A1(n3860), .A2(n_T_427[235]), .A3(n3866), .A4(
        n_T_427[363]), .Y(n6353) );
  AO22X1_LVT U7758 ( .A1(n_T_427[874]), .A2(n6871), .A3(n3839), .A4(
        n_T_427[43]), .Y(n6352) );
  NOR4X1_LVT U7759 ( .A1(n6355), .A2(n6354), .A3(n6353), .A4(n6352), .Y(n6356)
         );
  OA22X1_LVT U7760 ( .A1(n3554), .A2(n3881), .A3(n3877), .A4(n6356), .Y(n6359)
         );
  OA22X1_LVT U7761 ( .A1(n3150), .A2(n3803), .A3(n3502), .A4(n3799), .Y(n6358)
         );
  NAND2X0_LVT U7762 ( .A1(n4436), .A2(n3959), .Y(n6357) );
  AND3X1_LVT U7763 ( .A1(n6359), .A2(n6358), .A3(n6357), .Y(n6360) );
  NAND4X0_LVT U7764 ( .A1(n6362), .A2(n6363), .A3(n6361), .A4(n6360), .Y(
        id_rs_1[43]) );
  NAND2X0_LVT U7765 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[43]), .Y(n6367) );
  NAND2X0_LVT U7766 ( .A1(n6899), .A2(n_T_918[43]), .Y(n6366) );
  NAND2X0_LVT U7767 ( .A1(n6900), .A2(n_T_1165[43]), .Y(n6365) );
  NAND2X0_LVT U7768 ( .A1(n3243), .A2(n_T_635[43]), .Y(n6364) );
  NAND4X0_LVT U7769 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .Y(
        n_T_702[43]) );
  AOI22X1_LVT U7770 ( .A1(n6856), .A2(io_fpu_toint_data[44]), .A3(n6855), .A4(
        n_T_918[44]), .Y(n6368) );
  NAND2X0_LVT U7771 ( .A1(n6857), .A2(n6368), .Y(N642) );
  NAND2X0_LVT U7772 ( .A1(csr_io_rw_rdata[44]), .A2(n3845), .Y(n6371) );
  AOI22X1_LVT U7773 ( .A1(n3853), .A2(io_dmem_resp_bits_data[44]), .A3(n3846), 
        .A4(n_T_1165[44]), .Y(n6370) );
  NAND2X0_LVT U7774 ( .A1(div_io_resp_bits_data[44]), .A2(n3858), .Y(n6369) );
  NAND3X0_LVT U7775 ( .A1(n6371), .A2(n6370), .A3(n6369), .Y(
        n_T_427__T_1136_data[44]) );
  AOI22X1_LVT U7776 ( .A1(n3797), .A2(n_T_427[620]), .A3(n3867), .A4(
        n_T_427[364]), .Y(n6375) );
  AOI22X1_LVT U7777 ( .A1(n6871), .A2(n_T_427[875]), .A3(n3871), .A4(
        n_T_427[300]), .Y(n6374) );
  AOI22X1_LVT U7778 ( .A1(n6765), .A2(n_T_427[747]), .A3(n3864), .A4(
        n_T_427[108]), .Y(n6373) );
  AOI22X1_LVT U7779 ( .A1(n3863), .A2(n_T_427[684]), .A3(n3865), .A4(
        n_T_427[428]), .Y(n6372) );
  NAND4X0_LVT U7780 ( .A1(n6375), .A2(n6374), .A3(n6373), .A4(n6372), .Y(n6376) );
  AO22X1_LVT U7781 ( .A1(n3901), .A2(n_T_427[1067]), .A3(n_T_427[236]), .A4(
        n3807), .Y(n6380) );
  AO22X1_LVT U7782 ( .A1(n2860), .A2(n_T_427[811]), .A3(n_T_427[939]), .A4(
        n3895), .Y(n6379) );
  AO22X1_LVT U7783 ( .A1(n3912), .A2(n_T_427[492]), .A3(n_T_427[172]), .A4(
        n3909), .Y(n6378) );
  AO22X1_LVT U7784 ( .A1(n3818), .A2(n_T_427[556]), .A3(n_T_427[44]), .A4(
        n3914), .Y(n6377) );
  NOR4X1_LVT U7785 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .Y(n6387)
         );
  AO22X1_LVT U7786 ( .A1(n3925), .A2(n_T_427[1515]), .A3(n_T_427[1387]), .A4(
        n3920), .Y(n6384) );
  AO22X1_LVT U7787 ( .A1(n3935), .A2(n_T_427[1451]), .A3(n_T_427[1323]), .A4(
        n3930), .Y(n6383) );
  AO22X1_LVT U7788 ( .A1(n3945), .A2(n_T_427[1195]), .A3(n_T_427[1259]), .A4(
        n3940), .Y(n6382) );
  AO22X1_LVT U7789 ( .A1(n3955), .A2(n_T_427[1131]), .A3(n_T_427[1003]), .A4(
        n3950), .Y(n6381) );
  NOR4X1_LVT U7790 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .Y(n6386)
         );
  NAND2X0_LVT U7791 ( .A1(n3957), .A2(n4439), .Y(n6385) );
  NAND4X0_LVT U7792 ( .A1(n6387), .A2(n6388), .A3(n6386), .A4(n6385), .Y(
        id_rs_1[44]) );
  NAND2X0_LVT U7793 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[44]), .Y(n6392) );
  NAND2X0_LVT U7794 ( .A1(n6899), .A2(n_T_918[44]), .Y(n6391) );
  NAND2X0_LVT U7795 ( .A1(n6900), .A2(n_T_1165[44]), .Y(n6390) );
  NAND2X0_LVT U7796 ( .A1(n6901), .A2(n_T_635[44]), .Y(n6389) );
  NAND4X0_LVT U7797 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .Y(
        n_T_702[44]) );
  AOI22X1_LVT U7798 ( .A1(n6856), .A2(io_fpu_toint_data[45]), .A3(n6855), .A4(
        n_T_918[45]), .Y(n6393) );
  NAND2X0_LVT U7799 ( .A1(n6857), .A2(n6393), .Y(N643) );
  AO22X1_LVT U7800 ( .A1(n3851), .A2(io_dmem_resp_bits_data[45]), .A3(n3848), 
        .A4(n_T_1165[45]), .Y(n6394) );
  AO21X1_LVT U7801 ( .A1(n3857), .A2(div_io_resp_bits_data[45]), .A3(n6394), 
        .Y(n6395) );
  AO21X1_LVT U7802 ( .A1(n3842), .A2(csr_io_rw_rdata[45]), .A3(n6395), .Y(
        n_T_427__T_1136_data[45]) );
  AO22X1_LVT U7803 ( .A1(n3818), .A2(n_T_427[557]), .A3(n_T_427[45]), .A4(
        n2826), .Y(n6397) );
  AO22X1_LVT U7804 ( .A1(n3822), .A2(n_T_427[876]), .A3(n_T_427[685]), .A4(
        n3820), .Y(n6396) );
  NOR2X0_LVT U7805 ( .A1(n6397), .A2(n6396), .Y(n6407) );
  AO22X1_LVT U7806 ( .A1(n3815), .A2(n_T_427[173]), .A3(n_T_427[812]), .A4(
        n3812), .Y(n6401) );
  AO22X1_LVT U7807 ( .A1(n6765), .A2(n_T_427[748]), .A3(n3860), .A4(
        n_T_427[237]), .Y(n6400) );
  AO22X1_LVT U7808 ( .A1(n_T_427[621]), .A2(n3796), .A3(n3866), .A4(
        n_T_427[365]), .Y(n6399) );
  AO22X1_LVT U7809 ( .A1(n3838), .A2(n_T_427[493]), .A3(n3873), .A4(
        n_T_427[301]), .Y(n6398) );
  NOR4X1_LVT U7810 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .Y(n6402)
         );
  OA22X1_LVT U7811 ( .A1(n3151), .A2(n3803), .A3(n3503), .A4(n3800), .Y(n6404)
         );
  NAND2X0_LVT U7812 ( .A1(n4442), .A2(n3959), .Y(n6403) );
  AND3X1_LVT U7813 ( .A1(n6405), .A2(n6404), .A3(n6403), .Y(n6406) );
  NAND4X0_LVT U7814 ( .A1(n6408), .A2(n6409), .A3(n6407), .A4(n6406), .Y(
        id_rs_1[45]) );
  NAND2X0_LVT U7815 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[45]), .Y(n6413) );
  NAND2X0_LVT U7816 ( .A1(n6899), .A2(n_T_918[45]), .Y(n6412) );
  NAND2X0_LVT U7817 ( .A1(n6900), .A2(n_T_1165[45]), .Y(n6411) );
  NAND2X0_LVT U7818 ( .A1(n3243), .A2(n_T_635[45]), .Y(n6410) );
  NAND4X0_LVT U7819 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .Y(
        n_T_702[45]) );
  AOI22X1_LVT U7820 ( .A1(n6856), .A2(io_fpu_toint_data[46]), .A3(n6855), .A4(
        n_T_918[46]), .Y(n6414) );
  NAND2X0_LVT U7821 ( .A1(n6857), .A2(n6414), .Y(N644) );
  NAND2X0_LVT U7822 ( .A1(csr_io_rw_rdata[46]), .A2(n3845), .Y(n6417) );
  AOI22X1_LVT U7823 ( .A1(n3853), .A2(io_dmem_resp_bits_data[46]), .A3(n3847), 
        .A4(n_T_1165[46]), .Y(n6416) );
  NAND2X0_LVT U7824 ( .A1(div_io_resp_bits_data[46]), .A2(n3858), .Y(n6415) );
  NAND3X0_LVT U7825 ( .A1(n6417), .A2(n6416), .A3(n6415), .Y(
        n_T_427__T_1136_data[46]) );
  AO22X1_LVT U7826 ( .A1(n3925), .A2(n_T_427[1517]), .A3(n_T_427[1389]), .A4(
        n3920), .Y(n6421) );
  AO22X1_LVT U7827 ( .A1(n3935), .A2(n_T_427[1453]), .A3(n_T_427[1325]), .A4(
        n3930), .Y(n6420) );
  AO22X1_LVT U7828 ( .A1(n3945), .A2(n_T_427[1197]), .A3(n_T_427[1261]), .A4(
        n3940), .Y(n6419) );
  AO22X1_LVT U7829 ( .A1(n3955), .A2(n_T_427[1133]), .A3(n_T_427[1005]), .A4(
        n3950), .Y(n6418) );
  NOR4X1_LVT U7830 ( .A1(n6421), .A2(n6420), .A3(n6419), .A4(n6418), .Y(n6436)
         );
  AOI22X1_LVT U7831 ( .A1(n3870), .A2(n_T_427[558]), .A3(n6868), .A4(
        n_T_427[366]), .Y(n6427) );
  AOI22X1_LVT U7832 ( .A1(n3814), .A2(n_T_427[813]), .A3(n_T_427[877]), .A4(
        n3875), .Y(n6426) );
  OA22X1_LVT U7833 ( .A1(n3522), .A2(n6423), .A3(n3176), .A4(n6422), .Y(n6425)
         );
  AOI22X1_LVT U7834 ( .A1(n_T_427[941]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[622]), .Y(n6424) );
  NAND4X0_LVT U7835 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .Y(n6428) );
  AO22X1_LVT U7836 ( .A1(n2864), .A2(n_T_427[430]), .A3(n_T_427[1069]), .A4(
        n3898), .Y(n6432) );
  AO22X1_LVT U7837 ( .A1(n3911), .A2(n_T_427[494]), .A3(n_T_427[749]), .A4(
        n3905), .Y(n6431) );
  AO22X1_LVT U7838 ( .A1(n2879), .A2(n_T_427[46]), .A3(n_T_427[174]), .A4(
        n2862), .Y(n6430) );
  AO22X1_LVT U7839 ( .A1(n3810), .A2(n_T_427[302]), .A3(n_T_427[686]), .A4(
        n2829), .Y(n6429) );
  NOR4X1_LVT U7840 ( .A1(n6432), .A2(n6431), .A3(n6430), .A4(n6429), .Y(n6434)
         );
  NAND2X0_LVT U7841 ( .A1(n3957), .A2(n4445), .Y(n6433) );
  NAND4X0_LVT U7842 ( .A1(n6436), .A2(n6435), .A3(n6434), .A4(n6433), .Y(
        id_rs_1[46]) );
  NAND2X0_LVT U7843 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[46]), .Y(n6440) );
  NAND2X0_LVT U7844 ( .A1(n6899), .A2(n_T_918[46]), .Y(n6439) );
  NAND2X0_LVT U7845 ( .A1(n6900), .A2(n_T_1165[46]), .Y(n6438) );
  NAND2X0_LVT U7846 ( .A1(n6901), .A2(n_T_635[46]), .Y(n6437) );
  NAND4X0_LVT U7847 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .Y(
        n_T_702[46]) );
  AOI22X1_LVT U7848 ( .A1(n6856), .A2(io_fpu_toint_data[47]), .A3(n6855), .A4(
        n_T_918[47]), .Y(n6441) );
  NAND2X0_LVT U7849 ( .A1(n6857), .A2(n6441), .Y(N645) );
  NAND2X0_LVT U7850 ( .A1(csr_io_rw_rdata[47]), .A2(n3845), .Y(n6444) );
  AOI22X1_LVT U7851 ( .A1(n3853), .A2(io_dmem_resp_bits_data[47]), .A3(n3847), 
        .A4(n_T_1165[47]), .Y(n6443) );
  NAND2X0_LVT U7852 ( .A1(div_io_resp_bits_data[47]), .A2(n3858), .Y(n6442) );
  NAND3X0_LVT U7853 ( .A1(n6444), .A2(n6443), .A3(n6442), .Y(
        n_T_427__T_1136_data[47]) );
  AO22X1_LVT U7854 ( .A1(n3817), .A2(n_T_427[367]), .A3(n_T_427[495]), .A4(
        n3912), .Y(n6446) );
  AO22X1_LVT U7855 ( .A1(n3916), .A2(n_T_427[623]), .A3(n_T_427[878]), .A4(
        n3822), .Y(n6445) );
  NOR2X0_LVT U7856 ( .A1(n6446), .A2(n6445), .Y(n6456) );
  AO22X1_LVT U7857 ( .A1(n_T_427[942]), .A2(n6794), .A3(n3868), .A4(
        n_T_427[559]), .Y(n6450) );
  AO22X1_LVT U7858 ( .A1(n_T_427[687]), .A2(n3861), .A3(n6866), .A4(
        n_T_427[111]), .Y(n6449) );
  AO22X1_LVT U7859 ( .A1(n_T_427[814]), .A2(n3813), .A3(n3873), .A4(
        n_T_427[303]), .Y(n6448) );
  AO22X1_LVT U7860 ( .A1(n3815), .A2(n_T_427[175]), .A3(n3839), .A4(
        n_T_427[47]), .Y(n6447) );
  NOR4X1_LVT U7861 ( .A1(n6450), .A2(n6449), .A3(n6448), .A4(n6447), .Y(n6451)
         );
  OA22X1_LVT U7862 ( .A1(n3556), .A2(n3882), .A3(n3877), .A4(n6451), .Y(n6454)
         );
  NAND2X0_LVT U7863 ( .A1(n3957), .A2(n4448), .Y(n6453) );
  OA22X1_LVT U7864 ( .A1(n3152), .A2(n3803), .A3(n3504), .A4(n3800), .Y(n6452)
         );
  AND3X1_LVT U7865 ( .A1(n6454), .A2(n6453), .A3(n6452), .Y(n6455) );
  NAND4X0_LVT U7866 ( .A1(n6457), .A2(n6458), .A3(n6456), .A4(n6455), .Y(
        id_rs_1[47]) );
  NAND2X0_LVT U7867 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[47]), .Y(n6462) );
  NAND2X0_LVT U7868 ( .A1(n6899), .A2(n_T_918[47]), .Y(n6461) );
  NAND2X0_LVT U7869 ( .A1(n6900), .A2(n_T_1165[47]), .Y(n6460) );
  NAND2X0_LVT U7870 ( .A1(n3243), .A2(n_T_635[47]), .Y(n6459) );
  NAND4X0_LVT U7871 ( .A1(n6462), .A2(n6461), .A3(n6460), .A4(n6459), .Y(
        n_T_702[47]) );
  NAND2X0_LVT U7872 ( .A1(csr_io_rw_rdata[48]), .A2(n3845), .Y(n6465) );
  AOI22X1_LVT U7873 ( .A1(n3853), .A2(io_dmem_resp_bits_data[48]), .A3(n3847), 
        .A4(n_T_1165[48]), .Y(n6464) );
  NAND2X0_LVT U7874 ( .A1(div_io_resp_bits_data[48]), .A2(n3858), .Y(n6463) );
  NAND3X0_LVT U7875 ( .A1(n6465), .A2(n6464), .A3(n6463), .Y(
        n_T_427__T_1136_data[48]) );
  AO22X1_LVT U7876 ( .A1(n3828), .A2(n_T_427[1836]), .A3(n_T_427[1711]), .A4(
        n3824), .Y(n6469) );
  AO22X1_LVT U7877 ( .A1(n3893), .A2(n_T_427[1583]), .A3(n_T_427[1647]), .A4(
        n3888), .Y(n6468) );
  AO22X1_LVT U7878 ( .A1(n3925), .A2(n_T_427[1519]), .A3(n_T_427[1391]), .A4(
        n3920), .Y(n6467) );
  AO22X1_LVT U7879 ( .A1(n3935), .A2(n_T_427[1455]), .A3(n_T_427[1327]), .A4(
        n3930), .Y(n6466) );
  NOR4X1_LVT U7880 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .Y(n6483)
         );
  AO22X1_LVT U7881 ( .A1(n3911), .A2(n_T_427[496]), .A3(n_T_427[751]), .A4(
        n3903), .Y(n6471) );
  AO22X1_LVT U7882 ( .A1(n3915), .A2(n_T_427[624]), .A3(n_T_427[688]), .A4(
        n2829), .Y(n6470) );
  NOR2X0_LVT U7883 ( .A1(n6471), .A2(n6470), .Y(n6481) );
  AO22X1_LVT U7884 ( .A1(n3813), .A2(n_T_427[815]), .A3(n_T_427[879]), .A4(
        n3874), .Y(n6475) );
  AO22X1_LVT U7885 ( .A1(n_T_427[560]), .A2(n3869), .A3(n3873), .A4(
        n_T_427[304]), .Y(n6474) );
  AO22X1_LVT U7886 ( .A1(n3815), .A2(n_T_427[176]), .A3(n3839), .A4(
        n_T_427[48]), .Y(n6473) );
  AO22X1_LVT U7887 ( .A1(n6866), .A2(n_T_427[112]), .A3(n3867), .A4(
        n_T_427[368]), .Y(n6472) );
  NOR4X1_LVT U7888 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .Y(n6476)
         );
  OA22X1_LVT U7889 ( .A1(n3557), .A2(n3882), .A3(n1993), .A4(n6476), .Y(n6479)
         );
  NAND2X0_LVT U7890 ( .A1(n3957), .A2(n4451), .Y(n6478) );
  OA22X1_LVT U7891 ( .A1(n3153), .A2(n3803), .A3(n3505), .A4(n3800), .Y(n6477)
         );
  AND3X1_LVT U7892 ( .A1(n6479), .A2(n6478), .A3(n6477), .Y(n6480) );
  NAND4X0_LVT U7893 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .Y(
        id_rs_1[48]) );
  NAND2X0_LVT U7894 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[48]), .Y(n6487) );
  NAND2X0_LVT U7895 ( .A1(n6899), .A2(n_T_918[48]), .Y(n6486) );
  NAND2X0_LVT U7896 ( .A1(n6900), .A2(n_T_1165[48]), .Y(n6485) );
  NAND2X0_LVT U7897 ( .A1(n3243), .A2(n_T_635[48]), .Y(n6484) );
  NAND4X0_LVT U7898 ( .A1(n6487), .A2(n6486), .A3(n6485), .A4(n6484), .Y(
        n_T_702[48]) );
  AO22X1_LVT U7899 ( .A1(n6860), .A2(io_dmem_resp_bits_data[49]), .A3(n3848), 
        .A4(n_T_1165[49]), .Y(n6488) );
  AO21X1_LVT U7900 ( .A1(n3856), .A2(div_io_resp_bits_data[49]), .A3(n6488), 
        .Y(n6489) );
  AO21X1_LVT U7901 ( .A1(n3842), .A2(csr_io_rw_rdata[49]), .A3(n6489), .Y(
        n_T_427__T_1136_data[49]) );
  AO22X1_LVT U7902 ( .A1(n3830), .A2(n_T_427[1837]), .A3(n_T_427[1712]), .A4(
        n3824), .Y(n6493) );
  AO22X1_LVT U7903 ( .A1(n3893), .A2(n_T_427[1584]), .A3(n_T_427[1648]), .A4(
        n3887), .Y(n6492) );
  AO22X1_LVT U7904 ( .A1(n3925), .A2(n_T_427[1520]), .A3(n_T_427[1392]), .A4(
        n3919), .Y(n6491) );
  AO22X1_LVT U7905 ( .A1(n3935), .A2(n_T_427[1456]), .A3(n_T_427[1328]), .A4(
        n3930), .Y(n6490) );
  NOR4X1_LVT U7906 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .Y(n6507)
         );
  AO22X1_LVT U7907 ( .A1(n2857), .A2(n_T_427[369]), .A3(n_T_427[561]), .A4(
        n2850), .Y(n6495) );
  AO22X1_LVT U7908 ( .A1(n3822), .A2(n_T_427[880]), .A3(n_T_427[305]), .A4(
        n2828), .Y(n6494) );
  NAND2X0_LVT U7909 ( .A1(n4454), .A2(n3959), .Y(n6503) );
  AO22X1_LVT U7910 ( .A1(n_T_427[689]), .A2(n3861), .A3(n3796), .A4(
        n_T_427[625]), .Y(n6499) );
  AO22X1_LVT U7911 ( .A1(n_T_427[944]), .A2(n6794), .A3(n3812), .A4(
        n_T_427[816]), .Y(n6498) );
  AO22X1_LVT U7912 ( .A1(n6867), .A2(n_T_427[433]), .A3(n3860), .A4(
        n_T_427[241]), .Y(n6497) );
  AO22X1_LVT U7913 ( .A1(n3816), .A2(n_T_427[177]), .A3(n3839), .A4(
        n_T_427[49]), .Y(n6496) );
  NOR4X1_LVT U7914 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .Y(n6500)
         );
  OA22X1_LVT U7915 ( .A1(n3154), .A2(n3803), .A3(n3506), .A4(n3800), .Y(n6501)
         );
  AND3X1_LVT U7916 ( .A1(n6503), .A2(n6502), .A3(n6501), .Y(n6504) );
  NAND4X0_LVT U7917 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .Y(
        id_rs_1[49]) );
  NAND2X0_LVT U7918 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[49]), .Y(n6511) );
  NAND2X0_LVT U7919 ( .A1(n6899), .A2(n_T_918[49]), .Y(n6510) );
  NAND2X0_LVT U7920 ( .A1(n6900), .A2(n_T_1165[49]), .Y(n6509) );
  NAND2X0_LVT U7921 ( .A1(n6901), .A2(n_T_635[49]), .Y(n6508) );
  NAND4X0_LVT U7922 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .Y(
        n_T_702[49]) );
  NAND2X0_LVT U7923 ( .A1(csr_io_rw_rdata[50]), .A2(n3845), .Y(n6514) );
  AOI22X1_LVT U7924 ( .A1(n3853), .A2(io_dmem_resp_bits_data[50]), .A3(n3847), 
        .A4(n_T_1165[50]), .Y(n6513) );
  NAND2X0_LVT U7925 ( .A1(div_io_resp_bits_data[50]), .A2(n3857), .Y(n6512) );
  NAND3X0_LVT U7926 ( .A1(n6514), .A2(n6513), .A3(n6512), .Y(
        n_T_427__T_1136_data[50]) );
  AO22X1_LVT U7927 ( .A1(n3945), .A2(n_T_427[1201]), .A3(n_T_427[1265]), .A4(
        n3940), .Y(n6518) );
  AO22X1_LVT U7928 ( .A1(n3955), .A2(n_T_427[1137]), .A3(n_T_427[1009]), .A4(
        n3950), .Y(n6517) );
  AO22X1_LVT U7929 ( .A1(n3901), .A2(n_T_427[1073]), .A3(n_T_427[242]), .A4(
        n2830), .Y(n6516) );
  AO22X1_LVT U7930 ( .A1(n2864), .A2(n_T_427[434]), .A3(n_T_427[114]), .A4(
        n3831), .Y(n6515) );
  NOR4X1_LVT U7931 ( .A1(n6518), .A2(n6517), .A3(n6516), .A4(n6515), .Y(n6531)
         );
  AO22X1_LVT U7932 ( .A1(n3906), .A2(n_T_427[817]), .A3(n_T_427[753]), .A4(
        n3905), .Y(n6520) );
  AO22X1_LVT U7933 ( .A1(n2856), .A2(n_T_427[370]), .A3(n_T_427[306]), .A4(
        n2828), .Y(n6519) );
  NOR2X0_LVT U7934 ( .A1(n6520), .A2(n6519), .Y(n6530) );
  NAND2X0_LVT U7935 ( .A1(n3958), .A2(n4457), .Y(n6528) );
  AO22X1_LVT U7936 ( .A1(n_T_427[690]), .A2(n3861), .A3(n3868), .A4(
        n_T_427[562]), .Y(n6524) );
  AO22X1_LVT U7937 ( .A1(n_T_427[945]), .A2(n6794), .A3(n3875), .A4(
        n_T_427[881]), .Y(n6523) );
  AO22X1_LVT U7938 ( .A1(n3797), .A2(n_T_427[626]), .A3(n_T_427[498]), .A4(
        n3836), .Y(n6522) );
  AO22X1_LVT U7939 ( .A1(n3816), .A2(n_T_427[178]), .A3(n3840), .A4(
        n_T_427[50]), .Y(n6521) );
  NOR4X1_LVT U7940 ( .A1(n6524), .A2(n6523), .A3(n6522), .A4(n6521), .Y(n6525)
         );
  OA22X1_LVT U7941 ( .A1(n3155), .A2(n2027), .A3(n3507), .A4(n3800), .Y(n6526)
         );
  AND3X1_LVT U7942 ( .A1(n6528), .A2(n6527), .A3(n6526), .Y(n6529) );
  NAND4X0_LVT U7943 ( .A1(n6531), .A2(n6532), .A3(n6530), .A4(n6529), .Y(
        id_rs_1[50]) );
  NAND2X0_LVT U7944 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[50]), .Y(n6536) );
  NAND2X0_LVT U7945 ( .A1(n6899), .A2(n_T_918[50]), .Y(n6535) );
  NAND2X0_LVT U7946 ( .A1(n6900), .A2(n_T_1165[50]), .Y(n6534) );
  NAND2X0_LVT U7947 ( .A1(n3243), .A2(n_T_635[50]), .Y(n6533) );
  NAND4X0_LVT U7948 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .Y(
        n_T_702[50]) );
  AO22X1_LVT U7949 ( .A1(n6860), .A2(io_dmem_resp_bits_data[51]), .A3(n3848), 
        .A4(n_T_1165[51]), .Y(n6537) );
  AO21X1_LVT U7950 ( .A1(n3857), .A2(div_io_resp_bits_data[51]), .A3(n6537), 
        .Y(n6538) );
  AO21X1_LVT U7951 ( .A1(n3841), .A2(csr_io_rw_rdata[51]), .A3(n6538), .Y(
        n_T_427__T_1136_data[51]) );
  AO22X1_LVT U7952 ( .A1(n3828), .A2(n_T_427[1839]), .A3(n_T_427[1714]), .A4(
        n3824), .Y(n6542) );
  AO22X1_LVT U7953 ( .A1(n3893), .A2(n_T_427[1586]), .A3(n_T_427[1650]), .A4(
        n3888), .Y(n6541) );
  AO22X1_LVT U7954 ( .A1(n3925), .A2(n_T_427[1522]), .A3(n_T_427[1394]), .A4(
        n3920), .Y(n6540) );
  AO22X1_LVT U7955 ( .A1(n3935), .A2(n_T_427[1458]), .A3(n_T_427[1330]), .A4(
        n3930), .Y(n6539) );
  NOR4X1_LVT U7956 ( .A1(n6542), .A2(n6541), .A3(n6540), .A4(n6539), .Y(n6556)
         );
  AO22X1_LVT U7957 ( .A1(n2851), .A2(n_T_427[563]), .A3(n_T_427[51]), .A4(
        n2879), .Y(n6544) );
  AO22X1_LVT U7958 ( .A1(n3822), .A2(n_T_427[882]), .A3(n_T_427[691]), .A4(
        n3821), .Y(n6543) );
  NOR2X0_LVT U7959 ( .A1(n6544), .A2(n6543), .Y(n6554) );
  AO22X1_LVT U7960 ( .A1(n3815), .A2(n_T_427[179]), .A3(n_T_427[818]), .A4(
        n3812), .Y(n6548) );
  AO22X1_LVT U7961 ( .A1(n6867), .A2(n_T_427[435]), .A3(n6866), .A4(
        n_T_427[115]), .Y(n6547) );
  AO22X1_LVT U7962 ( .A1(n_T_427[627]), .A2(n3797), .A3(n3867), .A4(
        n_T_427[371]), .Y(n6546) );
  AO22X1_LVT U7963 ( .A1(n3838), .A2(n_T_427[499]), .A3(n3873), .A4(
        n_T_427[307]), .Y(n6545) );
  NOR4X1_LVT U7964 ( .A1(n6548), .A2(n6547), .A3(n6546), .A4(n6545), .Y(n6549)
         );
  OA22X1_LVT U7965 ( .A1(n3156), .A2(n3080), .A3(n3508), .A4(n3800), .Y(n6551)
         );
  NAND2X0_LVT U7966 ( .A1(n4460), .A2(n6898), .Y(n6550) );
  AND3X1_LVT U7967 ( .A1(n6552), .A2(n6551), .A3(n6550), .Y(n6553) );
  NAND4X0_LVT U7968 ( .A1(n6556), .A2(n6555), .A3(n6554), .A4(n6553), .Y(
        id_rs_1[51]) );
  NAND2X0_LVT U7969 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[51]), .Y(n6560) );
  NAND2X0_LVT U7970 ( .A1(n6899), .A2(n_T_918[51]), .Y(n6559) );
  NAND2X0_LVT U7971 ( .A1(n6900), .A2(n_T_1165[51]), .Y(n6558) );
  NAND2X0_LVT U7972 ( .A1(n6901), .A2(n_T_635[51]), .Y(n6557) );
  NAND4X0_LVT U7973 ( .A1(n6560), .A2(n6559), .A3(n6558), .A4(n6557), .Y(
        n_T_702[51]) );
  AO22X1_LVT U7974 ( .A1(n6860), .A2(io_dmem_resp_bits_data[52]), .A3(n3848), 
        .A4(n_T_1165[52]), .Y(n6561) );
  AO21X1_LVT U7975 ( .A1(n3856), .A2(div_io_resp_bits_data[52]), .A3(n6561), 
        .Y(n6562) );
  AO21X1_LVT U7976 ( .A1(n3841), .A2(csr_io_rw_rdata[52]), .A3(n6562), .Y(
        n_T_427__T_1136_data[52]) );
  AO22X1_LVT U7977 ( .A1(n3829), .A2(n_T_427[1840]), .A3(n_T_427[1715]), .A4(
        n3824), .Y(n6566) );
  AO22X1_LVT U7978 ( .A1(n3893), .A2(n_T_427[1587]), .A3(n_T_427[1651]), .A4(
        n3888), .Y(n6565) );
  AO22X1_LVT U7979 ( .A1(n3925), .A2(n_T_427[1523]), .A3(n_T_427[1395]), .A4(
        n3920), .Y(n6564) );
  AO22X1_LVT U7980 ( .A1(n3935), .A2(n_T_427[1459]), .A3(n_T_427[1331]), .A4(
        n3930), .Y(n6563) );
  NOR4X1_LVT U7981 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .Y(n6584)
         );
  AO22X1_LVT U7982 ( .A1(n3945), .A2(n_T_427[1203]), .A3(n_T_427[1267]), .A4(
        n3940), .Y(n6570) );
  AO22X1_LVT U7983 ( .A1(n3955), .A2(n_T_427[1139]), .A3(n_T_427[1011]), .A4(
        n3950), .Y(n6569) );
  AO22X1_LVT U7984 ( .A1(n3902), .A2(n_T_427[1075]), .A3(n_T_427[244]), .A4(
        n3806), .Y(n6568) );
  AO22X1_LVT U7985 ( .A1(n2871), .A2(n_T_427[116]), .A3(n_T_427[947]), .A4(
        n3895), .Y(n6567) );
  NOR4X1_LVT U7986 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .Y(n6583)
         );
  AO22X1_LVT U7987 ( .A1(n2860), .A2(n_T_427[819]), .A3(n_T_427[755]), .A4(
        n3904), .Y(n6572) );
  AO22X1_LVT U7988 ( .A1(n2879), .A2(n_T_427[52]), .A3(n_T_427[692]), .A4(
        n3820), .Y(n6571) );
  NOR2X0_LVT U7989 ( .A1(n6572), .A2(n6571), .Y(n6582) );
  AO22X1_LVT U7990 ( .A1(n3816), .A2(n_T_427[180]), .A3(n_T_427[883]), .A4(
        n3874), .Y(n6576) );
  AO22X1_LVT U7991 ( .A1(n3870), .A2(n_T_427[564]), .A3(n_T_427[628]), .A4(
        n3795), .Y(n6575) );
  AO22X1_LVT U7992 ( .A1(n6867), .A2(n_T_427[436]), .A3(n3867), .A4(
        n_T_427[372]), .Y(n6574) );
  AO22X1_LVT U7993 ( .A1(n3838), .A2(n_T_427[500]), .A3(n3873), .A4(
        n_T_427[308]), .Y(n6573) );
  NOR4X1_LVT U7994 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .Y(n6577)
         );
  OA22X1_LVT U7995 ( .A1(n3157), .A2(n1994), .A3(n3509), .A4(n3800), .Y(n6579)
         );
  NAND2X0_LVT U7996 ( .A1(n4463), .A2(n6898), .Y(n6578) );
  AND3X1_LVT U7997 ( .A1(n6580), .A2(n6579), .A3(n6578), .Y(n6581) );
  NAND4X0_LVT U7998 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .Y(
        id_rs_1[52]) );
  NAND2X0_LVT U7999 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[52]), .Y(n6588) );
  NAND2X0_LVT U8000 ( .A1(n6899), .A2(n_T_918[52]), .Y(n6587) );
  NAND2X0_LVT U8001 ( .A1(n6900), .A2(n_T_1165[52]), .Y(n6586) );
  NAND2X0_LVT U8002 ( .A1(n6901), .A2(n_T_635[52]), .Y(n6585) );
  NAND4X0_LVT U8003 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .Y(
        n_T_702[52]) );
  NAND2X0_LVT U8004 ( .A1(csr_io_rw_rdata[53]), .A2(n3845), .Y(n6591) );
  AOI22X1_LVT U8005 ( .A1(n3853), .A2(io_dmem_resp_bits_data[53]), .A3(n3847), 
        .A4(n_T_1165[53]), .Y(n6590) );
  NAND2X0_LVT U8006 ( .A1(div_io_resp_bits_data[53]), .A2(n3857), .Y(n6589) );
  NAND3X0_LVT U8007 ( .A1(n6591), .A2(n6590), .A3(n6589), .Y(
        n_T_427__T_1136_data[53]) );
  AO22X1_LVT U8008 ( .A1(n3946), .A2(n_T_427[1204]), .A3(n_T_427[1268]), .A4(
        n3940), .Y(n6595) );
  AO22X1_LVT U8009 ( .A1(n3956), .A2(n_T_427[1140]), .A3(n_T_427[1012]), .A4(
        n3950), .Y(n6594) );
  AO22X1_LVT U8010 ( .A1(n3902), .A2(n_T_427[1076]), .A3(n_T_427[245]), .A4(
        n3808), .Y(n6593) );
  AO22X1_LVT U8011 ( .A1(n2832), .A2(n_T_427[948]), .A3(n_T_427[756]), .A4(
        n2827), .Y(n6592) );
  NOR4X1_LVT U8012 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .Y(n6608)
         );
  AO22X1_LVT U8013 ( .A1(n3906), .A2(n_T_427[820]), .A3(n_T_427[373]), .A4(
        n1918), .Y(n6597) );
  AO22X1_LVT U8014 ( .A1(n2850), .A2(n_T_427[565]), .A3(n_T_427[693]), .A4(
        n3820), .Y(n6596) );
  NOR2X0_LVT U8015 ( .A1(n6597), .A2(n6596), .Y(n6607) );
  AO22X1_LVT U8016 ( .A1(n3797), .A2(n_T_427[629]), .A3(n_T_427[501]), .A4(
        n3836), .Y(n6601) );
  AO22X1_LVT U8017 ( .A1(n6867), .A2(n_T_427[437]), .A3(n3864), .A4(
        n_T_427[117]), .Y(n6600) );
  AO22X1_LVT U8018 ( .A1(n_T_427[884]), .A2(n6871), .A3(n3873), .A4(
        n_T_427[309]), .Y(n6599) );
  AO22X1_LVT U8019 ( .A1(n3816), .A2(n_T_427[181]), .A3(n3840), .A4(
        n_T_427[53]), .Y(n6598) );
  NOR4X1_LVT U8020 ( .A1(n6601), .A2(n6600), .A3(n6599), .A4(n6598), .Y(n6602)
         );
  OA22X1_LVT U8021 ( .A1(n3561), .A2(n3882), .A3(n1993), .A4(n6602), .Y(n6605)
         );
  NAND2X0_LVT U8022 ( .A1(n3958), .A2(n4466), .Y(n6604) );
  OA22X1_LVT U8023 ( .A1(n3158), .A2(n2027), .A3(n3510), .A4(n3800), .Y(n6603)
         );
  AND3X1_LVT U8024 ( .A1(n6605), .A2(n6604), .A3(n6603), .Y(n6606) );
  NAND4X0_LVT U8025 ( .A1(n6608), .A2(n6609), .A3(n6607), .A4(n6606), .Y(
        id_rs_1[53]) );
  NAND2X0_LVT U8026 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[53]), .Y(n6613) );
  NAND2X0_LVT U8027 ( .A1(n6899), .A2(n_T_918[53]), .Y(n6612) );
  NAND2X0_LVT U8028 ( .A1(n6900), .A2(n_T_1165[53]), .Y(n6611) );
  NAND2X0_LVT U8029 ( .A1(n6901), .A2(n_T_635[53]), .Y(n6610) );
  NAND4X0_LVT U8030 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .Y(
        n_T_702[53]) );
  AO22X1_LVT U8031 ( .A1(n6860), .A2(io_dmem_resp_bits_data[54]), .A3(n3848), 
        .A4(n_T_1165[54]), .Y(n6614) );
  AO21X1_LVT U8032 ( .A1(n3856), .A2(div_io_resp_bits_data[54]), .A3(n6614), 
        .Y(n6615) );
  AO21X1_LVT U8033 ( .A1(n3841), .A2(csr_io_rw_rdata[54]), .A3(n6615), .Y(
        n_T_427__T_1136_data[54]) );
  AO22X1_LVT U8034 ( .A1(n2856), .A2(n_T_427[374]), .A3(n_T_427[182]), .A4(
        n3908), .Y(n6617) );
  AO22X1_LVT U8035 ( .A1(n3809), .A2(n_T_427[310]), .A3(n_T_427[694]), .A4(
        n2829), .Y(n6616) );
  NOR2X0_LVT U8036 ( .A1(n6617), .A2(n6616), .Y(n6627) );
  AO22X1_LVT U8037 ( .A1(n3870), .A2(n_T_427[566]), .A3(n3860), .A4(
        n_T_427[246]), .Y(n6621) );
  AO22X1_LVT U8038 ( .A1(n_T_427[757]), .A2(n3804), .A3(n6866), .A4(
        n_T_427[118]), .Y(n6620) );
  AO22X1_LVT U8039 ( .A1(n3797), .A2(n_T_427[630]), .A3(n_T_427[502]), .A4(
        n3836), .Y(n6619) );
  AO22X1_LVT U8040 ( .A1(n_T_427[885]), .A2(n6871), .A3(n3840), .A4(
        n_T_427[54]), .Y(n6618) );
  NOR4X1_LVT U8041 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .Y(n6622)
         );
  OA22X1_LVT U8042 ( .A1(n3159), .A2(n3080), .A3(n3511), .A4(n3800), .Y(n6624)
         );
  NAND2X0_LVT U8043 ( .A1(n4469), .A2(n6898), .Y(n6623) );
  AND3X1_LVT U8044 ( .A1(n6625), .A2(n6624), .A3(n6623), .Y(n6626) );
  NAND4X0_LVT U8045 ( .A1(n6628), .A2(n6629), .A3(n6627), .A4(n6626), .Y(
        id_rs_1[54]) );
  NAND2X0_LVT U8046 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[54]), .Y(n6633) );
  NAND2X0_LVT U8047 ( .A1(n6899), .A2(n_T_918[54]), .Y(n6632) );
  NAND2X0_LVT U8048 ( .A1(n6900), .A2(n_T_1165[54]), .Y(n6631) );
  NAND2X0_LVT U8049 ( .A1(n3243), .A2(n_T_635[54]), .Y(n6630) );
  NAND4X0_LVT U8050 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .Y(
        n_T_702[54]) );
  NAND2X0_LVT U8051 ( .A1(csr_io_rw_rdata[55]), .A2(n3845), .Y(n6636) );
  AOI22X1_LVT U8052 ( .A1(n3853), .A2(io_dmem_resp_bits_data[55]), .A3(n3847), 
        .A4(n_T_1165[55]), .Y(n6635) );
  NAND2X0_LVT U8053 ( .A1(div_io_resp_bits_data[55]), .A2(n3857), .Y(n6634) );
  NAND3X0_LVT U8054 ( .A1(n6636), .A2(n6635), .A3(n6634), .Y(
        n_T_427__T_1136_data[55]) );
  AO22X1_LVT U8055 ( .A1(n_T_427[695]), .A2(n3862), .A3(n3860), .A4(
        n_T_427[247]), .Y(n6640) );
  AO22X1_LVT U8056 ( .A1(n3816), .A2(n_T_427[183]), .A3(n_T_427[886]), .A4(
        n3874), .Y(n6639) );
  AO22X1_LVT U8057 ( .A1(n6867), .A2(n_T_427[439]), .A3(n6866), .A4(
        n_T_427[119]), .Y(n6638) );
  AO22X1_LVT U8058 ( .A1(n3838), .A2(n_T_427[503]), .A3(n3867), .A4(
        n_T_427[375]), .Y(n6637) );
  NOR4X1_LVT U8059 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .Y(n6641)
         );
  OA22X1_LVT U8060 ( .A1(n3563), .A2(n3882), .A3(n3877), .A4(n6641), .Y(n6645)
         );
  OA22X1_LVT U8061 ( .A1(n3160), .A2(n3080), .A3(n3512), .A4(n3800), .Y(n6644)
         );
  AOI22X1_LVT U8062 ( .A1(n3894), .A2(n_T_427[1590]), .A3(n_T_427[1654]), .A4(
        n3889), .Y(n6643) );
  OA22X1_LVT U8063 ( .A1(n3161), .A2(n3081), .A3(n3513), .A4(n3082), .Y(n6642)
         );
  AND4X1_LVT U8064 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .Y(n6657)
         );
  AO22X1_LVT U8065 ( .A1(n3902), .A2(n_T_427[1078]), .A3(n_T_427[950]), .A4(
        n2832), .Y(n6649) );
  AO22X1_LVT U8066 ( .A1(n2861), .A2(n_T_427[822]), .A3(n_T_427[758]), .A4(
        n2827), .Y(n6648) );
  AO22X1_LVT U8067 ( .A1(n2869), .A2(n_T_427[631]), .A3(n_T_427[55]), .A4(
        n2826), .Y(n6647) );
  AO22X1_LVT U8068 ( .A1(n2850), .A2(n_T_427[567]), .A3(n_T_427[311]), .A4(
        n6774), .Y(n6646) );
  NOR4X1_LVT U8069 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .Y(n6656)
         );
  AO22X1_LVT U8070 ( .A1(n3926), .A2(n_T_427[1526]), .A3(n_T_427[1398]), .A4(
        n3919), .Y(n6653) );
  AO22X1_LVT U8071 ( .A1(n3936), .A2(n_T_427[1462]), .A3(n_T_427[1334]), .A4(
        n3930), .Y(n6652) );
  AO22X1_LVT U8072 ( .A1(n3946), .A2(n_T_427[1206]), .A3(n_T_427[1270]), .A4(
        n3939), .Y(n6651) );
  AO22X1_LVT U8073 ( .A1(n3956), .A2(n_T_427[1142]), .A3(n_T_427[1014]), .A4(
        n3949), .Y(n6650) );
  NOR4X1_LVT U8074 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .Y(n6655)
         );
  NAND2X0_LVT U8075 ( .A1(n3957), .A2(n4472), .Y(n6654) );
  NAND4X0_LVT U8076 ( .A1(n6656), .A2(n6657), .A3(n6655), .A4(n6654), .Y(
        id_rs_1[55]) );
  NAND2X0_LVT U8077 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[55]), .Y(n6661) );
  NAND2X0_LVT U8078 ( .A1(n6899), .A2(n_T_918[55]), .Y(n6660) );
  NAND2X0_LVT U8079 ( .A1(n6900), .A2(n_T_1165[55]), .Y(n6659) );
  NAND2X0_LVT U8080 ( .A1(n6901), .A2(n_T_635[55]), .Y(n6658) );
  NAND4X0_LVT U8081 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .Y(
        n_T_702[55]) );
  AO22X1_LVT U8082 ( .A1(n6860), .A2(io_dmem_resp_bits_data[56]), .A3(n3848), 
        .A4(n_T_1165[56]), .Y(n6662) );
  AO21X1_LVT U8083 ( .A1(n3856), .A2(div_io_resp_bits_data[56]), .A3(n6662), 
        .Y(n6663) );
  AO21X1_LVT U8084 ( .A1(n3841), .A2(csr_io_rw_rdata[56]), .A3(n6663), .Y(
        n_T_427__T_1136_data[56]) );
  AO22X1_LVT U8085 ( .A1(n3830), .A2(n_T_427[1843]), .A3(n_T_427[1719]), .A4(
        n3824), .Y(n6667) );
  AO22X1_LVT U8086 ( .A1(n3894), .A2(n_T_427[1591]), .A3(n_T_427[1655]), .A4(
        n3887), .Y(n6666) );
  AO22X1_LVT U8087 ( .A1(n3926), .A2(n_T_427[1527]), .A3(n_T_427[1399]), .A4(
        n3920), .Y(n6665) );
  AO22X1_LVT U8088 ( .A1(n3936), .A2(n_T_427[1463]), .A3(n_T_427[1335]), .A4(
        n3929), .Y(n6664) );
  NOR4X1_LVT U8089 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .Y(n6681)
         );
  AO22X1_LVT U8090 ( .A1(n1919), .A2(n_T_427[376]), .A3(n_T_427[632]), .A4(
        n2870), .Y(n6669) );
  AO22X1_LVT U8091 ( .A1(n3822), .A2(n_T_427[887]), .A3(n_T_427[696]), .A4(
        n2829), .Y(n6668) );
  NOR2X0_LVT U8092 ( .A1(n6669), .A2(n6668), .Y(n6679) );
  AO22X1_LVT U8093 ( .A1(n3870), .A2(n_T_427[568]), .A3(n3860), .A4(
        n_T_427[248]), .Y(n6673) );
  AO22X1_LVT U8094 ( .A1(n_T_427[759]), .A2(n3804), .A3(n6866), .A4(
        n_T_427[120]), .Y(n6672) );
  AO22X1_LVT U8095 ( .A1(n3838), .A2(n_T_427[504]), .A3(n3873), .A4(
        n_T_427[312]), .Y(n6671) );
  AO22X1_LVT U8096 ( .A1(n_T_427[823]), .A2(n3813), .A3(n3840), .A4(
        n_T_427[56]), .Y(n6670) );
  NOR4X1_LVT U8097 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .Y(n6674)
         );
  NAND2X0_LVT U8098 ( .A1(n4475), .A2(n6898), .Y(n6675) );
  AND3X1_LVT U8099 ( .A1(n6677), .A2(n6676), .A3(n6675), .Y(n6678) );
  NAND4X0_LVT U8100 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .Y(
        id_rs_1[56]) );
  NAND2X0_LVT U8101 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[56]), .Y(n6685) );
  NAND2X0_LVT U8102 ( .A1(n6899), .A2(n_T_918[56]), .Y(n6684) );
  NAND2X0_LVT U8103 ( .A1(n6900), .A2(n_T_1165[56]), .Y(n6683) );
  NAND2X0_LVT U8104 ( .A1(n6901), .A2(n_T_635[56]), .Y(n6682) );
  NAND4X0_LVT U8105 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .Y(
        n_T_702[56]) );
  NAND2X0_LVT U8106 ( .A1(csr_io_rw_rdata[57]), .A2(n3845), .Y(n6688) );
  AOI22X1_LVT U8107 ( .A1(n3853), .A2(io_dmem_resp_bits_data[57]), .A3(n3847), 
        .A4(n_T_1165[57]), .Y(n6687) );
  NAND2X0_LVT U8108 ( .A1(div_io_resp_bits_data[57]), .A2(n3857), .Y(n6686) );
  NAND3X0_LVT U8109 ( .A1(n6688), .A2(n6687), .A3(n6686), .Y(
        n_T_427__T_1136_data[57]) );
  AO22X1_LVT U8110 ( .A1(n3907), .A2(n_T_427[824]), .A3(n_T_427[185]), .A4(
        n3908), .Y(n6690) );
  AO22X1_LVT U8111 ( .A1(n2870), .A2(n_T_427[633]), .A3(n_T_427[888]), .A4(
        n3822), .Y(n6689) );
  NOR2X0_LVT U8112 ( .A1(n6690), .A2(n6689), .Y(n6700) );
  AO22X1_LVT U8113 ( .A1(n_T_427[697]), .A2(n3861), .A3(n3865), .A4(
        n_T_427[441]), .Y(n6694) );
  AO22X1_LVT U8114 ( .A1(n_T_427[952]), .A2(n6794), .A3(n3837), .A4(
        n_T_427[505]), .Y(n6693) );
  AO22X1_LVT U8115 ( .A1(n_T_427[569]), .A2(n3869), .A3(n3867), .A4(
        n_T_427[377]), .Y(n6692) );
  AO22X1_LVT U8116 ( .A1(n3871), .A2(n_T_427[313]), .A3(n3840), .A4(
        n_T_427[57]), .Y(n6691) );
  NOR4X1_LVT U8117 ( .A1(n6694), .A2(n6693), .A3(n6692), .A4(n6691), .Y(n6695)
         );
  NAND2X0_LVT U8118 ( .A1(n3958), .A2(n4478), .Y(n6697) );
  OA22X1_LVT U8119 ( .A1(n3163), .A2(n3080), .A3(n3515), .A4(n3800), .Y(n6696)
         );
  AND3X1_LVT U8120 ( .A1(n6698), .A2(n6697), .A3(n6696), .Y(n6699) );
  NAND4X0_LVT U8121 ( .A1(n6701), .A2(n6702), .A3(n6700), .A4(n6699), .Y(
        id_rs_1[57]) );
  NAND2X0_LVT U8122 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[57]), .Y(n6706) );
  NAND2X0_LVT U8123 ( .A1(n6899), .A2(n_T_918[57]), .Y(n6705) );
  NAND2X0_LVT U8124 ( .A1(n6900), .A2(n_T_1165[57]), .Y(n6704) );
  NAND2X0_LVT U8125 ( .A1(n3243), .A2(n_T_635[57]), .Y(n6703) );
  NAND4X0_LVT U8126 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .Y(
        n_T_702[57]) );
  AO22X1_LVT U8127 ( .A1(n6860), .A2(io_dmem_resp_bits_data[58]), .A3(n3849), 
        .A4(n_T_1165[58]), .Y(n6707) );
  AO21X1_LVT U8128 ( .A1(n3856), .A2(div_io_resp_bits_data[58]), .A3(n6707), 
        .Y(n6708) );
  AO21X1_LVT U8129 ( .A1(n3841), .A2(csr_io_rw_rdata[58]), .A3(n6708), .Y(
        n_T_427__T_1136_data[58]) );
  AO22X1_LVT U8130 ( .A1(n3828), .A2(n_T_427[1845]), .A3(n_T_427[1721]), .A4(
        n3824), .Y(n6712) );
  AO22X1_LVT U8131 ( .A1(n3894), .A2(n_T_427[1593]), .A3(n_T_427[1657]), .A4(
        n3888), .Y(n6711) );
  AO22X1_LVT U8132 ( .A1(n3926), .A2(n_T_427[1529]), .A3(n_T_427[1401]), .A4(
        n3921), .Y(n6710) );
  AO22X1_LVT U8133 ( .A1(n3936), .A2(n_T_427[1465]), .A3(n_T_427[1337]), .A4(
        n3931), .Y(n6709) );
  NOR4X1_LVT U8134 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .Y(n6727)
         );
  AO22X1_LVT U8135 ( .A1(n3912), .A2(n_T_427[506]), .A3(n_T_427[889]), .A4(
        n2833), .Y(n6714) );
  AO22X1_LVT U8136 ( .A1(n3810), .A2(n_T_427[314]), .A3(n_T_427[698]), .A4(
        n3820), .Y(n6713) );
  NOR2X0_LVT U8137 ( .A1(n6714), .A2(n6713), .Y(n6725) );
  AO22X1_LVT U8138 ( .A1(n_T_427[953]), .A2(n6794), .A3(n3796), .A4(
        n_T_427[634]), .Y(n6719) );
  AO22X1_LVT U8139 ( .A1(n6867), .A2(n_T_427[442]), .A3(n6866), .A4(
        n_T_427[122]), .Y(n6718) );
  AO22X1_LVT U8140 ( .A1(n_T_427[570]), .A2(n3869), .A3(n3867), .A4(
        n_T_427[378]), .Y(n6717) );
  AO22X1_LVT U8141 ( .A1(n3816), .A2(n_T_427[186]), .A3(n3840), .A4(
        n_T_427[58]), .Y(n6716) );
  NOR4X1_LVT U8142 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .Y(n6720)
         );
  OA22X1_LVT U8143 ( .A1(n3164), .A2(n3080), .A3(n3516), .A4(n3800), .Y(n6722)
         );
  NAND2X0_LVT U8144 ( .A1(n4481), .A2(n3958), .Y(n6721) );
  AND3X1_LVT U8145 ( .A1(n6723), .A2(n6722), .A3(n6721), .Y(n6724) );
  NAND4X0_LVT U8146 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .Y(
        id_rs_1[58]) );
  NAND2X0_LVT U8147 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[58]), .Y(n6731) );
  NAND2X0_LVT U8148 ( .A1(n6899), .A2(n_T_918[58]), .Y(n6730) );
  NAND2X0_LVT U8149 ( .A1(n6900), .A2(n_T_1165[58]), .Y(n6729) );
  NAND2X0_LVT U8150 ( .A1(n3243), .A2(n_T_635[58]), .Y(n6728) );
  NAND4X0_LVT U8151 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .Y(
        n_T_702[58]) );
  NAND2X0_LVT U8152 ( .A1(csr_io_rw_rdata[59]), .A2(n3845), .Y(n6734) );
  AOI22X1_LVT U8153 ( .A1(n3853), .A2(io_dmem_resp_bits_data[59]), .A3(n3847), 
        .A4(n_T_1165[59]), .Y(n6733) );
  NAND2X0_LVT U8154 ( .A1(div_io_resp_bits_data[59]), .A2(n3857), .Y(n6732) );
  NAND3X0_LVT U8155 ( .A1(n6734), .A2(n6733), .A3(n6732), .Y(
        n_T_427__T_1136_data[59]) );
  AO22X1_LVT U8156 ( .A1(n3814), .A2(n_T_427[826]), .A3(n_T_427[890]), .A4(
        n3874), .Y(n6738) );
  AO22X1_LVT U8157 ( .A1(n_T_427[699]), .A2(n3861), .A3(n6866), .A4(
        n_T_427[123]), .Y(n6737) );
  AO22X1_LVT U8158 ( .A1(n3838), .A2(n_T_427[507]), .A3(n3867), .A4(
        n_T_427[379]), .Y(n6736) );
  AO22X1_LVT U8159 ( .A1(n3816), .A2(n_T_427[187]), .A3(n3840), .A4(
        n_T_427[59]), .Y(n6735) );
  NOR4X1_LVT U8160 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .Y(n6739)
         );
  OA22X1_LVT U8161 ( .A1(n3165), .A2(n2027), .A3(n3517), .A4(n3800), .Y(n6742)
         );
  OA22X1_LVT U8162 ( .A1(n3166), .A2(n3081), .A3(n3518), .A4(n3082), .Y(n6741)
         );
  AOI22X1_LVT U8163 ( .A1(n3894), .A2(n_T_427[1594]), .A3(n_T_427[1658]), .A4(
        n3889), .Y(n6740) );
  AND4X1_LVT U8164 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .Y(n6755)
         );
  AO22X1_LVT U8165 ( .A1(n3902), .A2(n_T_427[1082]), .A3(n_T_427[251]), .A4(
        n3808), .Y(n6747) );
  AO22X1_LVT U8166 ( .A1(n2864), .A2(n_T_427[443]), .A3(n_T_427[954]), .A4(
        n3897), .Y(n6746) );
  AO22X1_LVT U8167 ( .A1(n3915), .A2(n_T_427[635]), .A3(n_T_427[762]), .A4(
        n2827), .Y(n6745) );
  AO22X1_LVT U8168 ( .A1(n2851), .A2(n_T_427[571]), .A3(n_T_427[315]), .A4(
        n2828), .Y(n6744) );
  NOR4X1_LVT U8169 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .Y(n6754)
         );
  AO22X1_LVT U8170 ( .A1(n3926), .A2(n_T_427[1530]), .A3(n_T_427[1402]), .A4(
        n3920), .Y(n6751) );
  AO22X1_LVT U8171 ( .A1(n3936), .A2(n_T_427[1466]), .A3(n_T_427[1338]), .A4(
        n3931), .Y(n6750) );
  AO22X1_LVT U8172 ( .A1(n3946), .A2(n_T_427[1210]), .A3(n_T_427[1274]), .A4(
        n3940), .Y(n6749) );
  AO22X1_LVT U8173 ( .A1(n3956), .A2(n_T_427[1146]), .A3(n_T_427[1018]), .A4(
        n3950), .Y(n6748) );
  NOR4X1_LVT U8174 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .Y(n6753)
         );
  NAND2X0_LVT U8175 ( .A1(n3957), .A2(n4484), .Y(n6752) );
  NAND4X0_LVT U8176 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .Y(
        id_rs_1[59]) );
  NAND2X0_LVT U8177 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[59]), .Y(n6759) );
  NAND2X0_LVT U8178 ( .A1(n6899), .A2(n_T_918[59]), .Y(n6758) );
  NAND2X0_LVT U8179 ( .A1(n6900), .A2(n_T_1165[59]), .Y(n6757) );
  NAND2X0_LVT U8180 ( .A1(n6901), .A2(n_T_635[59]), .Y(n6756) );
  NAND4X0_LVT U8181 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .Y(
        n_T_702[59]) );
  NAND2X0_LVT U8182 ( .A1(csr_io_rw_rdata[60]), .A2(n3845), .Y(n6762) );
  AOI22X1_LVT U8183 ( .A1(n3853), .A2(io_dmem_resp_bits_data[60]), .A3(n3847), 
        .A4(n_T_1165[60]), .Y(n6761) );
  NAND2X0_LVT U8184 ( .A1(div_io_resp_bits_data[60]), .A2(n3857), .Y(n6760) );
  NAND3X0_LVT U8185 ( .A1(n6762), .A2(n6761), .A3(n6760), .Y(
        n_T_427__T_1136_data[60]) );
  AOI22X1_LVT U8186 ( .A1(n6765), .A2(n_T_427[763]), .A3(n3864), .A4(
        n_T_427[124]), .Y(n6771) );
  AOI22X1_LVT U8187 ( .A1(n3814), .A2(n_T_427[827]), .A3(n6838), .A4(
        n_T_427[60]), .Y(n6770) );
  AOI22X1_LVT U8188 ( .A1(n3838), .A2(n_T_427[508]), .A3(n_T_427[572]), .A4(
        n3868), .Y(n6769) );
  OA22X1_LVT U8189 ( .A1(n6767), .A2(n3525), .A3(n3172), .A4(n6766), .Y(n6768)
         );
  NAND4X0_LVT U8190 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .Y(n6772) );
  AO22X1_LVT U8191 ( .A1(n3902), .A2(n_T_427[1083]), .A3(n_T_427[252]), .A4(
        n3807), .Y(n6778) );
  AO22X1_LVT U8192 ( .A1(n3915), .A2(n_T_427[636]), .A3(n_T_427[891]), .A4(
        n6813), .Y(n6777) );
  AO22X1_LVT U8193 ( .A1(n2831), .A2(n_T_427[955]), .A3(n_T_427[188]), .A4(
        n2862), .Y(n6776) );
  AO22X1_LVT U8194 ( .A1(n3810), .A2(n_T_427[316]), .A3(n_T_427[700]), .A4(
        n3821), .Y(n6775) );
  NOR4X1_LVT U8195 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .Y(n6785)
         );
  AO22X1_LVT U8196 ( .A1(n3926), .A2(n_T_427[1531]), .A3(n_T_427[1403]), .A4(
        n3921), .Y(n6782) );
  AO22X1_LVT U8197 ( .A1(n3936), .A2(n_T_427[1467]), .A3(n_T_427[1339]), .A4(
        n3931), .Y(n6781) );
  AO22X1_LVT U8198 ( .A1(n3946), .A2(n_T_427[1211]), .A3(n_T_427[1275]), .A4(
        n3941), .Y(n6780) );
  AO22X1_LVT U8199 ( .A1(n3956), .A2(n_T_427[1147]), .A3(n_T_427[1019]), .A4(
        n3951), .Y(n6779) );
  NOR4X1_LVT U8200 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .Y(n6784)
         );
  NAND2X0_LVT U8201 ( .A1(n3957), .A2(n4487), .Y(n6783) );
  NAND4X0_LVT U8202 ( .A1(n6785), .A2(n6786), .A3(n6784), .A4(n6783), .Y(
        id_rs_1[60]) );
  NAND2X0_LVT U8203 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[60]), .Y(n6790) );
  NAND2X0_LVT U8204 ( .A1(n6899), .A2(n_T_918[60]), .Y(n6789) );
  NAND2X0_LVT U8205 ( .A1(n6900), .A2(n_T_1165[60]), .Y(n6788) );
  NAND2X0_LVT U8206 ( .A1(n6901), .A2(n_T_635[60]), .Y(n6787) );
  NAND4X0_LVT U8207 ( .A1(n6790), .A2(n6789), .A3(n6788), .A4(n6787), .Y(
        n_T_702[60]) );
  NAND2X0_LVT U8208 ( .A1(csr_io_rw_rdata[61]), .A2(n3842), .Y(n6793) );
  AOI22X1_LVT U8209 ( .A1(n3853), .A2(io_dmem_resp_bits_data[61]), .A3(n3847), 
        .A4(n_T_1165[61]), .Y(n6792) );
  NAND2X0_LVT U8210 ( .A1(div_io_resp_bits_data[61]), .A2(n3857), .Y(n6791) );
  NAND3X0_LVT U8211 ( .A1(n6793), .A2(n6792), .A3(n6791), .Y(
        n_T_427__T_1136_data[61]) );
  AO22X1_LVT U8212 ( .A1(n_T_427[956]), .A2(n3811), .A3(n3837), .A4(
        n_T_427[509]), .Y(n6800) );
  AO22X1_LVT U8213 ( .A1(n_T_427[828]), .A2(n3813), .A3(n3873), .A4(
        n_T_427[317]), .Y(n6799) );
  AO22X1_LVT U8214 ( .A1(n3816), .A2(n_T_427[189]), .A3(n3840), .A4(
        n_T_427[61]), .Y(n6798) );
  AO22X1_LVT U8215 ( .A1(n3860), .A2(n_T_427[253]), .A3(n6866), .A4(
        n_T_427[125]), .Y(n6797) );
  NOR4X1_LVT U8216 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .Y(n6801)
         );
  OA22X1_LVT U8217 ( .A1(n3167), .A2(n1994), .A3(n3485), .A4(n3800), .Y(n6804)
         );
  OA22X1_LVT U8218 ( .A1(n3168), .A2(n3081), .A3(n3486), .A4(n3082), .Y(n6803)
         );
  AOI22X1_LVT U8219 ( .A1(n3894), .A2(n_T_427[1596]), .A3(n_T_427[1660]), .A4(
        n3889), .Y(n6802) );
  AND4X1_LVT U8220 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .Y(n6821)
         );
  AO22X1_LVT U8221 ( .A1(n3926), .A2(n_T_427[1532]), .A3(n_T_427[1404]), .A4(
        n3921), .Y(n6809) );
  AO22X1_LVT U8222 ( .A1(n3936), .A2(n_T_427[1468]), .A3(n_T_427[1340]), .A4(
        n3931), .Y(n6808) );
  AO22X1_LVT U8223 ( .A1(n3946), .A2(n_T_427[1212]), .A3(n_T_427[1276]), .A4(
        n3941), .Y(n6807) );
  AO22X1_LVT U8224 ( .A1(n3956), .A2(n_T_427[1148]), .A3(n_T_427[1020]), .A4(
        n3951), .Y(n6806) );
  NOR4X1_LVT U8225 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .Y(n6820)
         );
  AO22X1_LVT U8226 ( .A1(n3834), .A2(n_T_427[445]), .A3(n_T_427[1084]), .A4(
        n3898), .Y(n6817) );
  AO22X1_LVT U8227 ( .A1(n1918), .A2(n_T_427[381]), .A3(n_T_427[764]), .A4(
        n3903), .Y(n6816) );
  AO22X1_LVT U8228 ( .A1(n3818), .A2(n_T_427[573]), .A3(n_T_427[637]), .A4(
        n2869), .Y(n6815) );
  AO22X1_LVT U8229 ( .A1(n3823), .A2(n_T_427[892]), .A3(n_T_427[701]), .A4(
        n3821), .Y(n6814) );
  NOR4X1_LVT U8230 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(n6814), .Y(n6819)
         );
  NAND2X0_LVT U8231 ( .A1(n3958), .A2(n4490), .Y(n6818) );
  NAND4X0_LVT U8232 ( .A1(n6820), .A2(n6821), .A3(n6819), .A4(n6818), .Y(
        id_rs_1[61]) );
  NAND2X0_LVT U8233 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[61]), .Y(n6825) );
  NAND2X0_LVT U8234 ( .A1(n6899), .A2(n_T_918[61]), .Y(n6824) );
  NAND2X0_LVT U8235 ( .A1(n6900), .A2(n_T_1165[61]), .Y(n6823) );
  NAND2X0_LVT U8236 ( .A1(n3243), .A2(n_T_635[61]), .Y(n6822) );
  NAND4X0_LVT U8237 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .Y(
        n_T_702[61]) );
  NAND2X0_LVT U8238 ( .A1(csr_io_rw_rdata[62]), .A2(n3844), .Y(n6828) );
  AOI22X1_LVT U8239 ( .A1(n3852), .A2(io_dmem_resp_bits_data[62]), .A3(n3847), 
        .A4(n_T_1165[62]), .Y(n6827) );
  NAND2X0_LVT U8240 ( .A1(div_io_resp_bits_data[62]), .A2(n3857), .Y(n6826) );
  NAND3X0_LVT U8241 ( .A1(n6828), .A2(n6827), .A3(n6826), .Y(
        n_T_427__T_1136_data[62]) );
  AO22X1_LVT U8242 ( .A1(n3946), .A2(n_T_427[1213]), .A3(n_T_427[1277]), .A4(
        n3940), .Y(n6834) );
  AO22X1_LVT U8243 ( .A1(n3956), .A2(n_T_427[1149]), .A3(n_T_427[1021]), .A4(
        n3950), .Y(n6833) );
  AO22X1_LVT U8244 ( .A1(n3902), .A2(n_T_427[1085]), .A3(n_T_427[957]), .A4(
        n2832), .Y(n6832) );
  AO22X1_LVT U8245 ( .A1(n2864), .A2(n_T_427[446]), .A3(n_T_427[126]), .A4(
        n2872), .Y(n6831) );
  NOR4X1_LVT U8246 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .Y(n6849)
         );
  AO22X1_LVT U8247 ( .A1(n2860), .A2(n_T_427[829]), .A3(n_T_427[765]), .A4(
        n2827), .Y(n6836) );
  AO22X1_LVT U8248 ( .A1(n2869), .A2(n_T_427[638]), .A3(n_T_427[190]), .A4(
        n2863), .Y(n6835) );
  NOR2X0_LVT U8249 ( .A1(n6836), .A2(n6835), .Y(n6848) );
  AO22X1_LVT U8250 ( .A1(n_T_427[702]), .A2(n3861), .A3(n3860), .A4(
        n_T_427[254]), .Y(n6842) );
  AO22X1_LVT U8251 ( .A1(n_T_427[574]), .A2(n3868), .A3(n6868), .A4(
        n_T_427[382]), .Y(n6841) );
  AO22X1_LVT U8252 ( .A1(n3837), .A2(n_T_427[510]), .A3(n3873), .A4(
        n_T_427[318]), .Y(n6840) );
  AO22X1_LVT U8253 ( .A1(n_T_427[893]), .A2(n6871), .A3(n6838), .A4(
        n_T_427[62]), .Y(n6839) );
  NOR4X1_LVT U8254 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .Y(n6843)
         );
  NAND2X0_LVT U8255 ( .A1(n3957), .A2(n4493), .Y(n6845) );
  OA22X1_LVT U8256 ( .A1(n3169), .A2(n2027), .A3(n3487), .A4(n3800), .Y(n6844)
         );
  AND3X1_LVT U8257 ( .A1(n6846), .A2(n6845), .A3(n6844), .Y(n6847) );
  NAND4X0_LVT U8258 ( .A1(n6849), .A2(n6850), .A3(n6848), .A4(n6847), .Y(
        id_rs_1[62]) );
  NAND2X0_LVT U8259 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[62]), .Y(n6854) );
  NAND2X0_LVT U8260 ( .A1(n6899), .A2(n_T_918[62]), .Y(n6853) );
  NAND2X0_LVT U8261 ( .A1(n6900), .A2(n_T_1165[62]), .Y(n6852) );
  NAND2X0_LVT U8262 ( .A1(n6901), .A2(n_T_635[62]), .Y(n6851) );
  NAND4X0_LVT U8263 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .Y(
        n_T_702[62]) );
  NAND2X0_LVT U8264 ( .A1(csr_io_rw_rdata[63]), .A2(n3844), .Y(n6864) );
  AOI22X1_LVT U8265 ( .A1(n3852), .A2(io_dmem_resp_bits_data[63]), .A3(n3847), 
        .A4(n_T_1165[63]), .Y(n6863) );
  NAND2X0_LVT U8266 ( .A1(div_io_resp_bits_data[63]), .A2(n3858), .Y(n6862) );
  NAND3X0_LVT U8267 ( .A1(n6864), .A2(n6863), .A3(n6862), .Y(
        n_T_427__T_1136_data[63]) );
  AO22X1_LVT U8268 ( .A1(n_T_427[703]), .A2(n3861), .A3(n3859), .A4(
        n_T_427[255]), .Y(n6875) );
  AO22X1_LVT U8269 ( .A1(n6867), .A2(n_T_427[447]), .A3(n3864), .A4(
        n_T_427[127]), .Y(n6874) );
  AO22X1_LVT U8270 ( .A1(n_T_427[575]), .A2(n3869), .A3(n3866), .A4(
        n_T_427[383]), .Y(n6873) );
  AO22X1_LVT U8271 ( .A1(n_T_427[894]), .A2(n3875), .A3(n3871), .A4(
        n_T_427[319]), .Y(n6872) );
  NOR4X1_LVT U8272 ( .A1(n6875), .A2(n6874), .A3(n6873), .A4(n6872), .Y(n6876)
         );
  OA22X1_LVT U8273 ( .A1(n3529), .A2(n3882), .A3(n3878), .A4(n6876), .Y(n6881)
         );
  NAND2X0_LVT U8274 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[63]), .Y(n6905) );
  NAND2X0_LVT U8275 ( .A1(n6899), .A2(n_T_918[63]), .Y(n6904) );
  NAND2X0_LVT U8276 ( .A1(n_T_1165[63]), .A2(n6900), .Y(n6903) );
  NAND2X0_LVT U8277 ( .A1(n6901), .A2(n_T_635[63]), .Y(n6902) );
  NAND4X0_LVT U8278 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .Y(
        n_T_702[63]) );
  NAND2X0_LVT U8279 ( .A1(ibuf_io_inst_0_bits_rvc), .A2(n6912), .Y(n6913) );
  NAND2X0_LVT U8280 ( .A1(n4001), .A2(n_T_427[1728]), .Y(n6918) );
  OA21X1_LVT U8281 ( .A1(n3747), .A2(n3138), .A3(n6918), .Y(n6921) );
  NAND2X0_LVT U8282 ( .A1(n3648), .A2(n_T_427[1600]), .Y(n6920) );
  NAND2X0_LVT U8283 ( .A1(n3657), .A2(n_T_427[1664]), .Y(n6919) );
  NAND2X0_LVT U8284 ( .A1(n3670), .A2(n_T_427[1088]), .Y(n6925) );
  OA21X1_LVT U8285 ( .A1(n3416), .A2(n2897), .A3(n6925), .Y(n6929) );
  NAND2X0_LVT U8286 ( .A1(n3621), .A2(n_T_427[1536]), .Y(n6928) );
  NAND2X0_LVT U8287 ( .A1(n3641), .A2(n_T_427[1216]), .Y(n6927) );
  NAND2X0_LVT U8288 ( .A1(n2966), .A2(n_T_427[1408]), .Y(n6930) );
  OA21X1_LVT U8289 ( .A1(n3987), .A2(n3654), .A3(n6930), .Y(n6934) );
  NAND2X0_LVT U8290 ( .A1(n3606), .A2(n_T_427[1344]), .Y(n6933) );
  NAND2X0_LVT U8291 ( .A1(n3999), .A2(n_T_427[1280]), .Y(n6932) );
  AND2X1_LVT U8292 ( .A1(n6937), .A2(n6936), .Y(n6938) );
  NAND2X0_LVT U8293 ( .A1(n3991), .A2(n_T_427[1883]), .Y(n6942) );
  NAND2X0_LVT U8294 ( .A1(n3712), .A2(n_T_427[960]), .Y(n6970) );
  AND2X1_LVT U8295 ( .A1(n4051), .A2(n_T_427[1]), .Y(n6953) );
  AO22X1_LVT U8296 ( .A1(n4023), .A2(n_T_427[896]), .A3(n4020), .A4(
        n_T_427[641]), .Y(n6952) );
  AND2X1_LVT U8297 ( .A1(n6974), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n8980) );
  AO22X1_LVT U8298 ( .A1(n3977), .A2(n_T_427[513]), .A3(n4027), .A4(
        n_T_427[832]), .Y(n6951) );
  AO22X1_LVT U8299 ( .A1(n4033), .A2(n_T_427[577]), .A3(n3985), .A4(
        n_T_427[193]), .Y(n6950) );
  NOR4X1_LVT U8300 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .Y(n6968)
         );
  AO22X1_LVT U8301 ( .A1(n3968), .A2(n_T_427[385]), .A3(n3964), .A4(
        n_T_427[257]), .Y(n6961) );
  AO22X1_LVT U8302 ( .A1(n2858), .A2(n_T_427[129]), .A3(n4039), .A4(
        n_T_427[321]), .Y(n6960) );
  AND2X1_LVT U8303 ( .A1(n6954), .A2(n2825), .Y(n8981) );
  AO22X1_LVT U8304 ( .A1(n3981), .A2(n_T_427[768]), .A3(n4047), .A4(
        n_T_427[705]), .Y(n6959) );
  AND2X1_LVT U8305 ( .A1(n6957), .A2(ibuf_io_inst_0_bits_inst_rs1[3]), .Y(
        n8900) );
  AO22X1_LVT U8306 ( .A1(n3962), .A2(n_T_427[449]), .A3(n4044), .A4(
        n_T_427[65]), .Y(n6958) );
  NOR4X1_LVT U8307 ( .A1(n6961), .A2(n6960), .A3(n6959), .A4(n6958), .Y(n6967)
         );
  AND3X1_LVT U8308 ( .A1(n6971), .A2(n6970), .A3(n6969), .Y(n6978) );
  NAND2X0_LVT U8309 ( .A1(n2611), .A2(n_T_427[1152]), .Y(n6977) );
  NAND2X0_LVT U8310 ( .A1(n4014), .A2(n_T_427[1024]), .Y(n6976) );
  NAND2X0_LVT U8311 ( .A1(n4002), .A2(n_T_427[1727]), .Y(n6979) );
  OA21X1_LVT U8312 ( .A1(n3601), .A2(n3311), .A3(n6979), .Y(n6982) );
  NAND2X0_LVT U8313 ( .A1(n3651), .A2(n_T_427[1599]), .Y(n6981) );
  NAND2X0_LVT U8314 ( .A1(n2922), .A2(n_T_427[1663]), .Y(n6980) );
  NAND2X0_LVT U8315 ( .A1(n3671), .A2(n_T_427[1087]), .Y(n6983) );
  OA21X1_LVT U8316 ( .A1(n3417), .A2(n3653), .A3(n6983), .Y(n6986) );
  NAND2X0_LVT U8317 ( .A1(n3616), .A2(n_T_427[1535]), .Y(n6985) );
  NAND2X0_LVT U8318 ( .A1(n3636), .A2(n_T_427[1215]), .Y(n6984) );
  NAND2X0_LVT U8319 ( .A1(n3630), .A2(n_T_427[1407]), .Y(n6987) );
  OA21X1_LVT U8320 ( .A1(n2969), .A2(n3633), .A3(n6987), .Y(n6990) );
  NAND2X0_LVT U8321 ( .A1(n3607), .A2(n_T_427[1343]), .Y(n6989) );
  NAND2X0_LVT U8322 ( .A1(n3997), .A2(n_T_427[1279]), .Y(n6988) );
  NAND3X0_LVT U8323 ( .A1(n6995), .A2(n9288), .A3(n6994), .Y(n6998) );
  NAND2X0_LVT U8324 ( .A1(n2882), .A2(n_T_427[1882]), .Y(n6996) );
  NAND2X0_LVT U8325 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[0]), .Y(n7011)
         );
  NAND2X0_LVT U8326 ( .A1(n3712), .A2(n_T_427[959]), .Y(n7010) );
  AND2X1_LVT U8327 ( .A1(n4049), .A2(n_T_427[0]), .Y(n7002) );
  AO22X1_LVT U8328 ( .A1(n4026), .A2(n_T_427[895]), .A3(n4018), .A4(
        n_T_427[640]), .Y(n7001) );
  AO22X1_LVT U8329 ( .A1(n3976), .A2(n_T_427[512]), .A3(n4030), .A4(
        n_T_427[831]), .Y(n7000) );
  AO22X1_LVT U8330 ( .A1(n4032), .A2(n_T_427[576]), .A3(n3983), .A4(
        n_T_427[192]), .Y(n6999) );
  NOR4X1_LVT U8331 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .Y(n7008)
         );
  AO22X1_LVT U8332 ( .A1(n3968), .A2(n_T_427[384]), .A3(n3964), .A4(
        n_T_427[256]), .Y(n7006) );
  AO22X1_LVT U8333 ( .A1(n3975), .A2(n_T_427[128]), .A3(n4039), .A4(
        n_T_427[320]), .Y(n7005) );
  AO22X1_LVT U8334 ( .A1(n3979), .A2(n_T_427[767]), .A3(n4045), .A4(
        n_T_427[704]), .Y(n7004) );
  AO22X1_LVT U8335 ( .A1(n3960), .A2(n_T_427[448]), .A3(n2837), .A4(
        n_T_427[64]), .Y(n7003) );
  NOR4X1_LVT U8336 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .Y(n7007)
         );
  AND3X1_LVT U8337 ( .A1(n7011), .A2(n7010), .A3(n7009), .Y(n7014) );
  NAND2X0_LVT U8338 ( .A1(n2611), .A2(n_T_427[1151]), .Y(n7013) );
  NAND2X0_LVT U8339 ( .A1(n4014), .A2(n_T_427[1023]), .Y(n7012) );
  OR2X1_LVT U8340 ( .A1(n2497), .A2(n_T_918[0]), .Y(n7015) );
  AND2X1_LVT U8341 ( .A1(n3101), .A2(n_T_628[1]), .Y(n7017) );
  AO22X1_LVT U8342 ( .A1(n7019), .A2(n7015), .A3(n7017), .A4(
        io_imem_sfence_bits_addr[0]), .Y(n7016) );
  NAND2X0_LVT U8343 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[1]), .Y(n7022)
         );
  NAND3X0_LVT U8344 ( .A1(n7019), .A2(n_T_628[1]), .A3(
        io_fpu_dmem_resp_data[1]), .Y(n7018) );
  OA21X1_LVT U8345 ( .A1(n3101), .A2(n3255), .A3(n7018), .Y(n7021) );
  NAND2X0_LVT U8346 ( .A1(n9066), .A2(n_T_918[1]), .Y(n7020) );
  NAND3X0_LVT U8347 ( .A1(n7022), .A2(n7021), .A3(n7020), .Y(
        io_fpu_fromint_data[1]) );
  NAND2X0_LVT U8348 ( .A1(n3997), .A2(n_T_427[1281]), .Y(n7023) );
  OA21X1_LVT U8349 ( .A1(n3377), .A2(n3684), .A3(n7023), .Y(n7026) );
  NAND2X0_LVT U8350 ( .A1(n3990), .A2(n_T_427[1848]), .Y(n7025) );
  NAND2X0_LVT U8351 ( .A1(n_T_427[1792]), .A2(n3715), .Y(n7024) );
  NAND2X0_LVT U8352 ( .A1(n3619), .A2(n_T_427[1537]), .Y(n7027) );
  OA21X1_LVT U8353 ( .A1(n3418), .A2(n3653), .A3(n7027), .Y(n7030) );
  NAND2X0_LVT U8354 ( .A1(n4004), .A2(n_T_427[1729]), .Y(n7029) );
  NAND2X0_LVT U8355 ( .A1(n3652), .A2(n_T_427[1601]), .Y(n7028) );
  NAND2X0_LVT U8356 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[2]), .Y(n7043)
         );
  NAND2X0_LVT U8357 ( .A1(n3717), .A2(n_T_427[1025]), .Y(n7042) );
  AND2X1_LVT U8358 ( .A1(n4049), .A2(n_T_427[2]), .Y(n7034) );
  AO22X1_LVT U8359 ( .A1(n4024), .A2(n_T_427[897]), .A3(n4018), .A4(
        n_T_427[642]), .Y(n7033) );
  AO22X1_LVT U8360 ( .A1(n3976), .A2(n_T_427[514]), .A3(n4030), .A4(
        n_T_427[833]), .Y(n7032) );
  AO22X1_LVT U8361 ( .A1(n4031), .A2(n_T_427[578]), .A3(n3984), .A4(
        n_T_427[194]), .Y(n7031) );
  NOR4X1_LVT U8362 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .Y(n7040)
         );
  AO22X1_LVT U8363 ( .A1(n3968), .A2(n_T_427[386]), .A3(n3964), .A4(
        n_T_427[258]), .Y(n7038) );
  AO22X1_LVT U8364 ( .A1(n2858), .A2(n_T_427[130]), .A3(n4039), .A4(
        n_T_427[322]), .Y(n7037) );
  AO22X1_LVT U8365 ( .A1(n3979), .A2(n_T_427[769]), .A3(n4045), .A4(
        n_T_427[706]), .Y(n7036) );
  AO22X1_LVT U8366 ( .A1(n3960), .A2(n_T_427[450]), .A3(n4043), .A4(
        n_T_427[66]), .Y(n7035) );
  NOR4X1_LVT U8367 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .Y(n7039)
         );
  NAND2X0_LVT U8368 ( .A1(n3639), .A2(n_T_427[1217]), .Y(n7044) );
  NAND2X0_LVT U8369 ( .A1(n3673), .A2(n_T_427[1089]), .Y(n7046) );
  NAND2X0_LVT U8370 ( .A1(n3712), .A2(n_T_427[961]), .Y(n7045) );
  NAND2X0_LVT U8371 ( .A1(n2967), .A2(n_T_427[1409]), .Y(n7047) );
  OA21X1_LVT U8372 ( .A1(n3196), .A2(n2089), .A3(n7047), .Y(n7050) );
  NAND2X0_LVT U8373 ( .A1(n3609), .A2(n_T_427[1345]), .Y(n7049) );
  NAND2X0_LVT U8374 ( .A1(n3992), .A2(n_T_427[1884]), .Y(n7048) );
  NAND2X0_LVT U8375 ( .A1(n3996), .A2(n_T_427[1282]), .Y(n7051) );
  OA21X1_LVT U8376 ( .A1(n3378), .A2(n3684), .A3(n7051), .Y(n7054) );
  NAND2X0_LVT U8377 ( .A1(n_T_427[1849]), .A2(n3764), .Y(n7053) );
  NAND2X0_LVT U8378 ( .A1(n_T_427[1793]), .A2(n3715), .Y(n7052) );
  NAND2X0_LVT U8379 ( .A1(n3620), .A2(n_T_427[1538]), .Y(n7055) );
  OA21X1_LVT U8380 ( .A1(n3420), .A2(n2897), .A3(n7055), .Y(n7058) );
  NAND2X0_LVT U8381 ( .A1(n4004), .A2(n_T_427[1730]), .Y(n7057) );
  NAND2X0_LVT U8382 ( .A1(n3643), .A2(n_T_427[1602]), .Y(n7056) );
  NAND2X0_LVT U8383 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[3]), .Y(n7071)
         );
  NAND2X0_LVT U8384 ( .A1(n4014), .A2(n_T_427[1026]), .Y(n7070) );
  AND2X1_LVT U8385 ( .A1(n4049), .A2(n_T_427[3]), .Y(n7062) );
  AO22X1_LVT U8386 ( .A1(n4025), .A2(n_T_427[898]), .A3(n4018), .A4(
        n_T_427[643]), .Y(n7061) );
  AO22X1_LVT U8387 ( .A1(n3976), .A2(n_T_427[515]), .A3(n4030), .A4(
        n_T_427[834]), .Y(n7060) );
  AO22X1_LVT U8388 ( .A1(n4032), .A2(n_T_427[579]), .A3(n3983), .A4(
        n_T_427[195]), .Y(n7059) );
  NOR4X1_LVT U8389 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .Y(n7068)
         );
  AO22X1_LVT U8390 ( .A1(n3968), .A2(n_T_427[387]), .A3(n3964), .A4(
        n_T_427[259]), .Y(n7066) );
  AO22X1_LVT U8391 ( .A1(n3975), .A2(n_T_427[131]), .A3(n4038), .A4(
        n_T_427[323]), .Y(n7065) );
  AO22X1_LVT U8392 ( .A1(n3980), .A2(n_T_427[770]), .A3(n4045), .A4(
        n_T_427[707]), .Y(n7064) );
  AO22X1_LVT U8393 ( .A1(n3961), .A2(n_T_427[451]), .A3(n4042), .A4(
        n_T_427[67]), .Y(n7063) );
  NOR4X1_LVT U8394 ( .A1(n7066), .A2(n7065), .A3(n7064), .A4(n7063), .Y(n7067)
         );
  NAND2X0_LVT U8395 ( .A1(n_T_427[1218]), .A2(n3639), .Y(n7072) );
  OA21X1_LVT U8396 ( .A1(n3421), .A2(n3664), .A3(n7072), .Y(n7075) );
  NAND2X0_LVT U8397 ( .A1(n3667), .A2(n_T_427[1090]), .Y(n7074) );
  NAND2X0_LVT U8398 ( .A1(n3759), .A2(n_T_427[962]), .Y(n7073) );
  NAND2X0_LVT U8399 ( .A1(n2966), .A2(n_T_427[1410]), .Y(n7076) );
  OA21X1_LVT U8400 ( .A1(n3187), .A2(n2090), .A3(n7076), .Y(n7079) );
  NAND2X0_LVT U8401 ( .A1(n3602), .A2(n_T_427[1346]), .Y(n7078) );
  NAND2X0_LVT U8402 ( .A1(n2093), .A2(n_T_427[1283]), .Y(n7080) );
  OA21X1_LVT U8403 ( .A1(n3379), .A2(n3684), .A3(n7080), .Y(n7083) );
  NAND2X0_LVT U8404 ( .A1(n_T_427[1850]), .A2(n3990), .Y(n7082) );
  NAND2X0_LVT U8405 ( .A1(n_T_427[1794]), .A2(n3715), .Y(n7081) );
  NAND2X0_LVT U8406 ( .A1(n3615), .A2(n_T_427[1539]), .Y(n7084) );
  OA21X1_LVT U8407 ( .A1(n3422), .A2(n3653), .A3(n7084), .Y(n7087) );
  NAND2X0_LVT U8408 ( .A1(n4003), .A2(n_T_427[1731]), .Y(n7086) );
  NAND2X0_LVT U8409 ( .A1(n3643), .A2(n_T_427[1603]), .Y(n7085) );
  NAND2X0_LVT U8410 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[4]), .Y(n7100)
         );
  NAND2X0_LVT U8411 ( .A1(n3716), .A2(n_T_427[1027]), .Y(n7099) );
  AND2X1_LVT U8412 ( .A1(n4049), .A2(n_T_427[4]), .Y(n7091) );
  AO22X1_LVT U8413 ( .A1(n4026), .A2(n_T_427[899]), .A3(n4018), .A4(
        n_T_427[644]), .Y(n7090) );
  AO22X1_LVT U8414 ( .A1(n3976), .A2(n_T_427[516]), .A3(n4030), .A4(
        n_T_427[835]), .Y(n7089) );
  AO22X1_LVT U8415 ( .A1(n4032), .A2(n_T_427[580]), .A3(n3983), .A4(
        n_T_427[196]), .Y(n7088) );
  NOR4X1_LVT U8416 ( .A1(n7091), .A2(n7090), .A3(n7089), .A4(n7088), .Y(n7097)
         );
  AO22X1_LVT U8417 ( .A1(n3968), .A2(n_T_427[388]), .A3(n3964), .A4(
        n_T_427[260]), .Y(n7095) );
  AO22X1_LVT U8418 ( .A1(n2859), .A2(n_T_427[132]), .A3(n9040), .A4(
        n_T_427[324]), .Y(n7094) );
  AO22X1_LVT U8419 ( .A1(n3980), .A2(n_T_427[771]), .A3(n4045), .A4(
        n_T_427[708]), .Y(n7093) );
  AO22X1_LVT U8420 ( .A1(n3961), .A2(n_T_427[452]), .A3(n4042), .A4(
        n_T_427[68]), .Y(n7092) );
  NOR4X1_LVT U8421 ( .A1(n7095), .A2(n7094), .A3(n7093), .A4(n7092), .Y(n7096)
         );
  NAND3X0_LVT U8422 ( .A1(n7100), .A2(n7099), .A3(n7098), .Y(n7107) );
  NAND2X0_LVT U8423 ( .A1(n3674), .A2(n_T_427[1091]), .Y(n7102) );
  NAND2X0_LVT U8424 ( .A1(n3758), .A2(n_T_427[963]), .Y(n7101) );
  NAND2X0_LVT U8425 ( .A1(n_T_427[1347]), .A2(n3611), .Y(n7104) );
  NAND2X0_LVT U8426 ( .A1(n2986), .A2(n_T_427[1885]), .Y(n7103) );
  OR3X1_LVT U8427 ( .A1(n7108), .A2(n7109), .A3(n7110), .Y(N684) );
  NAND2X0_LVT U8428 ( .A1(n3999), .A2(n_T_427[1284]), .Y(n7111) );
  OA21X1_LVT U8429 ( .A1(n3380), .A2(n3684), .A3(n7111), .Y(n7114) );
  NAND2X0_LVT U8430 ( .A1(n_T_427[1851]), .A2(n3764), .Y(n7113) );
  NAND2X0_LVT U8431 ( .A1(n_T_427[1795]), .A2(n3715), .Y(n7112) );
  NAND2X0_LVT U8432 ( .A1(n3616), .A2(n_T_427[1540]), .Y(n7115) );
  OA21X1_LVT U8433 ( .A1(n3423), .A2(n2897), .A3(n7115), .Y(n7118) );
  NAND2X0_LVT U8434 ( .A1(n4002), .A2(n_T_427[1732]), .Y(n7117) );
  NAND2X0_LVT U8435 ( .A1(n3642), .A2(n_T_427[1604]), .Y(n7116) );
  NAND2X0_LVT U8436 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[5]), .Y(n7131)
         );
  NAND2X0_LVT U8437 ( .A1(n3717), .A2(n_T_427[1028]), .Y(n7130) );
  AND2X1_LVT U8438 ( .A1(n4049), .A2(n_T_427[5]), .Y(n7122) );
  AO22X1_LVT U8439 ( .A1(n4026), .A2(n_T_427[900]), .A3(n4018), .A4(
        n_T_427[645]), .Y(n7121) );
  AO22X1_LVT U8440 ( .A1(n3976), .A2(n_T_427[517]), .A3(n4030), .A4(
        n_T_427[836]), .Y(n7120) );
  AO22X1_LVT U8441 ( .A1(n4032), .A2(n_T_427[581]), .A3(n3984), .A4(
        n_T_427[197]), .Y(n7119) );
  NOR4X1_LVT U8442 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .Y(n7128)
         );
  AO22X1_LVT U8443 ( .A1(n3968), .A2(n_T_427[389]), .A3(n3964), .A4(
        n_T_427[261]), .Y(n7126) );
  AO22X1_LVT U8444 ( .A1(n3974), .A2(n_T_427[133]), .A3(n4037), .A4(
        n_T_427[325]), .Y(n7125) );
  AO22X1_LVT U8445 ( .A1(n3980), .A2(n_T_427[772]), .A3(n4045), .A4(
        n_T_427[709]), .Y(n7124) );
  AO22X1_LVT U8446 ( .A1(n3961), .A2(n_T_427[453]), .A3(n4042), .A4(
        n_T_427[69]), .Y(n7123) );
  NOR4X1_LVT U8447 ( .A1(n7126), .A2(n7125), .A3(n7124), .A4(n7123), .Y(n7127)
         );
  AO21X1_LVT U8448 ( .A1(n7128), .A2(n7127), .A3(n2645), .Y(n7129) );
  NAND2X0_LVT U8449 ( .A1(n3641), .A2(n_T_427[1220]), .Y(n7132) );
  NAND2X0_LVT U8450 ( .A1(n3674), .A2(n_T_427[1092]), .Y(n7134) );
  NAND2X0_LVT U8451 ( .A1(n3756), .A2(n_T_427[964]), .Y(n7133) );
  NAND2X0_LVT U8452 ( .A1(n3629), .A2(n_T_427[1412]), .Y(n7135) );
  OA21X1_LVT U8453 ( .A1(n3197), .A2(n2089), .A3(n7135), .Y(n7138) );
  NAND2X0_LVT U8454 ( .A1(n3608), .A2(n_T_427[1348]), .Y(n7137) );
  NAND2X0_LVT U8455 ( .A1(n2986), .A2(n_T_427[1886]), .Y(n7136) );
  NAND2X0_LVT U8456 ( .A1(n4000), .A2(n_T_427[1285]), .Y(n7139) );
  OA21X1_LVT U8457 ( .A1(n3381), .A2(n3684), .A3(n7139), .Y(n7142) );
  NAND2X0_LVT U8458 ( .A1(n_T_427[1852]), .A2(n3990), .Y(n7141) );
  NAND2X0_LVT U8459 ( .A1(n_T_427[1796]), .A2(n3715), .Y(n7140) );
  NAND2X0_LVT U8460 ( .A1(n3617), .A2(n_T_427[1541]), .Y(n7143) );
  OA21X1_LVT U8461 ( .A1(n3425), .A2(n3653), .A3(n7143), .Y(n7146) );
  NAND2X0_LVT U8462 ( .A1(n4002), .A2(n_T_427[1733]), .Y(n7145) );
  NAND2X0_LVT U8463 ( .A1(n3651), .A2(n_T_427[1605]), .Y(n7144) );
  NAND2X0_LVT U8464 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[6]), .Y(n7159)
         );
  NAND2X0_LVT U8465 ( .A1(n4014), .A2(n_T_427[1029]), .Y(n7158) );
  AND2X1_LVT U8466 ( .A1(n4049), .A2(n_T_427[6]), .Y(n7150) );
  AO22X1_LVT U8467 ( .A1(n4023), .A2(n_T_427[901]), .A3(n4018), .A4(
        n_T_427[646]), .Y(n7149) );
  AO22X1_LVT U8468 ( .A1(n3977), .A2(n_T_427[518]), .A3(n4030), .A4(
        n_T_427[837]), .Y(n7148) );
  AO22X1_LVT U8469 ( .A1(n4032), .A2(n_T_427[582]), .A3(n3983), .A4(
        n_T_427[198]), .Y(n7147) );
  NOR4X1_LVT U8470 ( .A1(n7150), .A2(n7149), .A3(n7148), .A4(n7147), .Y(n7156)
         );
  AO22X1_LVT U8471 ( .A1(n3968), .A2(n_T_427[390]), .A3(n3964), .A4(
        n_T_427[262]), .Y(n7154) );
  AO22X1_LVT U8472 ( .A1(n2859), .A2(n_T_427[134]), .A3(n4039), .A4(
        n_T_427[326]), .Y(n7153) );
  AO22X1_LVT U8473 ( .A1(n3980), .A2(n_T_427[773]), .A3(n4045), .A4(
        n_T_427[710]), .Y(n7152) );
  AO22X1_LVT U8474 ( .A1(n3961), .A2(n_T_427[454]), .A3(n4041), .A4(
        n_T_427[70]), .Y(n7151) );
  NOR4X1_LVT U8475 ( .A1(n7154), .A2(n7153), .A3(n7152), .A4(n7151), .Y(n7155)
         );
  AO21X1_LVT U8476 ( .A1(n7156), .A2(n7155), .A3(n2154), .Y(n7157) );
  NAND2X0_LVT U8477 ( .A1(n_T_427[1221]), .A2(n3640), .Y(n7160) );
  OA21X1_LVT U8478 ( .A1(n3426), .A2(n2081), .A3(n7160), .Y(n7163) );
  NAND2X0_LVT U8479 ( .A1(n3675), .A2(n_T_427[1093]), .Y(n7162) );
  NAND2X0_LVT U8480 ( .A1(n3760), .A2(n_T_427[965]), .Y(n7161) );
  NAND2X0_LVT U8481 ( .A1(n3629), .A2(n_T_427[1413]), .Y(n7164) );
  OA21X1_LVT U8482 ( .A1(n3194), .A2(n2090), .A3(n7164), .Y(n7167) );
  NAND2X0_LVT U8483 ( .A1(n3605), .A2(n_T_427[1349]), .Y(n7166) );
  NAND2X0_LVT U8484 ( .A1(n2985), .A2(n_T_427[1887]), .Y(n7165) );
  NAND2X0_LVT U8485 ( .A1(n2093), .A2(n_T_427[1286]), .Y(n7168) );
  OA21X1_LVT U8486 ( .A1(n3382), .A2(n3684), .A3(n7168), .Y(n7171) );
  NAND2X0_LVT U8487 ( .A1(n_T_427[1853]), .A2(n3990), .Y(n7170) );
  NAND2X0_LVT U8488 ( .A1(n_T_427[1797]), .A2(n3715), .Y(n7169) );
  NAND2X0_LVT U8489 ( .A1(n3618), .A2(n_T_427[1542]), .Y(n7172) );
  NAND2X0_LVT U8490 ( .A1(n4005), .A2(n_T_427[1734]), .Y(n7174) );
  NAND2X0_LVT U8491 ( .A1(n3651), .A2(n_T_427[1606]), .Y(n7173) );
  NAND2X0_LVT U8492 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[7]), .Y(n7187)
         );
  NAND2X0_LVT U8493 ( .A1(n3717), .A2(n_T_427[1030]), .Y(n7186) );
  AND2X1_LVT U8494 ( .A1(n4049), .A2(n_T_427[7]), .Y(n7178) );
  AO22X1_LVT U8495 ( .A1(n4026), .A2(n_T_427[902]), .A3(n4018), .A4(
        n_T_427[647]), .Y(n7177) );
  AO22X1_LVT U8496 ( .A1(n3977), .A2(n_T_427[519]), .A3(n4030), .A4(
        n_T_427[838]), .Y(n7176) );
  AO22X1_LVT U8497 ( .A1(n4032), .A2(n_T_427[583]), .A3(n3983), .A4(
        n_T_427[199]), .Y(n7175) );
  NOR4X1_LVT U8498 ( .A1(n7178), .A2(n7177), .A3(n7176), .A4(n7175), .Y(n7184)
         );
  AO22X1_LVT U8499 ( .A1(n3968), .A2(n_T_427[391]), .A3(n3964), .A4(
        n_T_427[263]), .Y(n7182) );
  AO22X1_LVT U8500 ( .A1(n3975), .A2(n_T_427[135]), .A3(n4037), .A4(
        n_T_427[327]), .Y(n7181) );
  AO22X1_LVT U8501 ( .A1(n3980), .A2(n_T_427[774]), .A3(n4045), .A4(
        n_T_427[711]), .Y(n7180) );
  AO22X1_LVT U8502 ( .A1(n3961), .A2(n_T_427[455]), .A3(n4043), .A4(
        n_T_427[71]), .Y(n7179) );
  NOR4X1_LVT U8503 ( .A1(n7182), .A2(n7181), .A3(n7180), .A4(n7179), .Y(n7183)
         );
  AO21X1_LVT U8504 ( .A1(n7184), .A2(n7183), .A3(n3631), .Y(n7185) );
  NAND2X0_LVT U8505 ( .A1(n_T_427[1222]), .A2(n3638), .Y(n7188) );
  NAND2X0_LVT U8506 ( .A1(n3667), .A2(n_T_427[1094]), .Y(n7190) );
  NAND2X0_LVT U8507 ( .A1(n3756), .A2(n_T_427[966]), .Y(n7189) );
  NAND2X0_LVT U8508 ( .A1(n2967), .A2(n_T_427[1414]), .Y(n7191) );
  NAND2X0_LVT U8509 ( .A1(n3607), .A2(n_T_427[1350]), .Y(n7193) );
  NAND2X0_LVT U8510 ( .A1(n2985), .A2(n_T_427[1888]), .Y(n7192) );
  NAND2X0_LVT U8511 ( .A1(n4000), .A2(n_T_427[1287]), .Y(n7194) );
  OA21X1_LVT U8512 ( .A1(n3383), .A2(n3684), .A3(n7194), .Y(n7197) );
  NAND2X0_LVT U8513 ( .A1(n_T_427[1854]), .A2(n3764), .Y(n7196) );
  NAND2X0_LVT U8514 ( .A1(n_T_427[1798]), .A2(n3715), .Y(n7195) );
  NAND2X0_LVT U8515 ( .A1(n3619), .A2(n_T_427[1543]), .Y(n7198) );
  OA21X1_LVT U8516 ( .A1(n3429), .A2(n2897), .A3(n7198), .Y(n7201) );
  NAND2X0_LVT U8517 ( .A1(n4001), .A2(n_T_427[1735]), .Y(n7200) );
  NAND2X0_LVT U8518 ( .A1(n3643), .A2(n_T_427[1607]), .Y(n7199) );
  NAND2X0_LVT U8519 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[8]), .Y(n7214)
         );
  NAND2X0_LVT U8520 ( .A1(n3716), .A2(n_T_427[1031]), .Y(n7213) );
  AND2X1_LVT U8521 ( .A1(n4049), .A2(n_T_427[8]), .Y(n7205) );
  AO22X1_LVT U8522 ( .A1(n4026), .A2(n_T_427[903]), .A3(n4018), .A4(
        n_T_427[648]), .Y(n7204) );
  AO22X1_LVT U8523 ( .A1(n3977), .A2(n_T_427[520]), .A3(n4030), .A4(
        n_T_427[839]), .Y(n7203) );
  AO22X1_LVT U8524 ( .A1(n4032), .A2(n_T_427[584]), .A3(n3983), .A4(
        n_T_427[200]), .Y(n7202) );
  NOR4X1_LVT U8525 ( .A1(n7205), .A2(n7204), .A3(n7203), .A4(n7202), .Y(n7211)
         );
  AO22X1_LVT U8526 ( .A1(n3968), .A2(n_T_427[392]), .A3(n3964), .A4(
        n_T_427[264]), .Y(n7209) );
  AO22X1_LVT U8527 ( .A1(n3974), .A2(n_T_427[136]), .A3(n4039), .A4(
        n_T_427[328]), .Y(n7208) );
  AO22X1_LVT U8528 ( .A1(n3980), .A2(n_T_427[775]), .A3(n4045), .A4(
        n_T_427[712]), .Y(n7207) );
  AO22X1_LVT U8529 ( .A1(n3961), .A2(n_T_427[456]), .A3(n4044), .A4(
        n_T_427[72]), .Y(n7206) );
  NOR4X1_LVT U8530 ( .A1(n7209), .A2(n7208), .A3(n7207), .A4(n7206), .Y(n7210)
         );
  AO21X1_LVT U8531 ( .A1(n7211), .A2(n7210), .A3(n3656), .Y(n7212) );
  NAND2X0_LVT U8532 ( .A1(n3637), .A2(n_T_427[1223]), .Y(n7215) );
  OA21X1_LVT U8533 ( .A1(n3430), .A2(n4010), .A3(n7215), .Y(n7218) );
  NAND2X0_LVT U8534 ( .A1(n3675), .A2(n_T_427[1095]), .Y(n7217) );
  NAND2X0_LVT U8535 ( .A1(n3756), .A2(n_T_427[967]), .Y(n7216) );
  NAND2X0_LVT U8536 ( .A1(n3629), .A2(n_T_427[1415]), .Y(n7219) );
  OA21X1_LVT U8537 ( .A1(n3192), .A2(n2089), .A3(n7219), .Y(n7222) );
  NAND2X0_LVT U8538 ( .A1(n3608), .A2(n_T_427[1351]), .Y(n7221) );
  NAND2X0_LVT U8539 ( .A1(n2986), .A2(n_T_427[1889]), .Y(n7220) );
  NAND2X0_LVT U8540 ( .A1(n2093), .A2(n_T_427[1288]), .Y(n7223) );
  OA21X1_LVT U8541 ( .A1(n3384), .A2(n3684), .A3(n7223), .Y(n7226) );
  NAND2X0_LVT U8542 ( .A1(n_T_427[1855]), .A2(n3990), .Y(n7225) );
  NAND2X0_LVT U8543 ( .A1(n_T_427[1799]), .A2(n3715), .Y(n7224) );
  NAND2X0_LVT U8544 ( .A1(n3620), .A2(n_T_427[1544]), .Y(n7227) );
  OA21X1_LVT U8545 ( .A1(n3431), .A2(n2897), .A3(n7227), .Y(n7230) );
  NAND2X0_LVT U8546 ( .A1(n4001), .A2(n_T_427[1736]), .Y(n7229) );
  NAND2X0_LVT U8547 ( .A1(n3652), .A2(n_T_427[1608]), .Y(n7228) );
  NAND2X0_LVT U8548 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[9]), .Y(n7243)
         );
  NAND2X0_LVT U8549 ( .A1(n4014), .A2(n_T_427[1032]), .Y(n7242) );
  AND2X1_LVT U8550 ( .A1(n4049), .A2(n_T_427[9]), .Y(n7234) );
  AO22X1_LVT U8551 ( .A1(n4026), .A2(n_T_427[904]), .A3(n4019), .A4(
        n_T_427[649]), .Y(n7233) );
  AO22X1_LVT U8552 ( .A1(n3977), .A2(n_T_427[521]), .A3(n4029), .A4(
        n_T_427[840]), .Y(n7232) );
  AO22X1_LVT U8553 ( .A1(n4032), .A2(n_T_427[585]), .A3(n3984), .A4(
        n_T_427[201]), .Y(n7231) );
  NOR4X1_LVT U8554 ( .A1(n7234), .A2(n7233), .A3(n7232), .A4(n7231), .Y(n7240)
         );
  AO22X1_LVT U8555 ( .A1(n3969), .A2(n_T_427[393]), .A3(n3965), .A4(
        n_T_427[265]), .Y(n7238) );
  AO22X1_LVT U8556 ( .A1(n3975), .A2(n_T_427[137]), .A3(n4039), .A4(
        n_T_427[329]), .Y(n7237) );
  AO22X1_LVT U8557 ( .A1(n3980), .A2(n_T_427[776]), .A3(n4045), .A4(
        n_T_427[713]), .Y(n7236) );
  AO22X1_LVT U8558 ( .A1(n3961), .A2(n_T_427[457]), .A3(n2837), .A4(
        n_T_427[73]), .Y(n7235) );
  NOR4X1_LVT U8559 ( .A1(n7238), .A2(n7237), .A3(n7236), .A4(n7235), .Y(n7239)
         );
  AO21X1_LVT U8560 ( .A1(n7240), .A2(n7239), .A3(n2155), .Y(n7241) );
  NAND2X0_LVT U8561 ( .A1(n3636), .A2(n_T_427[1224]), .Y(n7244) );
  NAND2X0_LVT U8562 ( .A1(n3672), .A2(n_T_427[1096]), .Y(n7246) );
  NAND2X0_LVT U8563 ( .A1(n3761), .A2(n_T_427[968]), .Y(n7245) );
  NAND2X0_LVT U8564 ( .A1(n3626), .A2(n_T_427[1416]), .Y(n7247) );
  NAND2X0_LVT U8565 ( .A1(n2882), .A2(n_T_427[1890]), .Y(n7248) );
  NAND2X0_LVT U8566 ( .A1(n3998), .A2(n_T_427[1289]), .Y(n7249) );
  OA21X1_LVT U8567 ( .A1(n3385), .A2(n3684), .A3(n7249), .Y(n7252) );
  NAND2X0_LVT U8568 ( .A1(n_T_427[1856]), .A2(n3764), .Y(n7251) );
  NAND2X0_LVT U8569 ( .A1(n_T_427[1800]), .A2(n3715), .Y(n7250) );
  NAND2X0_LVT U8570 ( .A1(n3621), .A2(n_T_427[1545]), .Y(n7253) );
  OA21X1_LVT U8571 ( .A1(n3433), .A2(n3653), .A3(n7253), .Y(n7256) );
  NAND2X0_LVT U8572 ( .A1(n2091), .A2(n_T_427[1737]), .Y(n7255) );
  NAND2X0_LVT U8573 ( .A1(n3648), .A2(n_T_427[1609]), .Y(n7254) );
  NAND2X0_LVT U8574 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[10]), .Y(n7269)
         );
  NAND2X0_LVT U8575 ( .A1(n3717), .A2(n_T_427[1033]), .Y(n7268) );
  AND2X1_LVT U8576 ( .A1(n4049), .A2(n_T_427[10]), .Y(n7260) );
  AO22X1_LVT U8577 ( .A1(n4026), .A2(n_T_427[905]), .A3(n4018), .A4(
        n_T_427[650]), .Y(n7259) );
  AO22X1_LVT U8578 ( .A1(n3977), .A2(n_T_427[522]), .A3(n4029), .A4(
        n_T_427[841]), .Y(n7258) );
  AO22X1_LVT U8579 ( .A1(n4032), .A2(n_T_427[586]), .A3(n3984), .A4(
        n_T_427[202]), .Y(n7257) );
  NOR4X1_LVT U8580 ( .A1(n7260), .A2(n7259), .A3(n7258), .A4(n7257), .Y(n7266)
         );
  AO22X1_LVT U8581 ( .A1(n3968), .A2(n_T_427[394]), .A3(n3964), .A4(
        n_T_427[266]), .Y(n7264) );
  AO22X1_LVT U8582 ( .A1(n3973), .A2(n_T_427[138]), .A3(n4039), .A4(
        n_T_427[330]), .Y(n7263) );
  AO22X1_LVT U8583 ( .A1(n3980), .A2(n_T_427[777]), .A3(n4045), .A4(
        n_T_427[714]), .Y(n7262) );
  AO22X1_LVT U8584 ( .A1(n3961), .A2(n_T_427[458]), .A3(n2836), .A4(
        n_T_427[74]), .Y(n7261) );
  NOR4X1_LVT U8585 ( .A1(n7264), .A2(n7263), .A3(n7262), .A4(n7261), .Y(n7265)
         );
  AO21X1_LVT U8586 ( .A1(n7266), .A2(n7265), .A3(n2645), .Y(n7267) );
  NAND2X0_LVT U8587 ( .A1(n3637), .A2(n_T_427[1225]), .Y(n7270) );
  OA21X1_LVT U8588 ( .A1(n3434), .A2(n3664), .A3(n7270), .Y(n7273) );
  NAND2X0_LVT U8589 ( .A1(n3671), .A2(n_T_427[1097]), .Y(n7272) );
  NAND2X0_LVT U8590 ( .A1(n3757), .A2(n_T_427[969]), .Y(n7271) );
  NAND2X0_LVT U8591 ( .A1(n2966), .A2(n_T_427[1417]), .Y(n7274) );
  OA21X1_LVT U8592 ( .A1(n3188), .A2(n2090), .A3(n7274), .Y(n7277) );
  NAND2X0_LVT U8593 ( .A1(n3602), .A2(n_T_427[1353]), .Y(n7276) );
  NAND2X0_LVT U8594 ( .A1(n2998), .A2(n_T_427[1891]), .Y(n7275) );
  NAND2X0_LVT U8595 ( .A1(n4000), .A2(n_T_427[1290]), .Y(n7278) );
  OA21X1_LVT U8596 ( .A1(n3435), .A2(n3684), .A3(n7278), .Y(n7281) );
  NAND2X0_LVT U8597 ( .A1(n_T_427[1857]), .A2(n3764), .Y(n7280) );
  NAND2X0_LVT U8598 ( .A1(n_T_427[1801]), .A2(n3715), .Y(n7279) );
  NAND2X0_LVT U8599 ( .A1(n3619), .A2(n_T_427[1546]), .Y(n7282) );
  OA21X1_LVT U8600 ( .A1(n3386), .A2(n3653), .A3(n7282), .Y(n7285) );
  NAND2X0_LVT U8601 ( .A1(n2092), .A2(n_T_427[1738]), .Y(n7284) );
  NAND2X0_LVT U8602 ( .A1(n3642), .A2(n_T_427[1610]), .Y(n7283) );
  NAND2X0_LVT U8603 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[11]), .Y(n7298)
         );
  NAND2X0_LVT U8604 ( .A1(n4014), .A2(n_T_427[1034]), .Y(n7297) );
  AND2X1_LVT U8605 ( .A1(n4049), .A2(n_T_427[11]), .Y(n7289) );
  AO22X1_LVT U8606 ( .A1(n4026), .A2(n_T_427[906]), .A3(n4019), .A4(
        n_T_427[651]), .Y(n7288) );
  AO22X1_LVT U8607 ( .A1(n3977), .A2(n_T_427[523]), .A3(n4029), .A4(
        n_T_427[842]), .Y(n7287) );
  AO22X1_LVT U8608 ( .A1(n4032), .A2(n_T_427[587]), .A3(n3984), .A4(
        n_T_427[203]), .Y(n7286) );
  NOR4X1_LVT U8609 ( .A1(n7289), .A2(n7288), .A3(n7287), .A4(n7286), .Y(n7295)
         );
  AO22X1_LVT U8610 ( .A1(n3969), .A2(n_T_427[395]), .A3(n3964), .A4(
        n_T_427[267]), .Y(n7293) );
  AO22X1_LVT U8611 ( .A1(n3973), .A2(n_T_427[139]), .A3(n4037), .A4(
        n_T_427[331]), .Y(n7292) );
  AO22X1_LVT U8612 ( .A1(n3980), .A2(n_T_427[778]), .A3(n4045), .A4(
        n_T_427[715]), .Y(n7291) );
  AO22X1_LVT U8613 ( .A1(n3961), .A2(n_T_427[459]), .A3(n4042), .A4(
        n_T_427[75]), .Y(n7290) );
  NOR4X1_LVT U8614 ( .A1(n7293), .A2(n7292), .A3(n7291), .A4(n7290), .Y(n7294)
         );
  AO21X1_LVT U8615 ( .A1(n7295), .A2(n7294), .A3(n3631), .Y(n7296) );
  NAND2X0_LVT U8616 ( .A1(n3667), .A2(n_T_427[1098]), .Y(n7300) );
  NAND2X0_LVT U8617 ( .A1(n3758), .A2(n_T_427[970]), .Y(n7299) );
  NAND2X0_LVT U8618 ( .A1(n3630), .A2(n_T_427[1418]), .Y(n7302) );
  NAND2X0_LVT U8619 ( .A1(n3603), .A2(n_T_427[1354]), .Y(n7304) );
  NAND2X0_LVT U8620 ( .A1(n2985), .A2(n_T_427[1892]), .Y(n7303) );
  NAND2X0_LVT U8621 ( .A1(n2093), .A2(n_T_427[1291]), .Y(n7305) );
  OA21X1_LVT U8622 ( .A1(n3387), .A2(n3684), .A3(n7305), .Y(n7308) );
  NAND2X0_LVT U8623 ( .A1(n_T_427[1858]), .A2(n3990), .Y(n7307) );
  NAND2X0_LVT U8624 ( .A1(n_T_427[1802]), .A2(n3995), .Y(n7306) );
  NAND2X0_LVT U8625 ( .A1(n3615), .A2(n_T_427[1547]), .Y(n7309) );
  OA21X1_LVT U8626 ( .A1(n3436), .A2(n2897), .A3(n7309), .Y(n7312) );
  NAND2X0_LVT U8627 ( .A1(n4005), .A2(n_T_427[1739]), .Y(n7311) );
  NAND2X0_LVT U8628 ( .A1(n3648), .A2(n_T_427[1611]), .Y(n7310) );
  NAND2X0_LVT U8629 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[12]), .Y(n7325)
         );
  NAND2X0_LVT U8630 ( .A1(n3716), .A2(n_T_427[1035]), .Y(n7324) );
  AND2X1_LVT U8631 ( .A1(n4049), .A2(n_T_427[12]), .Y(n7316) );
  AO22X1_LVT U8632 ( .A1(n4026), .A2(n_T_427[907]), .A3(n4019), .A4(
        n_T_427[652]), .Y(n7315) );
  AO22X1_LVT U8633 ( .A1(n3977), .A2(n_T_427[524]), .A3(n4029), .A4(
        n_T_427[843]), .Y(n7314) );
  AO22X1_LVT U8634 ( .A1(n4032), .A2(n_T_427[588]), .A3(n3984), .A4(
        n_T_427[204]), .Y(n7313) );
  NOR4X1_LVT U8635 ( .A1(n7316), .A2(n7315), .A3(n7314), .A4(n7313), .Y(n7322)
         );
  AO22X1_LVT U8636 ( .A1(n3968), .A2(n_T_427[396]), .A3(n3965), .A4(
        n_T_427[268]), .Y(n7320) );
  AO22X1_LVT U8637 ( .A1(n3973), .A2(n_T_427[140]), .A3(n4036), .A4(
        n_T_427[332]), .Y(n7319) );
  AO22X1_LVT U8638 ( .A1(n3980), .A2(n_T_427[779]), .A3(n4046), .A4(
        n_T_427[716]), .Y(n7318) );
  AO22X1_LVT U8639 ( .A1(n3961), .A2(n_T_427[460]), .A3(n4044), .A4(
        n_T_427[76]), .Y(n7317) );
  NOR4X1_LVT U8640 ( .A1(n7320), .A2(n7319), .A3(n7318), .A4(n7317), .Y(n7321)
         );
  NAND2X0_LVT U8641 ( .A1(n_T_427[1227]), .A2(n3640), .Y(n7326) );
  OA21X1_LVT U8642 ( .A1(n3437), .A2(n4008), .A3(n7326), .Y(n7329) );
  NAND2X0_LVT U8643 ( .A1(n3674), .A2(n_T_427[1099]), .Y(n7328) );
  NAND2X0_LVT U8644 ( .A1(n3761), .A2(n_T_427[971]), .Y(n7327) );
  NAND2X0_LVT U8645 ( .A1(n2966), .A2(n_T_427[1419]), .Y(n7330) );
  OA21X1_LVT U8646 ( .A1(n3193), .A2(n2089), .A3(n7330), .Y(n7333) );
  NAND2X0_LVT U8647 ( .A1(n3604), .A2(n_T_427[1355]), .Y(n7332) );
  NAND2X0_LVT U8648 ( .A1(n2986), .A2(n_T_427[1893]), .Y(n7331) );
  NAND2X0_LVT U8649 ( .A1(n2094), .A2(n_T_427[1292]), .Y(n7334) );
  OA21X1_LVT U8650 ( .A1(n3388), .A2(n3684), .A3(n7334), .Y(n7337) );
  NAND2X0_LVT U8651 ( .A1(n_T_427[1859]), .A2(n3990), .Y(n7336) );
  NAND2X0_LVT U8652 ( .A1(n_T_427[1803]), .A2(n3995), .Y(n7335) );
  NAND2X0_LVT U8653 ( .A1(n3616), .A2(n_T_427[1548]), .Y(n7338) );
  OA21X1_LVT U8654 ( .A1(n3438), .A2(n3653), .A3(n7338), .Y(n7341) );
  NAND2X0_LVT U8655 ( .A1(n2092), .A2(n_T_427[1740]), .Y(n7340) );
  NAND2X0_LVT U8656 ( .A1(n3652), .A2(n_T_427[1612]), .Y(n7339) );
  NAND2X0_LVT U8657 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[13]), .Y(n7354)
         );
  NAND2X0_LVT U8658 ( .A1(n3716), .A2(n_T_427[1036]), .Y(n7353) );
  AND2X1_LVT U8659 ( .A1(n4050), .A2(n_T_427[13]), .Y(n7345) );
  AO22X1_LVT U8660 ( .A1(n4026), .A2(n_T_427[908]), .A3(n4019), .A4(
        n_T_427[653]), .Y(n7344) );
  AO22X1_LVT U8661 ( .A1(n3977), .A2(n_T_427[525]), .A3(n4029), .A4(
        n_T_427[844]), .Y(n7343) );
  AO22X1_LVT U8662 ( .A1(n4032), .A2(n_T_427[589]), .A3(n3984), .A4(
        n_T_427[205]), .Y(n7342) );
  NOR4X1_LVT U8663 ( .A1(n7345), .A2(n7344), .A3(n7343), .A4(n7342), .Y(n7351)
         );
  AO22X1_LVT U8664 ( .A1(n3969), .A2(n_T_427[397]), .A3(n3965), .A4(
        n_T_427[269]), .Y(n7349) );
  AO22X1_LVT U8665 ( .A1(n3974), .A2(n_T_427[141]), .A3(n4037), .A4(
        n_T_427[333]), .Y(n7348) );
  AO22X1_LVT U8666 ( .A1(n3980), .A2(n_T_427[780]), .A3(n4046), .A4(
        n_T_427[717]), .Y(n7347) );
  AO22X1_LVT U8667 ( .A1(n3961), .A2(n_T_427[461]), .A3(n2836), .A4(
        n_T_427[77]), .Y(n7346) );
  NOR4X1_LVT U8668 ( .A1(n7349), .A2(n7348), .A3(n7347), .A4(n7346), .Y(n7350)
         );
  NAND2X0_LVT U8669 ( .A1(n_T_427[1228]), .A2(n3638), .Y(n7355) );
  NAND2X0_LVT U8670 ( .A1(n_T_427[1100]), .A2(n3674), .Y(n7357) );
  NAND2X0_LVT U8671 ( .A1(n3757), .A2(n_T_427[972]), .Y(n7356) );
  NAND2X0_LVT U8672 ( .A1(n3610), .A2(n_T_427[1356]), .Y(n7359) );
  NAND2X0_LVT U8673 ( .A1(n2998), .A2(n_T_427[1894]), .Y(n7358) );
  NAND2X0_LVT U8674 ( .A1(n3998), .A2(n_T_427[1293]), .Y(n7361) );
  OA21X1_LVT U8675 ( .A1(n3389), .A2(n3684), .A3(n7361), .Y(n7364) );
  NAND2X0_LVT U8676 ( .A1(n_T_427[1860]), .A2(n3990), .Y(n7363) );
  NAND2X0_LVT U8677 ( .A1(n_T_427[1804]), .A2(n3995), .Y(n7362) );
  NAND2X0_LVT U8678 ( .A1(n3617), .A2(n_T_427[1549]), .Y(n7365) );
  OA21X1_LVT U8679 ( .A1(n3440), .A2(n2897), .A3(n7365), .Y(n7368) );
  NAND2X0_LVT U8680 ( .A1(n4001), .A2(n_T_427[1741]), .Y(n7367) );
  NAND2X0_LVT U8681 ( .A1(n3651), .A2(n_T_427[1613]), .Y(n7366) );
  NAND2X0_LVT U8682 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[14]), .Y(n7381)
         );
  NAND2X0_LVT U8683 ( .A1(n3716), .A2(n_T_427[1037]), .Y(n7380) );
  AND2X1_LVT U8684 ( .A1(n4050), .A2(n_T_427[14]), .Y(n7372) );
  AO22X1_LVT U8685 ( .A1(n4026), .A2(n_T_427[909]), .A3(n4019), .A4(
        n_T_427[654]), .Y(n7371) );
  AO22X1_LVT U8686 ( .A1(n3977), .A2(n_T_427[526]), .A3(n4029), .A4(
        n_T_427[845]), .Y(n7370) );
  AO22X1_LVT U8687 ( .A1(n4032), .A2(n_T_427[590]), .A3(n3984), .A4(
        n_T_427[206]), .Y(n7369) );
  NOR4X1_LVT U8688 ( .A1(n7372), .A2(n7371), .A3(n7370), .A4(n7369), .Y(n7378)
         );
  AO22X1_LVT U8689 ( .A1(n3969), .A2(n_T_427[398]), .A3(n3965), .A4(
        n_T_427[270]), .Y(n7376) );
  AO22X1_LVT U8690 ( .A1(n2859), .A2(n_T_427[142]), .A3(n4036), .A4(
        n_T_427[334]), .Y(n7375) );
  AO22X1_LVT U8691 ( .A1(n3980), .A2(n_T_427[781]), .A3(n4046), .A4(
        n_T_427[718]), .Y(n7374) );
  AO22X1_LVT U8692 ( .A1(n3961), .A2(n_T_427[462]), .A3(n2837), .A4(
        n_T_427[78]), .Y(n7373) );
  NOR4X1_LVT U8693 ( .A1(n7376), .A2(n7375), .A3(n7374), .A4(n7373), .Y(n7377)
         );
  NAND2X0_LVT U8694 ( .A1(n_T_427[1229]), .A2(n3636), .Y(n7382) );
  OA21X1_LVT U8695 ( .A1(n3441), .A2(n3664), .A3(n7382), .Y(n7385) );
  NAND2X0_LVT U8696 ( .A1(n3673), .A2(n_T_427[1101]), .Y(n7384) );
  NAND2X0_LVT U8697 ( .A1(n3758), .A2(n_T_427[973]), .Y(n7383) );
  NAND2X0_LVT U8698 ( .A1(n3629), .A2(n_T_427[1421]), .Y(n7386) );
  OA21X1_LVT U8699 ( .A1(n3195), .A2(n2089), .A3(n7386), .Y(n7389) );
  NAND2X0_LVT U8700 ( .A1(n3604), .A2(n_T_427[1357]), .Y(n7388) );
  NAND2X0_LVT U8701 ( .A1(n3992), .A2(n_T_427[1895]), .Y(n7387) );
  NAND2X0_LVT U8702 ( .A1(n3996), .A2(n_T_427[1294]), .Y(n7390) );
  OA21X1_LVT U8703 ( .A1(n3390), .A2(n3684), .A3(n7390), .Y(n7393) );
  NAND2X0_LVT U8704 ( .A1(n_T_427[1861]), .A2(n3764), .Y(n7392) );
  NAND2X0_LVT U8705 ( .A1(n_T_427[1805]), .A2(n3995), .Y(n7391) );
  NAND2X0_LVT U8706 ( .A1(n3618), .A2(n_T_427[1550]), .Y(n7394) );
  OA21X1_LVT U8707 ( .A1(n3442), .A2(n3653), .A3(n7394), .Y(n7397) );
  NAND2X0_LVT U8708 ( .A1(n4005), .A2(n_T_427[1742]), .Y(n7396) );
  NAND2X0_LVT U8709 ( .A1(n3649), .A2(n_T_427[1614]), .Y(n7395) );
  NAND2X0_LVT U8710 ( .A1(n3625), .A2(ibuf_io_inst_0_bits_raw[15]), .Y(n7410)
         );
  NAND2X0_LVT U8711 ( .A1(n3716), .A2(n_T_427[1038]), .Y(n7409) );
  AND2X1_LVT U8712 ( .A1(n4050), .A2(n_T_427[15]), .Y(n7401) );
  AO22X1_LVT U8713 ( .A1(n4026), .A2(n_T_427[910]), .A3(n4019), .A4(
        n_T_427[655]), .Y(n7400) );
  AO22X1_LVT U8714 ( .A1(n3977), .A2(n_T_427[527]), .A3(n4029), .A4(
        n_T_427[846]), .Y(n7399) );
  AO22X1_LVT U8715 ( .A1(n4033), .A2(n_T_427[591]), .A3(n3984), .A4(
        n_T_427[207]), .Y(n7398) );
  NOR4X1_LVT U8716 ( .A1(n7401), .A2(n7400), .A3(n7399), .A4(n7398), .Y(n7407)
         );
  AO22X1_LVT U8717 ( .A1(n3969), .A2(n_T_427[399]), .A3(n3965), .A4(
        n_T_427[271]), .Y(n7405) );
  AO22X1_LVT U8718 ( .A1(n3973), .A2(n_T_427[143]), .A3(n4039), .A4(
        n_T_427[335]), .Y(n7404) );
  AO22X1_LVT U8719 ( .A1(n3980), .A2(n_T_427[782]), .A3(n4046), .A4(
        n_T_427[719]), .Y(n7403) );
  AO22X1_LVT U8720 ( .A1(n3961), .A2(n_T_427[463]), .A3(n4043), .A4(
        n_T_427[79]), .Y(n7402) );
  NOR4X1_LVT U8721 ( .A1(n7405), .A2(n7404), .A3(n7403), .A4(n7402), .Y(n7406)
         );
  AO21X1_LVT U8722 ( .A1(n7407), .A2(n7406), .A3(n3632), .Y(n7408) );
  NAND2X0_LVT U8723 ( .A1(n3641), .A2(n_T_427[1230]), .Y(n7411) );
  NAND2X0_LVT U8724 ( .A1(n3673), .A2(n_T_427[1102]), .Y(n7413) );
  NAND2X0_LVT U8725 ( .A1(n3756), .A2(n_T_427[974]), .Y(n7412) );
  NAND2X0_LVT U8726 ( .A1(n3627), .A2(n_T_427[1422]), .Y(n7414) );
  NAND2X0_LVT U8727 ( .A1(n3607), .A2(n_T_427[1358]), .Y(n7416) );
  NAND2X0_LVT U8728 ( .A1(n2985), .A2(n_T_427[1896]), .Y(n7415) );
  NAND2X0_LVT U8729 ( .A1(n2093), .A2(n_T_427[1295]), .Y(n7417) );
  OA21X1_LVT U8730 ( .A1(n3444), .A2(n3601), .A3(n7417), .Y(n7420) );
  NAND2X0_LVT U8731 ( .A1(n3744), .A2(n_T_427[1679]), .Y(n7419) );
  NAND2X0_LVT U8732 ( .A1(n4005), .A2(n_T_427[1743]), .Y(n7418) );
  NAND2X0_LVT U8733 ( .A1(n3619), .A2(n_T_427[1551]), .Y(n7421) );
  OA21X1_LVT U8734 ( .A1(n3664), .A2(n3312), .A3(n7421), .Y(n7424) );
  NAND2X0_LVT U8735 ( .A1(n3649), .A2(n_T_427[1615]), .Y(n7423) );
  NAND2X0_LVT U8736 ( .A1(n4006), .A2(n_T_427[1487]), .Y(n7422) );
  NAND2X0_LVT U8737 ( .A1(n3757), .A2(n_T_427[975]), .Y(n7425) );
  NAND2X0_LVT U8738 ( .A1(n3636), .A2(n_T_427[1231]), .Y(n7427) );
  NAND2X0_LVT U8739 ( .A1(n3667), .A2(n_T_427[1103]), .Y(n7426) );
  NAND2X0_LVT U8740 ( .A1(n2966), .A2(n_T_427[1423]), .Y(n7429) );
  NAND2X0_LVT U8741 ( .A1(n3608), .A2(n_T_427[1359]), .Y(n7428) );
  AND2X1_LVT U8742 ( .A1(n4050), .A2(n_T_427[16]), .Y(n7433) );
  AO22X1_LVT U8743 ( .A1(n4026), .A2(n_T_427[911]), .A3(n4019), .A4(
        n_T_427[656]), .Y(n7432) );
  AO22X1_LVT U8744 ( .A1(n3977), .A2(n_T_427[528]), .A3(n4029), .A4(
        n_T_427[847]), .Y(n7431) );
  AO22X1_LVT U8745 ( .A1(n4032), .A2(n_T_427[592]), .A3(n3984), .A4(
        n_T_427[208]), .Y(n7430) );
  NOR4X1_LVT U8746 ( .A1(n7433), .A2(n7432), .A3(n7431), .A4(n7430), .Y(n7439)
         );
  AO22X1_LVT U8747 ( .A1(n3969), .A2(n_T_427[400]), .A3(n3965), .A4(
        n_T_427[272]), .Y(n7437) );
  AO22X1_LVT U8748 ( .A1(n3974), .A2(n_T_427[144]), .A3(n4036), .A4(
        n_T_427[336]), .Y(n7436) );
  AO22X1_LVT U8749 ( .A1(n3980), .A2(n_T_427[783]), .A3(n4046), .A4(
        n_T_427[720]), .Y(n7435) );
  AO22X1_LVT U8750 ( .A1(n3961), .A2(n_T_427[464]), .A3(n2836), .A4(
        n_T_427[80]), .Y(n7434) );
  NOR4X1_LVT U8751 ( .A1(n7437), .A2(n7436), .A3(n7435), .A4(n7434), .Y(n7438)
         );
  AO21X1_LVT U8752 ( .A1(n7439), .A2(n7438), .A3(n2154), .Y(n7440) );
  NAND2X0_LVT U8753 ( .A1(n4000), .A2(n_T_427[1296]), .Y(n7443) );
  OA21X1_LVT U8754 ( .A1(n3142), .A2(n3747), .A3(n7443), .Y(n7446) );
  NAND2X0_LVT U8755 ( .A1(n3744), .A2(n_T_427[1680]), .Y(n7445) );
  NAND2X0_LVT U8756 ( .A1(n2092), .A2(n_T_427[1744]), .Y(n7444) );
  NAND2X0_LVT U8757 ( .A1(n3615), .A2(n_T_427[1552]), .Y(n7447) );
  OA21X1_LVT U8758 ( .A1(n4010), .A2(n3313), .A3(n7447), .Y(n7450) );
  NAND2X0_LVT U8759 ( .A1(n3652), .A2(n_T_427[1616]), .Y(n7449) );
  NAND2X0_LVT U8760 ( .A1(n4007), .A2(n_T_427[1488]), .Y(n7448) );
  NAND2X0_LVT U8761 ( .A1(n3758), .A2(n_T_427[976]), .Y(n7451) );
  OA21X1_LVT U8762 ( .A1(n3752), .A2(n3283), .A3(n7451), .Y(n7454) );
  NAND2X0_LVT U8763 ( .A1(n3639), .A2(n_T_427[1232]), .Y(n7453) );
  NAND2X0_LVT U8764 ( .A1(n3669), .A2(n_T_427[1104]), .Y(n7452) );
  NAND2X0_LVT U8765 ( .A1(n3992), .A2(n_T_427[1898]), .Y(n7455) );
  NAND2X0_LVT U8766 ( .A1(n3628), .A2(n_T_427[1424]), .Y(n7457) );
  NAND2X0_LVT U8767 ( .A1(n3605), .A2(n_T_427[1360]), .Y(n7456) );
  NAND2X0_LVT U8768 ( .A1(n3665), .A2(n4367), .Y(n7469) );
  AND2X1_LVT U8769 ( .A1(n4050), .A2(n_T_427[17]), .Y(n7461) );
  AO22X1_LVT U8770 ( .A1(n4025), .A2(n_T_427[912]), .A3(n4019), .A4(
        n_T_427[657]), .Y(n7460) );
  AO22X1_LVT U8771 ( .A1(n3977), .A2(n_T_427[529]), .A3(n4029), .A4(
        n_T_427[848]), .Y(n7459) );
  AO22X1_LVT U8772 ( .A1(n4033), .A2(n_T_427[593]), .A3(n3984), .A4(
        n_T_427[209]), .Y(n7458) );
  NOR4X1_LVT U8773 ( .A1(n7461), .A2(n7460), .A3(n7459), .A4(n7458), .Y(n7467)
         );
  AO22X1_LVT U8774 ( .A1(n3969), .A2(n_T_427[401]), .A3(n3965), .A4(
        n_T_427[273]), .Y(n7465) );
  AO22X1_LVT U8775 ( .A1(n3973), .A2(n_T_427[145]), .A3(n9040), .A4(
        n_T_427[337]), .Y(n7464) );
  AO22X1_LVT U8776 ( .A1(n3981), .A2(n_T_427[784]), .A3(n4046), .A4(
        n_T_427[721]), .Y(n7463) );
  AO22X1_LVT U8777 ( .A1(n3962), .A2(n_T_427[465]), .A3(n4042), .A4(
        n_T_427[81]), .Y(n7462) );
  NOR4X1_LVT U8778 ( .A1(n7465), .A2(n7464), .A3(n7463), .A4(n7462), .Y(n7466)
         );
  NAND2X0_LVT U8779 ( .A1(n3996), .A2(n_T_427[1297]), .Y(n7471) );
  OA21X1_LVT U8780 ( .A1(n3445), .A2(n3601), .A3(n7471), .Y(n7474) );
  NAND2X0_LVT U8781 ( .A1(n3744), .A2(n_T_427[1681]), .Y(n7473) );
  NAND2X0_LVT U8782 ( .A1(n2092), .A2(n_T_427[1745]), .Y(n7472) );
  NAND2X0_LVT U8783 ( .A1(n3620), .A2(n_T_427[1553]), .Y(n7475) );
  OA21X1_LVT U8784 ( .A1(n3663), .A2(n3314), .A3(n7475), .Y(n7478) );
  NAND2X0_LVT U8785 ( .A1(n3649), .A2(n_T_427[1617]), .Y(n7477) );
  NAND2X0_LVT U8786 ( .A1(n4007), .A2(n_T_427[1489]), .Y(n7476) );
  NAND2X0_LVT U8787 ( .A1(n3757), .A2(n_T_427[977]), .Y(n7479) );
  OA21X1_LVT U8788 ( .A1(n3752), .A2(n3315), .A3(n7479), .Y(n7482) );
  NAND2X0_LVT U8789 ( .A1(n3637), .A2(n_T_427[1233]), .Y(n7481) );
  NAND2X0_LVT U8790 ( .A1(n3673), .A2(n_T_427[1105]), .Y(n7480) );
  OA21X1_LVT U8791 ( .A1(n3988), .A2(n3316), .A3(n7483), .Y(n7486) );
  NAND2X0_LVT U8792 ( .A1(n3628), .A2(n_T_427[1425]), .Y(n7485) );
  NAND2X0_LVT U8793 ( .A1(n3602), .A2(n_T_427[1361]), .Y(n7484) );
  NAND2X0_LVT U8794 ( .A1(n4015), .A2(n4370), .Y(n7498) );
  AND2X1_LVT U8795 ( .A1(n4050), .A2(n_T_427[18]), .Y(n7490) );
  AO22X1_LVT U8796 ( .A1(n4026), .A2(n_T_427[913]), .A3(n4019), .A4(
        n_T_427[658]), .Y(n7489) );
  AO22X1_LVT U8797 ( .A1(n3977), .A2(n_T_427[530]), .A3(n4029), .A4(
        n_T_427[849]), .Y(n7488) );
  AO22X1_LVT U8798 ( .A1(n4033), .A2(n_T_427[594]), .A3(n3984), .A4(
        n_T_427[210]), .Y(n7487) );
  NOR4X1_LVT U8799 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .Y(n7496)
         );
  AO22X1_LVT U8800 ( .A1(n3969), .A2(n_T_427[402]), .A3(n3965), .A4(
        n_T_427[274]), .Y(n7494) );
  AO22X1_LVT U8801 ( .A1(n2858), .A2(n_T_427[146]), .A3(n4039), .A4(
        n_T_427[338]), .Y(n7493) );
  AO22X1_LVT U8802 ( .A1(n3981), .A2(n_T_427[785]), .A3(n4046), .A4(
        n_T_427[722]), .Y(n7492) );
  AO22X1_LVT U8803 ( .A1(n3962), .A2(n_T_427[466]), .A3(n2836), .A4(
        n_T_427[82]), .Y(n7491) );
  NOR4X1_LVT U8804 ( .A1(n7494), .A2(n7493), .A3(n7492), .A4(n7491), .Y(n7495)
         );
  AO21X1_LVT U8805 ( .A1(n7496), .A2(n7495), .A3(n2154), .Y(n7497) );
  NAND2X0_LVT U8806 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[18]), .Y(n7503) );
  NAND2X0_LVT U8807 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[18]), .Y(n7502)
         );
  NAND2X0_LVT U8808 ( .A1(n2497), .A2(n_T_628[18]), .Y(n7501) );
  NAND2X0_LVT U8809 ( .A1(n9066), .A2(n_T_918[18]), .Y(n7500) );
  NAND4X0_LVT U8810 ( .A1(n7503), .A2(n7502), .A3(n7501), .A4(n7500), .Y(
        io_fpu_fromint_data[18]) );
  NAND2X0_LVT U8811 ( .A1(n3997), .A2(n_T_427[1298]), .Y(n7504) );
  OA21X1_LVT U8812 ( .A1(n3446), .A2(n3751), .A3(n7504), .Y(n7507) );
  NAND2X0_LVT U8813 ( .A1(n3744), .A2(n_T_427[1682]), .Y(n7506) );
  NAND2X0_LVT U8814 ( .A1(n4002), .A2(n_T_427[1746]), .Y(n7505) );
  NAND2X0_LVT U8815 ( .A1(n3616), .A2(n_T_427[1554]), .Y(n7508) );
  OA21X1_LVT U8816 ( .A1(n4008), .A2(n3317), .A3(n7508), .Y(n7511) );
  NAND2X0_LVT U8817 ( .A1(n3648), .A2(n_T_427[1618]), .Y(n7510) );
  NAND2X0_LVT U8818 ( .A1(n4006), .A2(n_T_427[1490]), .Y(n7509) );
  NAND2X0_LVT U8819 ( .A1(n3712), .A2(n_T_427[978]), .Y(n7512) );
  OA21X1_LVT U8820 ( .A1(n3752), .A2(n3318), .A3(n7512), .Y(n7515) );
  NAND2X0_LVT U8821 ( .A1(n3640), .A2(n_T_427[1234]), .Y(n7514) );
  NAND2X0_LVT U8822 ( .A1(n3668), .A2(n_T_427[1106]), .Y(n7513) );
  NAND2X0_LVT U8823 ( .A1(n2882), .A2(n_T_427[1900]), .Y(n7516) );
  OA21X1_LVT U8824 ( .A1(n3987), .A2(n3319), .A3(n7516), .Y(n7519) );
  NAND2X0_LVT U8825 ( .A1(n3630), .A2(n_T_427[1426]), .Y(n7518) );
  NAND2X0_LVT U8826 ( .A1(n3608), .A2(n_T_427[1362]), .Y(n7517) );
  NAND2X0_LVT U8827 ( .A1(n3665), .A2(n4373), .Y(n7531) );
  AND2X1_LVT U8828 ( .A1(n4050), .A2(n_T_427[19]), .Y(n7523) );
  AO22X1_LVT U8829 ( .A1(n4025), .A2(n_T_427[914]), .A3(n4019), .A4(
        n_T_427[659]), .Y(n7522) );
  AO22X1_LVT U8830 ( .A1(n3978), .A2(n_T_427[531]), .A3(n4029), .A4(
        n_T_427[850]), .Y(n7521) );
  AO22X1_LVT U8831 ( .A1(n4033), .A2(n_T_427[595]), .A3(n3984), .A4(
        n_T_427[211]), .Y(n7520) );
  NOR4X1_LVT U8832 ( .A1(n7523), .A2(n7522), .A3(n7521), .A4(n7520), .Y(n7529)
         );
  AO22X1_LVT U8833 ( .A1(n3969), .A2(n_T_427[403]), .A3(n3965), .A4(
        n_T_427[275]), .Y(n7527) );
  AO22X1_LVT U8834 ( .A1(n3975), .A2(n_T_427[147]), .A3(n4038), .A4(
        n_T_427[339]), .Y(n7526) );
  AO22X1_LVT U8835 ( .A1(n3981), .A2(n_T_427[786]), .A3(n4046), .A4(
        n_T_427[723]), .Y(n7525) );
  AO22X1_LVT U8836 ( .A1(n3962), .A2(n_T_427[467]), .A3(n2837), .A4(
        n_T_427[83]), .Y(n7524) );
  NOR4X1_LVT U8837 ( .A1(n7527), .A2(n7526), .A3(n7525), .A4(n7524), .Y(n7528)
         );
  AO21X1_LVT U8838 ( .A1(n7529), .A2(n7528), .A3(n3632), .Y(n7530) );
  NAND2X0_LVT U8839 ( .A1(n3999), .A2(n_T_427[1299]), .Y(n7533) );
  OA21X1_LVT U8840 ( .A1(n3447), .A2(n3601), .A3(n7533), .Y(n7536) );
  NAND2X0_LVT U8841 ( .A1(n3744), .A2(n_T_427[1683]), .Y(n7535) );
  NAND2X0_LVT U8842 ( .A1(n4005), .A2(n_T_427[1747]), .Y(n7534) );
  NAND2X0_LVT U8843 ( .A1(n3617), .A2(n_T_427[1555]), .Y(n7537) );
  OA21X1_LVT U8844 ( .A1(n3663), .A2(n3320), .A3(n7537), .Y(n7540) );
  NAND2X0_LVT U8845 ( .A1(n3651), .A2(n_T_427[1619]), .Y(n7539) );
  NAND2X0_LVT U8846 ( .A1(n4007), .A2(n_T_427[1491]), .Y(n7538) );
  NAND2X0_LVT U8847 ( .A1(n3755), .A2(n_T_427[979]), .Y(n7541) );
  OA21X1_LVT U8848 ( .A1(n3752), .A2(n3321), .A3(n7541), .Y(n7544) );
  NAND2X0_LVT U8849 ( .A1(n3641), .A2(n_T_427[1235]), .Y(n7543) );
  NAND2X0_LVT U8850 ( .A1(n3670), .A2(n_T_427[1107]), .Y(n7542) );
  NAND2X0_LVT U8851 ( .A1(n3628), .A2(n_T_427[1427]), .Y(n7546) );
  NAND2X0_LVT U8852 ( .A1(n3604), .A2(n_T_427[1363]), .Y(n7545) );
  NAND2X0_LVT U8853 ( .A1(n2982), .A2(n4376), .Y(n7558) );
  AND2X1_LVT U8854 ( .A1(n4050), .A2(n_T_427[20]), .Y(n7550) );
  AO22X1_LVT U8855 ( .A1(n4025), .A2(n_T_427[915]), .A3(n4019), .A4(
        n_T_427[660]), .Y(n7549) );
  AO22X1_LVT U8856 ( .A1(n3978), .A2(n_T_427[532]), .A3(n4029), .A4(
        n_T_427[851]), .Y(n7548) );
  AO22X1_LVT U8857 ( .A1(n4033), .A2(n_T_427[596]), .A3(n3985), .A4(
        n_T_427[212]), .Y(n7547) );
  NOR4X1_LVT U8858 ( .A1(n7550), .A2(n7549), .A3(n7548), .A4(n7547), .Y(n7556)
         );
  AO22X1_LVT U8859 ( .A1(n3969), .A2(n_T_427[404]), .A3(n3965), .A4(
        n_T_427[276]), .Y(n7554) );
  AO22X1_LVT U8860 ( .A1(n2858), .A2(n_T_427[148]), .A3(n4038), .A4(
        n_T_427[340]), .Y(n7553) );
  AO22X1_LVT U8861 ( .A1(n3981), .A2(n_T_427[787]), .A3(n4046), .A4(
        n_T_427[724]), .Y(n7552) );
  AO22X1_LVT U8862 ( .A1(n3962), .A2(n_T_427[468]), .A3(n2836), .A4(
        n_T_427[84]), .Y(n7551) );
  NOR4X1_LVT U8863 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .Y(n7555)
         );
  AO21X1_LVT U8864 ( .A1(n7556), .A2(n7555), .A3(n3632), .Y(n7557) );
  NAND2X0_LVT U8865 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[20]), .Y(n7563) );
  NAND2X0_LVT U8866 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[20]), .Y(n7562)
         );
  NAND2X0_LVT U8867 ( .A1(n2497), .A2(n_T_628[20]), .Y(n7561) );
  NAND2X0_LVT U8868 ( .A1(n9066), .A2(n_T_918[20]), .Y(n7560) );
  NAND4X0_LVT U8869 ( .A1(n7563), .A2(n7562), .A3(n7561), .A4(n7560), .Y(
        io_fpu_fromint_data[20]) );
  NAND2X0_LVT U8870 ( .A1(n3996), .A2(n_T_427[1300]), .Y(n7564) );
  OA21X1_LVT U8871 ( .A1(n3391), .A2(n3601), .A3(n7564), .Y(n7567) );
  NAND2X0_LVT U8872 ( .A1(n3744), .A2(n_T_427[1684]), .Y(n7566) );
  NAND2X0_LVT U8873 ( .A1(n2091), .A2(n_T_427[1748]), .Y(n7565) );
  NAND2X0_LVT U8874 ( .A1(n3618), .A2(n_T_427[1556]), .Y(n7568) );
  OA21X1_LVT U8875 ( .A1(n3664), .A2(n3284), .A3(n7568), .Y(n7571) );
  NAND2X0_LVT U8876 ( .A1(n3648), .A2(n_T_427[1620]), .Y(n7570) );
  NAND2X0_LVT U8877 ( .A1(n4006), .A2(n_T_427[1492]), .Y(n7569) );
  NAND2X0_LVT U8878 ( .A1(n3758), .A2(n_T_427[980]), .Y(n7572) );
  OA21X1_LVT U8879 ( .A1(n3752), .A2(n3285), .A3(n7572), .Y(n7575) );
  NAND2X0_LVT U8880 ( .A1(n3639), .A2(n_T_427[1236]), .Y(n7574) );
  NAND2X0_LVT U8881 ( .A1(n3671), .A2(n_T_427[1108]), .Y(n7573) );
  NAND2X0_LVT U8882 ( .A1(n3992), .A2(n_T_427[1902]), .Y(n7576) );
  NAND2X0_LVT U8883 ( .A1(n3630), .A2(n_T_427[1428]), .Y(n7578) );
  NAND2X0_LVT U8884 ( .A1(n3602), .A2(n_T_427[1364]), .Y(n7577) );
  NAND2X0_LVT U8885 ( .A1(n3060), .A2(n4378), .Y(n7590) );
  AND2X1_LVT U8886 ( .A1(n4050), .A2(n_T_427[21]), .Y(n7582) );
  AO22X1_LVT U8887 ( .A1(n4025), .A2(n_T_427[916]), .A3(n4019), .A4(
        n_T_427[661]), .Y(n7581) );
  AO22X1_LVT U8888 ( .A1(n3978), .A2(n_T_427[533]), .A3(n4029), .A4(
        n_T_427[852]), .Y(n7580) );
  AO22X1_LVT U8889 ( .A1(n4033), .A2(n_T_427[597]), .A3(n3985), .A4(
        n_T_427[213]), .Y(n7579) );
  NOR4X1_LVT U8890 ( .A1(n7582), .A2(n7581), .A3(n7580), .A4(n7579), .Y(n7588)
         );
  AO22X1_LVT U8891 ( .A1(n3969), .A2(n_T_427[405]), .A3(n3965), .A4(
        n_T_427[277]), .Y(n7586) );
  AO22X1_LVT U8892 ( .A1(n2859), .A2(n_T_427[149]), .A3(n4038), .A4(
        n_T_427[341]), .Y(n7585) );
  AO22X1_LVT U8893 ( .A1(n3981), .A2(n_T_427[788]), .A3(n4046), .A4(
        n_T_427[725]), .Y(n7584) );
  AO22X1_LVT U8894 ( .A1(n3962), .A2(n_T_427[469]), .A3(n4041), .A4(
        n_T_427[85]), .Y(n7583) );
  NOR4X1_LVT U8895 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .Y(n7587)
         );
  NAND2X0_LVT U8896 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[21]), .Y(n7595) );
  NAND2X0_LVT U8897 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[21]), .Y(n7594)
         );
  NAND2X0_LVT U8898 ( .A1(n2497), .A2(n_T_628[21]), .Y(n7593) );
  NAND2X0_LVT U8899 ( .A1(n9066), .A2(n_T_918[21]), .Y(n7592) );
  NAND4X0_LVT U8900 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .Y(
        io_fpu_fromint_data[21]) );
  NAND2X0_LVT U8901 ( .A1(n2094), .A2(n_T_427[1301]), .Y(n7596) );
  OA21X1_LVT U8902 ( .A1(n3392), .A2(n3601), .A3(n7596), .Y(n7599) );
  NAND2X0_LVT U8903 ( .A1(n3744), .A2(n_T_427[1685]), .Y(n7598) );
  NAND2X0_LVT U8904 ( .A1(n4004), .A2(n_T_427[1749]), .Y(n7597) );
  NAND2X0_LVT U8905 ( .A1(n3619), .A2(n_T_427[1557]), .Y(n7600) );
  OA21X1_LVT U8906 ( .A1(n4010), .A2(n3286), .A3(n7600), .Y(n7603) );
  NAND2X0_LVT U8907 ( .A1(n3649), .A2(n_T_427[1621]), .Y(n7602) );
  NAND2X0_LVT U8908 ( .A1(n4006), .A2(n_T_427[1493]), .Y(n7601) );
  NAND2X0_LVT U8909 ( .A1(n3755), .A2(n_T_427[981]), .Y(n7604) );
  OA21X1_LVT U8910 ( .A1(n3752), .A2(n3287), .A3(n7604), .Y(n7607) );
  NAND2X0_LVT U8911 ( .A1(n_T_427[1237]), .A2(n3638), .Y(n7606) );
  NAND2X0_LVT U8912 ( .A1(n3670), .A2(n_T_427[1109]), .Y(n7605) );
  NAND2X0_LVT U8913 ( .A1(n2967), .A2(n_T_427[1429]), .Y(n7609) );
  NAND2X0_LVT U8914 ( .A1(n3609), .A2(n_T_427[1365]), .Y(n7608) );
  NAND2X0_LVT U8915 ( .A1(n3060), .A2(n4380), .Y(n7621) );
  AND2X1_LVT U8916 ( .A1(n4050), .A2(n_T_427[22]), .Y(n7613) );
  AO22X1_LVT U8917 ( .A1(n4025), .A2(n_T_427[917]), .A3(n4019), .A4(
        n_T_427[662]), .Y(n7612) );
  AO22X1_LVT U8918 ( .A1(n3978), .A2(n_T_427[534]), .A3(n4028), .A4(
        n_T_427[853]), .Y(n7611) );
  AO22X1_LVT U8919 ( .A1(n4033), .A2(n_T_427[598]), .A3(n3985), .A4(
        n_T_427[214]), .Y(n7610) );
  NOR4X1_LVT U8920 ( .A1(n7613), .A2(n7612), .A3(n7611), .A4(n7610), .Y(n7619)
         );
  AO22X1_LVT U8921 ( .A1(n3969), .A2(n_T_427[406]), .A3(n3965), .A4(
        n_T_427[278]), .Y(n7617) );
  AO22X1_LVT U8922 ( .A1(n2859), .A2(n_T_427[150]), .A3(n4038), .A4(
        n_T_427[342]), .Y(n7616) );
  AO22X1_LVT U8923 ( .A1(n3981), .A2(n_T_427[789]), .A3(n4046), .A4(
        n_T_427[726]), .Y(n7615) );
  AO22X1_LVT U8924 ( .A1(n3962), .A2(n_T_427[470]), .A3(n2837), .A4(
        n_T_427[86]), .Y(n7614) );
  NOR4X1_LVT U8925 ( .A1(n7617), .A2(n7616), .A3(n7615), .A4(n7614), .Y(n7618)
         );
  AO21X1_LVT U8926 ( .A1(n7619), .A2(n7618), .A3(n2155), .Y(n7620) );
  NAND2X0_LVT U8927 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[22]), .Y(n7626) );
  NAND2X0_LVT U8928 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[22]), .Y(n7625)
         );
  NAND2X0_LVT U8929 ( .A1(n2497), .A2(n_T_628[22]), .Y(n7624) );
  NAND2X0_LVT U8930 ( .A1(n9066), .A2(n_T_918[22]), .Y(n7623) );
  NAND4X0_LVT U8931 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .Y(
        io_fpu_fromint_data[22]) );
  NAND2X0_LVT U8932 ( .A1(n2094), .A2(n_T_427[1302]), .Y(n7627) );
  OA21X1_LVT U8933 ( .A1(n3448), .A2(n3751), .A3(n7627), .Y(n7630) );
  NAND2X0_LVT U8934 ( .A1(n3657), .A2(n_T_427[1686]), .Y(n7629) );
  NAND2X0_LVT U8935 ( .A1(n2092), .A2(n_T_427[1750]), .Y(n7628) );
  NAND2X0_LVT U8936 ( .A1(n3621), .A2(n_T_427[1558]), .Y(n7631) );
  OA21X1_LVT U8937 ( .A1(n2081), .A2(n3323), .A3(n7631), .Y(n7634) );
  NAND2X0_LVT U8938 ( .A1(n3642), .A2(n_T_427[1622]), .Y(n7633) );
  NAND2X0_LVT U8939 ( .A1(n4006), .A2(n_T_427[1494]), .Y(n7632) );
  NAND2X0_LVT U8940 ( .A1(n3760), .A2(n_T_427[982]), .Y(n7635) );
  OA21X1_LVT U8941 ( .A1(n3752), .A2(n3324), .A3(n7635), .Y(n7638) );
  NAND2X0_LVT U8942 ( .A1(n_T_427[1238]), .A2(n3638), .Y(n7637) );
  NAND2X0_LVT U8943 ( .A1(n3672), .A2(n_T_427[1110]), .Y(n7636) );
  NAND2X0_LVT U8944 ( .A1(n3991), .A2(n_T_427[1904]), .Y(n7639) );
  OA21X1_LVT U8945 ( .A1(n3989), .A2(n3325), .A3(n7639), .Y(n7642) );
  NAND2X0_LVT U8946 ( .A1(n3626), .A2(n_T_427[1430]), .Y(n7641) );
  NAND2X0_LVT U8947 ( .A1(n3602), .A2(n_T_427[1366]), .Y(n7640) );
  NAND2X0_LVT U8948 ( .A1(n4015), .A2(n4383), .Y(n7654) );
  AND2X1_LVT U8949 ( .A1(n4050), .A2(n_T_427[23]), .Y(n7646) );
  AO22X1_LVT U8950 ( .A1(n4025), .A2(n_T_427[918]), .A3(n4020), .A4(
        n_T_427[663]), .Y(n7645) );
  AO22X1_LVT U8951 ( .A1(n3978), .A2(n_T_427[535]), .A3(n4028), .A4(
        n_T_427[854]), .Y(n7644) );
  AO22X1_LVT U8952 ( .A1(n4033), .A2(n_T_427[599]), .A3(n3985), .A4(
        n_T_427[215]), .Y(n7643) );
  NOR4X1_LVT U8953 ( .A1(n7646), .A2(n7645), .A3(n7644), .A4(n7643), .Y(n7652)
         );
  AO22X1_LVT U8954 ( .A1(n3969), .A2(n_T_427[407]), .A3(n3965), .A4(
        n_T_427[279]), .Y(n7650) );
  AO22X1_LVT U8955 ( .A1(n3973), .A2(n_T_427[151]), .A3(n4038), .A4(
        n_T_427[343]), .Y(n7649) );
  AO22X1_LVT U8956 ( .A1(n3981), .A2(n_T_427[790]), .A3(n4046), .A4(
        n_T_427[727]), .Y(n7648) );
  AO22X1_LVT U8957 ( .A1(n3962), .A2(n_T_427[471]), .A3(n2837), .A4(
        n_T_427[87]), .Y(n7647) );
  NOR4X1_LVT U8958 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .Y(n7651)
         );
  AO21X1_LVT U8959 ( .A1(n7652), .A2(n7651), .A3(n2155), .Y(n7653) );
  NAND2X0_LVT U8960 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[23]), .Y(n7659) );
  NAND2X0_LVT U8961 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[23]), .Y(n7658)
         );
  NAND2X0_LVT U8962 ( .A1(n2497), .A2(n_T_628[23]), .Y(n7657) );
  NAND2X0_LVT U8963 ( .A1(n9066), .A2(n_T_918[23]), .Y(n7656) );
  NAND4X0_LVT U8964 ( .A1(n7659), .A2(n7658), .A3(n7657), .A4(n7656), .Y(
        io_fpu_fromint_data[23]) );
  NAND2X0_LVT U8965 ( .A1(n4000), .A2(n_T_427[1303]), .Y(n7660) );
  OA21X1_LVT U8966 ( .A1(n3449), .A2(n3747), .A3(n7660), .Y(n7663) );
  NAND2X0_LVT U8967 ( .A1(n2922), .A2(n_T_427[1687]), .Y(n7662) );
  NAND2X0_LVT U8968 ( .A1(n2091), .A2(n_T_427[1751]), .Y(n7661) );
  NAND3X0_LVT U8969 ( .A1(n7663), .A2(n7662), .A3(n7661), .Y(n7685) );
  NAND2X0_LVT U8970 ( .A1(n3620), .A2(n_T_427[1559]), .Y(n7664) );
  OA21X1_LVT U8971 ( .A1(n4010), .A2(n3326), .A3(n7664), .Y(n7667) );
  NAND2X0_LVT U8972 ( .A1(n3651), .A2(n_T_427[1623]), .Y(n7666) );
  NAND2X0_LVT U8973 ( .A1(n4006), .A2(n_T_427[1495]), .Y(n7665) );
  NAND3X0_LVT U8974 ( .A1(n7667), .A2(n7666), .A3(n7665), .Y(n7684) );
  NAND2X0_LVT U8975 ( .A1(n3759), .A2(n_T_427[983]), .Y(n7668) );
  NAND2X0_LVT U8976 ( .A1(n3640), .A2(n_T_427[1239]), .Y(n7670) );
  NAND2X0_LVT U8977 ( .A1(n3672), .A2(n_T_427[1111]), .Y(n7669) );
  NAND2X0_LVT U8978 ( .A1(n2882), .A2(n_T_427[1905]), .Y(n7671) );
  NAND2X0_LVT U8979 ( .A1(n3604), .A2(n_T_427[1367]), .Y(n7672) );
  NAND2X0_LVT U8980 ( .A1(n3665), .A2(n4386), .Y(n7682) );
  AND2X1_LVT U8981 ( .A1(n4050), .A2(n_T_427[24]), .Y(n7676) );
  AO22X1_LVT U8982 ( .A1(n4025), .A2(n_T_427[919]), .A3(n4020), .A4(
        n_T_427[664]), .Y(n7675) );
  AO22X1_LVT U8983 ( .A1(n3978), .A2(n_T_427[536]), .A3(n4028), .A4(
        n_T_427[855]), .Y(n7674) );
  AO22X1_LVT U8984 ( .A1(n4033), .A2(n_T_427[600]), .A3(n3985), .A4(
        n_T_427[216]), .Y(n7673) );
  AO22X1_LVT U8985 ( .A1(n3969), .A2(n_T_427[408]), .A3(n3966), .A4(
        n_T_427[280]), .Y(n7680) );
  AO22X1_LVT U8986 ( .A1(n3973), .A2(n_T_427[152]), .A3(n4038), .A4(
        n_T_427[344]), .Y(n7679) );
  AO22X1_LVT U8987 ( .A1(n3981), .A2(n_T_427[791]), .A3(n4047), .A4(
        n_T_427[728]), .Y(n7678) );
  AO22X1_LVT U8988 ( .A1(n3962), .A2(n_T_427[472]), .A3(n4042), .A4(
        n_T_427[88]), .Y(n7677) );
  NAND2X0_LVT U8989 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[24]), .Y(n7689) );
  NAND2X0_LVT U8990 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[24]), .Y(n7688)
         );
  NAND2X0_LVT U8991 ( .A1(n2497), .A2(n_T_628[24]), .Y(n7687) );
  NAND2X0_LVT U8992 ( .A1(n9066), .A2(n_T_918[24]), .Y(n7686) );
  NAND4X0_LVT U8993 ( .A1(n7689), .A2(n7688), .A3(n7687), .A4(n7686), .Y(
        io_fpu_fromint_data[24]) );
  NAND2X0_LVT U8994 ( .A1(n3999), .A2(n_T_427[1304]), .Y(n7690) );
  OA21X1_LVT U8995 ( .A1(n3393), .A2(n3747), .A3(n7690), .Y(n7693) );
  NAND2X0_LVT U8996 ( .A1(n3744), .A2(n_T_427[1688]), .Y(n7692) );
  NAND2X0_LVT U8997 ( .A1(n2091), .A2(n_T_427[1752]), .Y(n7691) );
  NAND2X0_LVT U8998 ( .A1(n3621), .A2(n_T_427[1560]), .Y(n7694) );
  OA21X1_LVT U8999 ( .A1(n4009), .A2(n3288), .A3(n7694), .Y(n7697) );
  NAND2X0_LVT U9000 ( .A1(n3643), .A2(n_T_427[1624]), .Y(n7696) );
  NAND2X0_LVT U9001 ( .A1(n4007), .A2(n_T_427[1496]), .Y(n7695) );
  NAND2X0_LVT U9002 ( .A1(n3758), .A2(n_T_427[984]), .Y(n7698) );
  OA21X1_LVT U9003 ( .A1(n3752), .A2(n3289), .A3(n7698), .Y(n7701) );
  NAND2X0_LVT U9004 ( .A1(n3636), .A2(n_T_427[1240]), .Y(n7700) );
  NAND2X0_LVT U9005 ( .A1(n3674), .A2(n_T_427[1112]), .Y(n7699) );
  NAND2X0_LVT U9006 ( .A1(n2998), .A2(n_T_427[1906]), .Y(n7702) );
  OA21X1_LVT U9007 ( .A1(n3989), .A2(n3372), .A3(n7702), .Y(n7705) );
  NAND2X0_LVT U9008 ( .A1(n3626), .A2(n_T_427[1432]), .Y(n7704) );
  NAND2X0_LVT U9009 ( .A1(n3603), .A2(n_T_427[1368]), .Y(n7703) );
  NAND2X0_LVT U9010 ( .A1(n3060), .A2(n4388), .Y(n7717) );
  AND2X1_LVT U9011 ( .A1(n4051), .A2(n_T_427[25]), .Y(n7709) );
  AO22X1_LVT U9012 ( .A1(n4025), .A2(n_T_427[920]), .A3(n4020), .A4(
        n_T_427[665]), .Y(n7708) );
  AO22X1_LVT U9013 ( .A1(n3976), .A2(n_T_427[537]), .A3(n4028), .A4(
        n_T_427[856]), .Y(n7707) );
  AO22X1_LVT U9014 ( .A1(n4033), .A2(n_T_427[601]), .A3(n3985), .A4(
        n_T_427[217]), .Y(n7706) );
  NOR4X1_LVT U9015 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .Y(n7715)
         );
  AO22X1_LVT U9016 ( .A1(n3970), .A2(n_T_427[409]), .A3(n3966), .A4(
        n_T_427[281]), .Y(n7713) );
  AO22X1_LVT U9017 ( .A1(n2858), .A2(n_T_427[153]), .A3(n4038), .A4(
        n_T_427[345]), .Y(n7712) );
  AO22X1_LVT U9018 ( .A1(n3981), .A2(n_T_427[792]), .A3(n4047), .A4(
        n_T_427[729]), .Y(n7711) );
  AO22X1_LVT U9019 ( .A1(n3962), .A2(n_T_427[473]), .A3(n4044), .A4(
        n_T_427[89]), .Y(n7710) );
  NOR4X1_LVT U9020 ( .A1(n7713), .A2(n7712), .A3(n7711), .A4(n7710), .Y(n7714)
         );
  AO21X1_LVT U9021 ( .A1(n7715), .A2(n7714), .A3(n2645), .Y(n7716) );
  NAND2X0_LVT U9022 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[25]), .Y(n7722) );
  NAND2X0_LVT U9023 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[25]), .Y(n7721)
         );
  NAND2X0_LVT U9024 ( .A1(n2497), .A2(n_T_628[25]), .Y(n7720) );
  NAND2X0_LVT U9025 ( .A1(n9066), .A2(n_T_918[25]), .Y(n7719) );
  NAND4X0_LVT U9026 ( .A1(n7722), .A2(n7721), .A3(n7720), .A4(n7719), .Y(
        io_fpu_fromint_data[25]) );
  NAND2X0_LVT U9027 ( .A1(n3997), .A2(n_T_427[1305]), .Y(n7723) );
  OA21X1_LVT U9028 ( .A1(n3394), .A2(n3747), .A3(n7723), .Y(n7726) );
  NAND2X0_LVT U9029 ( .A1(n3744), .A2(n_T_427[1689]), .Y(n7725) );
  NAND2X0_LVT U9030 ( .A1(n4001), .A2(n_T_427[1753]), .Y(n7724) );
  NAND2X0_LVT U9031 ( .A1(n3621), .A2(n_T_427[1561]), .Y(n7727) );
  OA21X1_LVT U9032 ( .A1(n2081), .A2(n3290), .A3(n7727), .Y(n7730) );
  NAND2X0_LVT U9033 ( .A1(n3652), .A2(n_T_427[1625]), .Y(n7729) );
  NAND2X0_LVT U9034 ( .A1(n4006), .A2(n_T_427[1497]), .Y(n7728) );
  NAND2X0_LVT U9035 ( .A1(n3756), .A2(n_T_427[985]), .Y(n7731) );
  OA21X1_LVT U9036 ( .A1(n3752), .A2(n3291), .A3(n7731), .Y(n7734) );
  NAND2X0_LVT U9037 ( .A1(n3637), .A2(n_T_427[1241]), .Y(n7733) );
  NAND2X0_LVT U9038 ( .A1(n3675), .A2(n_T_427[1113]), .Y(n7732) );
  NAND2X0_LVT U9039 ( .A1(n2998), .A2(n_T_427[1907]), .Y(n7735) );
  OA21X1_LVT U9040 ( .A1(n3987), .A2(n3373), .A3(n7735), .Y(n7738) );
  NAND2X0_LVT U9041 ( .A1(n3628), .A2(n_T_427[1433]), .Y(n7737) );
  NAND2X0_LVT U9042 ( .A1(n3603), .A2(n_T_427[1369]), .Y(n7736) );
  NAND2X0_LVT U9043 ( .A1(n2982), .A2(n4390), .Y(n7750) );
  AND2X1_LVT U9044 ( .A1(n4051), .A2(n_T_427[26]), .Y(n7742) );
  AO22X1_LVT U9045 ( .A1(n4025), .A2(n_T_427[921]), .A3(n4020), .A4(
        n_T_427[666]), .Y(n7741) );
  AO22X1_LVT U9046 ( .A1(n3978), .A2(n_T_427[538]), .A3(n4028), .A4(
        n_T_427[857]), .Y(n7740) );
  AO22X1_LVT U9047 ( .A1(n4033), .A2(n_T_427[602]), .A3(n3985), .A4(
        n_T_427[218]), .Y(n7739) );
  NOR4X1_LVT U9048 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .Y(n7748)
         );
  AO22X1_LVT U9049 ( .A1(n3970), .A2(n_T_427[410]), .A3(n3966), .A4(
        n_T_427[282]), .Y(n7746) );
  AO22X1_LVT U9050 ( .A1(n3975), .A2(n_T_427[154]), .A3(n4038), .A4(
        n_T_427[346]), .Y(n7745) );
  AO22X1_LVT U9051 ( .A1(n3981), .A2(n_T_427[793]), .A3(n4047), .A4(
        n_T_427[730]), .Y(n7744) );
  AO22X1_LVT U9052 ( .A1(n3962), .A2(n_T_427[474]), .A3(n4041), .A4(
        n_T_427[90]), .Y(n7743) );
  NOR4X1_LVT U9053 ( .A1(n7746), .A2(n7745), .A3(n7744), .A4(n7743), .Y(n7747)
         );
  NAND2X0_LVT U9054 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[26]), .Y(n7755) );
  NAND2X0_LVT U9055 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[26]), .Y(n7754)
         );
  NAND2X0_LVT U9056 ( .A1(n2497), .A2(n_T_628[26]), .Y(n7753) );
  NAND2X0_LVT U9057 ( .A1(n9066), .A2(n_T_918[26]), .Y(n7752) );
  NAND4X0_LVT U9058 ( .A1(n7755), .A2(n7754), .A3(n7753), .A4(n7752), .Y(
        io_fpu_fromint_data[26]) );
  NAND2X0_LVT U9059 ( .A1(n3999), .A2(n_T_427[1306]), .Y(n7756) );
  OA21X1_LVT U9060 ( .A1(n3450), .A2(n3751), .A3(n7756), .Y(n7759) );
  NAND2X0_LVT U9061 ( .A1(n3744), .A2(n_T_427[1690]), .Y(n7758) );
  NAND2X0_LVT U9062 ( .A1(n4002), .A2(n_T_427[1754]), .Y(n7757) );
  NAND2X0_LVT U9063 ( .A1(n3618), .A2(n_T_427[1562]), .Y(n7760) );
  OA21X1_LVT U9064 ( .A1(n2081), .A2(n3328), .A3(n7760), .Y(n7762) );
  NAND2X0_LVT U9065 ( .A1(n4007), .A2(n_T_427[1498]), .Y(n7761) );
  NAND2X0_LVT U9066 ( .A1(n3757), .A2(n_T_427[986]), .Y(n7763) );
  OA21X1_LVT U9067 ( .A1(n3752), .A2(n3329), .A3(n7763), .Y(n7766) );
  NAND2X0_LVT U9068 ( .A1(n3636), .A2(n_T_427[1242]), .Y(n7765) );
  NAND2X0_LVT U9069 ( .A1(n3672), .A2(n_T_427[1114]), .Y(n7764) );
  NAND2X0_LVT U9070 ( .A1(n2985), .A2(n_T_427[1908]), .Y(n7767) );
  OA21X1_LVT U9071 ( .A1(n2120), .A2(n3330), .A3(n7767), .Y(n7770) );
  NAND2X0_LVT U9072 ( .A1(n2966), .A2(n_T_427[1434]), .Y(n7769) );
  NAND2X0_LVT U9073 ( .A1(n3607), .A2(n_T_427[1370]), .Y(n7768) );
  NAND2X0_LVT U9074 ( .A1(n4015), .A2(n4393), .Y(n7782) );
  AND2X1_LVT U9075 ( .A1(n4051), .A2(n_T_427[27]), .Y(n7774) );
  AO22X1_LVT U9076 ( .A1(n4025), .A2(n_T_427[922]), .A3(n4020), .A4(
        n_T_427[667]), .Y(n7773) );
  AO22X1_LVT U9077 ( .A1(n3978), .A2(n_T_427[539]), .A3(n4028), .A4(
        n_T_427[858]), .Y(n7772) );
  AO22X1_LVT U9078 ( .A1(n4033), .A2(n_T_427[603]), .A3(n3985), .A4(
        n_T_427[219]), .Y(n7771) );
  NOR4X1_LVT U9079 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .Y(n7780)
         );
  AO22X1_LVT U9080 ( .A1(n3970), .A2(n_T_427[411]), .A3(n3966), .A4(
        n_T_427[283]), .Y(n7778) );
  AO22X1_LVT U9081 ( .A1(n3973), .A2(n_T_427[155]), .A3(n4038), .A4(
        n_T_427[347]), .Y(n7777) );
  AO22X1_LVT U9082 ( .A1(n3981), .A2(n_T_427[794]), .A3(n4047), .A4(
        n_T_427[731]), .Y(n7776) );
  AO22X1_LVT U9083 ( .A1(n3962), .A2(n_T_427[475]), .A3(n2836), .A4(
        n_T_427[91]), .Y(n7775) );
  NOR4X1_LVT U9084 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .Y(n7779)
         );
  NAND2X0_LVT U9085 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[27]), .Y(n7787) );
  NAND2X0_LVT U9086 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[27]), .Y(n7786)
         );
  NAND2X0_LVT U9087 ( .A1(n2497), .A2(n_T_628[27]), .Y(n7785) );
  NAND2X0_LVT U9088 ( .A1(n9066), .A2(n_T_918[27]), .Y(n7784) );
  NAND4X0_LVT U9089 ( .A1(n7787), .A2(n7786), .A3(n7785), .A4(n7784), .Y(
        io_fpu_fromint_data[27]) );
  NAND2X0_LVT U9090 ( .A1(n2093), .A2(n_T_427[1307]), .Y(n7788) );
  OA21X1_LVT U9091 ( .A1(n3395), .A2(n3601), .A3(n7788), .Y(n7791) );
  NAND2X0_LVT U9092 ( .A1(n3744), .A2(n_T_427[1691]), .Y(n7790) );
  NAND2X0_LVT U9093 ( .A1(n4004), .A2(n_T_427[1755]), .Y(n7789) );
  NAND2X0_LVT U9094 ( .A1(n3615), .A2(n_T_427[1563]), .Y(n7792) );
  OA21X1_LVT U9095 ( .A1(n4008), .A2(n3292), .A3(n7792), .Y(n7794) );
  NAND2X0_LVT U9096 ( .A1(n4007), .A2(n_T_427[1499]), .Y(n7793) );
  NAND2X0_LVT U9097 ( .A1(n3760), .A2(n_T_427[987]), .Y(n7795) );
  OA21X1_LVT U9098 ( .A1(n4012), .A2(n3293), .A3(n7795), .Y(n7798) );
  NAND2X0_LVT U9099 ( .A1(n3639), .A2(n_T_427[1243]), .Y(n7797) );
  NAND2X0_LVT U9100 ( .A1(n3672), .A2(n_T_427[1115]), .Y(n7796) );
  NAND2X0_LVT U9101 ( .A1(n3992), .A2(n_T_427[1909]), .Y(n7799) );
  OA21X1_LVT U9102 ( .A1(n3767), .A2(n3374), .A3(n7799), .Y(n7802) );
  NAND2X0_LVT U9103 ( .A1(n3630), .A2(n_T_427[1435]), .Y(n7801) );
  NAND2X0_LVT U9104 ( .A1(n3604), .A2(n_T_427[1371]), .Y(n7800) );
  AND2X1_LVT U9105 ( .A1(n4051), .A2(n_T_427[28]), .Y(n7806) );
  AO22X1_LVT U9106 ( .A1(n4025), .A2(n_T_427[923]), .A3(n4020), .A4(
        n_T_427[668]), .Y(n7805) );
  AO22X1_LVT U9107 ( .A1(n3978), .A2(n_T_427[540]), .A3(n4028), .A4(
        n_T_427[859]), .Y(n7804) );
  AO22X1_LVT U9108 ( .A1(n4033), .A2(n_T_427[604]), .A3(n3985), .A4(
        n_T_427[220]), .Y(n7803) );
  NOR4X1_LVT U9109 ( .A1(n7806), .A2(n7805), .A3(n7804), .A4(n7803), .Y(n7812)
         );
  AO22X1_LVT U9110 ( .A1(n3970), .A2(n_T_427[412]), .A3(n3966), .A4(
        n_T_427[284]), .Y(n7810) );
  AO22X1_LVT U9111 ( .A1(n3974), .A2(n_T_427[156]), .A3(n4038), .A4(
        n_T_427[348]), .Y(n7809) );
  AO22X1_LVT U9112 ( .A1(n3981), .A2(n_T_427[795]), .A3(n4047), .A4(
        n_T_427[732]), .Y(n7808) );
  AO22X1_LVT U9113 ( .A1(n3962), .A2(n_T_427[476]), .A3(n4043), .A4(
        n_T_427[92]), .Y(n7807) );
  NOR4X1_LVT U9114 ( .A1(n7810), .A2(n7809), .A3(n7808), .A4(n7807), .Y(n7811)
         );
  NAND2X0_LVT U9115 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[28]), .Y(n7819) );
  NAND2X0_LVT U9116 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[28]), .Y(n7818)
         );
  NAND2X0_LVT U9117 ( .A1(n2493), .A2(n_T_628[28]), .Y(n7817) );
  NAND2X0_LVT U9118 ( .A1(n9066), .A2(n_T_918[28]), .Y(n7816) );
  NAND4X0_LVT U9119 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .Y(
        io_fpu_fromint_data[28]) );
  NAND2X0_LVT U9120 ( .A1(n4000), .A2(n_T_427[1308]), .Y(n7820) );
  OA21X1_LVT U9121 ( .A1(n3396), .A2(n3601), .A3(n7820), .Y(n7823) );
  NAND2X0_LVT U9122 ( .A1(n3744), .A2(n_T_427[1692]), .Y(n7822) );
  NAND2X0_LVT U9123 ( .A1(n4003), .A2(n_T_427[1756]), .Y(n7821) );
  NAND2X0_LVT U9124 ( .A1(n3616), .A2(n_T_427[1564]), .Y(n7824) );
  OA21X1_LVT U9125 ( .A1(n4008), .A2(n3294), .A3(n7824), .Y(n7827) );
  NAND2X0_LVT U9126 ( .A1(n3642), .A2(n_T_427[1628]), .Y(n7826) );
  NAND2X0_LVT U9127 ( .A1(n4007), .A2(n_T_427[1500]), .Y(n7825) );
  NAND2X0_LVT U9128 ( .A1(n3755), .A2(n_T_427[988]), .Y(n7828) );
  OA21X1_LVT U9129 ( .A1(n4013), .A2(n3295), .A3(n7828), .Y(n7831) );
  NAND2X0_LVT U9130 ( .A1(n3640), .A2(n_T_427[1244]), .Y(n7830) );
  NAND2X0_LVT U9131 ( .A1(n3675), .A2(n_T_427[1116]), .Y(n7829) );
  NAND2X0_LVT U9132 ( .A1(n2986), .A2(n_T_427[1910]), .Y(n7832) );
  OA21X1_LVT U9133 ( .A1(n2120), .A2(n3375), .A3(n7832), .Y(n7835) );
  NAND2X0_LVT U9134 ( .A1(n2967), .A2(n_T_427[1436]), .Y(n7834) );
  NAND2X0_LVT U9135 ( .A1(n3603), .A2(n_T_427[1372]), .Y(n7833) );
  AND2X1_LVT U9136 ( .A1(n4051), .A2(n_T_427[29]), .Y(n7839) );
  AO22X1_LVT U9137 ( .A1(n4025), .A2(n_T_427[924]), .A3(n4020), .A4(
        n_T_427[669]), .Y(n7838) );
  AO22X1_LVT U9138 ( .A1(n3978), .A2(n_T_427[541]), .A3(n4028), .A4(
        n_T_427[860]), .Y(n7837) );
  AO22X1_LVT U9139 ( .A1(n4034), .A2(n_T_427[605]), .A3(n3985), .A4(
        n_T_427[221]), .Y(n7836) );
  NOR4X1_LVT U9140 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .Y(n7845)
         );
  AO22X1_LVT U9141 ( .A1(n3970), .A2(n_T_427[413]), .A3(n3966), .A4(
        n_T_427[285]), .Y(n7843) );
  AO22X1_LVT U9142 ( .A1(n3974), .A2(n_T_427[157]), .A3(n4038), .A4(
        n_T_427[349]), .Y(n7842) );
  AO22X1_LVT U9143 ( .A1(n3981), .A2(n_T_427[796]), .A3(n4047), .A4(
        n_T_427[733]), .Y(n7841) );
  AO22X1_LVT U9144 ( .A1(n3962), .A2(n_T_427[477]), .A3(n4041), .A4(
        n_T_427[93]), .Y(n7840) );
  NOR4X1_LVT U9145 ( .A1(n7843), .A2(n7842), .A3(n7841), .A4(n7840), .Y(n7844)
         );
  AO21X1_LVT U9146 ( .A1(n7845), .A2(n7844), .A3(n3656), .Y(n7846) );
  NAND2X0_LVT U9147 ( .A1(n3998), .A2(n_T_427[1309]), .Y(n7849) );
  OA21X1_LVT U9148 ( .A1(n3451), .A2(n3601), .A3(n7849), .Y(n7852) );
  NAND2X0_LVT U9149 ( .A1(n3744), .A2(n_T_427[1693]), .Y(n7851) );
  NAND2X0_LVT U9150 ( .A1(n2091), .A2(n_T_427[1757]), .Y(n7850) );
  NAND2X0_LVT U9151 ( .A1(n3617), .A2(n_T_427[1565]), .Y(n7853) );
  OA21X1_LVT U9152 ( .A1(n4010), .A2(n3331), .A3(n7853), .Y(n7856) );
  NAND2X0_LVT U9153 ( .A1(n3651), .A2(n_T_427[1629]), .Y(n7855) );
  NAND2X0_LVT U9154 ( .A1(n3769), .A2(n_T_427[1501]), .Y(n7854) );
  NAND2X0_LVT U9155 ( .A1(n_T_427[1245]), .A2(n3638), .Y(n7858) );
  NAND2X0_LVT U9156 ( .A1(n3671), .A2(n_T_427[1117]), .Y(n7857) );
  NAND2X0_LVT U9157 ( .A1(n3992), .A2(n_T_427[1911]), .Y(n7860) );
  NAND2X0_LVT U9158 ( .A1(n3627), .A2(n_T_427[1437]), .Y(n7862) );
  NAND2X0_LVT U9159 ( .A1(n3605), .A2(n_T_427[1373]), .Y(n7861) );
  AND2X1_LVT U9160 ( .A1(n4051), .A2(n_T_427[30]), .Y(n7866) );
  AO22X1_LVT U9161 ( .A1(n4024), .A2(n_T_427[925]), .A3(n4020), .A4(
        n_T_427[670]), .Y(n7865) );
  AO22X1_LVT U9162 ( .A1(n3978), .A2(n_T_427[542]), .A3(n4028), .A4(
        n_T_427[861]), .Y(n7864) );
  AO22X1_LVT U9163 ( .A1(n4034), .A2(n_T_427[606]), .A3(n3985), .A4(
        n_T_427[222]), .Y(n7863) );
  NOR4X1_LVT U9164 ( .A1(n7866), .A2(n7865), .A3(n7864), .A4(n7863), .Y(n7872)
         );
  AO22X1_LVT U9165 ( .A1(n3970), .A2(n_T_427[414]), .A3(n3966), .A4(
        n_T_427[286]), .Y(n7870) );
  AO22X1_LVT U9166 ( .A1(n3974), .A2(n_T_427[158]), .A3(n4037), .A4(
        n_T_427[350]), .Y(n7869) );
  AO22X1_LVT U9167 ( .A1(n3982), .A2(n_T_427[797]), .A3(n4047), .A4(
        n_T_427[734]), .Y(n7868) );
  AO22X1_LVT U9168 ( .A1(n3963), .A2(n_T_427[478]), .A3(n4044), .A4(
        n_T_427[94]), .Y(n7867) );
  NOR4X1_LVT U9169 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .Y(n7871)
         );
  NAND2X0_LVT U9170 ( .A1(n2094), .A2(n_T_427[1310]), .Y(n7876) );
  OA21X1_LVT U9171 ( .A1(n3397), .A2(n3751), .A3(n7876), .Y(n7879) );
  NAND2X0_LVT U9172 ( .A1(n3689), .A2(n_T_427[1694]), .Y(n7878) );
  NAND2X0_LVT U9173 ( .A1(n4001), .A2(n_T_427[1758]), .Y(n7877) );
  NAND2X0_LVT U9174 ( .A1(n3618), .A2(n_T_427[1566]), .Y(n7880) );
  OA21X1_LVT U9175 ( .A1(n3664), .A2(n3296), .A3(n7880), .Y(n7882) );
  NAND2X0_LVT U9176 ( .A1(n4007), .A2(n_T_427[1502]), .Y(n7881) );
  NAND2X0_LVT U9177 ( .A1(n3759), .A2(n_T_427[990]), .Y(n7883) );
  OA21X1_LVT U9178 ( .A1(n4011), .A2(n3297), .A3(n7883), .Y(n7886) );
  NAND2X0_LVT U9179 ( .A1(n3641), .A2(n_T_427[1246]), .Y(n7885) );
  NAND2X0_LVT U9180 ( .A1(n3672), .A2(n_T_427[1118]), .Y(n7884) );
  NAND2X0_LVT U9181 ( .A1(n2985), .A2(n_T_427[1912]), .Y(n7887) );
  OA21X1_LVT U9182 ( .A1(n3767), .A2(n3376), .A3(n7887), .Y(n7890) );
  NAND2X0_LVT U9183 ( .A1(n3630), .A2(n_T_427[1438]), .Y(n7889) );
  NAND2X0_LVT U9184 ( .A1(n_T_427[1374]), .A2(n3611), .Y(n7888) );
  NAND2X0_LVT U9185 ( .A1(n4015), .A2(n4403), .Y(n7902) );
  AND2X1_LVT U9186 ( .A1(n4051), .A2(n_T_427[31]), .Y(n7894) );
  AO22X1_LVT U9187 ( .A1(n4024), .A2(n_T_427[926]), .A3(n4020), .A4(
        n_T_427[671]), .Y(n7893) );
  AO22X1_LVT U9188 ( .A1(n3978), .A2(n_T_427[543]), .A3(n4028), .A4(
        n_T_427[862]), .Y(n7892) );
  AO22X1_LVT U9189 ( .A1(n4034), .A2(n_T_427[607]), .A3(n3985), .A4(
        n_T_427[223]), .Y(n7891) );
  NOR4X1_LVT U9190 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .Y(n7900)
         );
  AO22X1_LVT U9191 ( .A1(n3970), .A2(n_T_427[415]), .A3(n3966), .A4(
        n_T_427[287]), .Y(n7898) );
  AO22X1_LVT U9192 ( .A1(n2858), .A2(n_T_427[159]), .A3(n4037), .A4(
        n_T_427[351]), .Y(n7897) );
  AO22X1_LVT U9193 ( .A1(n3982), .A2(n_T_427[798]), .A3(n4047), .A4(
        n_T_427[735]), .Y(n7896) );
  AO22X1_LVT U9194 ( .A1(n3963), .A2(n_T_427[479]), .A3(n4043), .A4(
        n_T_427[95]), .Y(n7895) );
  NOR4X1_LVT U9195 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .Y(n7899)
         );
  AO21X1_LVT U9196 ( .A1(n7900), .A2(n7899), .A3(n3632), .Y(n7901) );
  AO22X1_LVT U9197 ( .A1(n2497), .A2(n_T_628[31]), .A3(n9064), .A4(
        io_fpu_dmem_resp_data[31]), .Y(n7905) );
  AO22X1_LVT U9198 ( .A1(n9066), .A2(n_T_918[31]), .A3(n9065), .A4(
        io_imem_sfence_bits_addr[31]), .Y(n7904) );
  NAND2X0_LVT U9199 ( .A1(n3757), .A2(n_T_427[991]), .Y(n7906) );
  OA21X1_LVT U9200 ( .A1(n4012), .A2(n3333), .A3(n7906), .Y(n7909) );
  NAND2X0_LVT U9201 ( .A1(n3637), .A2(n_T_427[1247]), .Y(n7908) );
  NAND2X0_LVT U9202 ( .A1(n3672), .A2(n_T_427[1119]), .Y(n7907) );
  AND2X1_LVT U9203 ( .A1(n3976), .A2(n8105), .Y(n9035) );
  NAND2X0_LVT U9204 ( .A1(n3786), .A2(n_T_427[544]), .Y(n7921) );
  NAND2X0_LVT U9205 ( .A1(n3060), .A2(n4406), .Y(n7920) );
  AO22X1_LVT U9206 ( .A1(n4024), .A2(n_T_427[927]), .A3(n4041), .A4(
        n_T_427[96]), .Y(n7917) );
  AO22X1_LVT U9207 ( .A1(n3970), .A2(n_T_427[416]), .A3(n4037), .A4(
        n_T_427[352]), .Y(n7916) );
  AOI22X1_LVT U9208 ( .A1(n4035), .A2(n_T_427[608]), .A3(n4027), .A4(
        n_T_427[863]), .Y(n7914) );
  AOI22X1_LVT U9209 ( .A1(n2858), .A2(n_T_427[160]), .A3(n4051), .A4(
        n_T_427[32]), .Y(n7913) );
  AOI22X1_LVT U9210 ( .A1(n4022), .A2(n_T_427[672]), .A3(n3983), .A4(
        n_T_427[224]), .Y(n7912) );
  NAND3X0_LVT U9211 ( .A1(n7914), .A2(n7913), .A3(n7912), .Y(n7915) );
  OR3X1_LVT U9212 ( .A1(n7917), .A2(n7916), .A3(n7915), .Y(n7918) );
  NAND2X0_LVT U9213 ( .A1(n4053), .A2(n7918), .Y(n7919) );
  AND3X1_LVT U9214 ( .A1(n7921), .A2(n7920), .A3(n7919), .Y(n7924) );
  AND2X1_LVT U9215 ( .A1(n3964), .A2(n8105), .Y(n9053) );
  NAND2X0_LVT U9216 ( .A1(n3789), .A2(n_T_427[288]), .Y(n7922) );
  NAND2X0_LVT U9217 ( .A1(n3689), .A2(n_T_427[1695]), .Y(n7925) );
  OA21X1_LVT U9218 ( .A1(n3143), .A2(n3751), .A3(n7925), .Y(n7928) );
  NAND2X0_LVT U9219 ( .A1(n4000), .A2(n_T_427[1311]), .Y(n7927) );
  NAND2X0_LVT U9220 ( .A1(n2091), .A2(n_T_427[1759]), .Y(n7926) );
  NAND2X0_LVT U9221 ( .A1(n3769), .A2(n_T_427[1503]), .Y(n7929) );
  OA21X1_LVT U9222 ( .A1(n2081), .A2(n3334), .A3(n7929), .Y(n7932) );
  NAND2X0_LVT U9223 ( .A1(n3616), .A2(n_T_427[1567]), .Y(n7931) );
  NAND2X0_LVT U9224 ( .A1(n3652), .A2(n_T_427[1631]), .Y(n7930) );
  NAND2X0_LVT U9225 ( .A1(n9056), .A2(n_T_427[799]), .Y(n7933) );
  OA21X1_LVT U9226 ( .A1(n3398), .A2(n3691), .A3(n7933), .Y(n7938) );
  NAND2X0_LVT U9227 ( .A1(n3629), .A2(n_T_427[1439]), .Y(n7934) );
  NAND2X0_LVT U9228 ( .A1(n3603), .A2(n_T_427[1375]), .Y(n7935) );
  NAND2X0_LVT U9229 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[32]), .Y(n7942) );
  NAND2X0_LVT U9230 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[32]), .Y(n7941)
         );
  NAND2X0_LVT U9231 ( .A1(n2497), .A2(n_T_628[32]), .Y(n7940) );
  NAND2X0_LVT U9232 ( .A1(n9066), .A2(n_T_918[32]), .Y(n7939) );
  NAND4X0_LVT U9233 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .Y(
        io_fpu_fromint_data[32]) );
  NAND2X0_LVT U9234 ( .A1(n3787), .A2(n_T_427[545]), .Y(n7952) );
  NAND2X0_LVT U9235 ( .A1(n3665), .A2(n4408), .Y(n7951) );
  AO22X1_LVT U9236 ( .A1(n4021), .A2(n_T_427[673]), .A3(n3966), .A4(
        n_T_427[289]), .Y(n7948) );
  AO22X1_LVT U9237 ( .A1(n4036), .A2(n_T_427[353]), .A3(n4047), .A4(
        n_T_427[737]), .Y(n7947) );
  AO22X1_LVT U9238 ( .A1(n4024), .A2(n_T_427[928]), .A3(n4031), .A4(
        n_T_427[609]), .Y(n7945) );
  AO22X1_LVT U9239 ( .A1(n2858), .A2(n_T_427[161]), .A3(n4051), .A4(
        n_T_427[33]), .Y(n7944) );
  AO22X1_LVT U9240 ( .A1(n3963), .A2(n_T_427[481]), .A3(n2836), .A4(
        n_T_427[97]), .Y(n7943) );
  OR3X1_LVT U9241 ( .A1(n7945), .A2(n7944), .A3(n7943), .Y(n7946) );
  OR3X1_LVT U9242 ( .A1(n7948), .A2(n7947), .A3(n7946), .Y(n7949) );
  NAND2X0_LVT U9243 ( .A1(n4053), .A2(n7949), .Y(n7950) );
  AND2X1_LVT U9244 ( .A1(n3983), .A2(n8105), .Y(n9058) );
  NAND2X0_LVT U9245 ( .A1(n3624), .A2(n_T_427[225]), .Y(n7954) );
  NAND2X0_LVT U9246 ( .A1(n3661), .A2(n_T_427[864]), .Y(n7953) );
  NAND2X0_LVT U9247 ( .A1(n3635), .A2(n_T_427[1248]), .Y(n7956) );
  NAND2X0_LVT U9248 ( .A1(n3668), .A2(n_T_427[1120]), .Y(n7955) );
  NAND2X0_LVT U9249 ( .A1(n3760), .A2(n_T_427[992]), .Y(n7958) );
  NAND2X0_LVT U9250 ( .A1(n4014), .A2(n_T_427[1056]), .Y(n7957) );
  NAND2X0_LVT U9251 ( .A1(n3605), .A2(n_T_427[1376]), .Y(n7959) );
  NAND2X0_LVT U9252 ( .A1(n2966), .A2(n_T_427[1440]), .Y(n7961) );
  NAND2X0_LVT U9253 ( .A1(n3991), .A2(n_T_427[1913]), .Y(n7960) );
  AND3X1_LVT U9254 ( .A1(n7962), .A2(n7961), .A3(n7960), .Y(n7965) );
  NAND2X0_LVT U9255 ( .A1(n3600), .A2(n_T_427[800]), .Y(n7964) );
  OA21X1_LVT U9256 ( .A1(n3399), .A2(n3601), .A3(n7966), .Y(n7969) );
  NAND2X0_LVT U9257 ( .A1(n2093), .A2(n_T_427[1312]), .Y(n7968) );
  NAND2X0_LVT U9258 ( .A1(n2092), .A2(n_T_427[1760]), .Y(n7967) );
  NAND3X0_LVT U9259 ( .A1(n7969), .A2(n7968), .A3(n7967), .Y(n7974) );
  NAND2X0_LVT U9260 ( .A1(n3769), .A2(n_T_427[1504]), .Y(n7970) );
  NAND2X0_LVT U9261 ( .A1(n3621), .A2(n_T_427[1568]), .Y(n7972) );
  NAND2X0_LVT U9262 ( .A1(n3650), .A2(n_T_427[1632]), .Y(n7971) );
  NAND2X0_LVT U9263 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[33]), .Y(n7978) );
  NAND2X0_LVT U9264 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[33]), .Y(n7977)
         );
  NAND2X0_LVT U9265 ( .A1(n2493), .A2(n_T_628[33]), .Y(n7976) );
  NAND2X0_LVT U9266 ( .A1(n9066), .A2(n_T_918[33]), .Y(n7975) );
  NAND4X0_LVT U9267 ( .A1(n7978), .A2(n7977), .A3(n7976), .A4(n7975), .Y(
        io_fpu_fromint_data[33]) );
  AND2X1_LVT U9268 ( .A1(n4031), .A2(n2135), .Y(n8837) );
  NAND2X0_LVT U9269 ( .A1(n8837), .A2(n_T_427[610]), .Y(n7986) );
  NAND2X0_LVT U9270 ( .A1(n3665), .A2(n4411), .Y(n7985) );
  AO22X1_LVT U9271 ( .A1(n3970), .A2(n_T_427[418]), .A3(n4020), .A4(
        n_T_427[674]), .Y(n7982) );
  AO22X1_LVT U9272 ( .A1(n4024), .A2(n_T_427[929]), .A3(n3986), .A4(
        n_T_427[226]), .Y(n7981) );
  AO22X1_LVT U9273 ( .A1(n2837), .A2(n_T_427[98]), .A3(n4037), .A4(
        n_T_427[354]), .Y(n7980) );
  AO22X1_LVT U9274 ( .A1(n3982), .A2(n_T_427[801]), .A3(n4051), .A4(
        n_T_427[34]), .Y(n7979) );
  NOR4X1_LVT U9275 ( .A1(n7982), .A2(n7981), .A3(n7980), .A4(n7979), .Y(n7983)
         );
  OR2X1_LVT U9276 ( .A1(n7983), .A2(n2154), .Y(n7984) );
  AND3X1_LVT U9277 ( .A1(n7986), .A2(n7985), .A3(n7984), .Y(n7989) );
  NAND2X0_LVT U9278 ( .A1(n3788), .A2(n_T_427[546]), .Y(n7988) );
  NAND2X0_LVT U9279 ( .A1(n_T_427[482]), .A2(n3614), .Y(n7987) );
  NAND2X0_LVT U9280 ( .A1(n8991), .A2(n_T_427[865]), .Y(n7990) );
  OA21X1_LVT U9281 ( .A1(n3691), .A2(n3141), .A3(n7990), .Y(n7993) );
  NAND2X0_LVT U9282 ( .A1(n3790), .A2(n_T_427[290]), .Y(n7992) );
  NAND2X0_LVT U9283 ( .A1(n3713), .A2(n_T_427[162]), .Y(n7991) );
  NAND2X0_LVT U9284 ( .A1(n3605), .A2(n_T_427[1377]), .Y(n7994) );
  OA21X1_LVT U9285 ( .A1(n3452), .A2(n3767), .A3(n7994), .Y(n7997) );
  NAND2X0_LVT U9286 ( .A1(n3628), .A2(n_T_427[1441]), .Y(n7996) );
  NAND2X0_LVT U9287 ( .A1(n2998), .A2(n_T_427[1914]), .Y(n7995) );
  NAND2X0_LVT U9288 ( .A1(n2922), .A2(n_T_427[1697]), .Y(n7998) );
  OA21X1_LVT U9289 ( .A1(n3453), .A2(n3601), .A3(n7998), .Y(n8001) );
  NAND2X0_LVT U9290 ( .A1(n2094), .A2(n_T_427[1313]), .Y(n8000) );
  NAND2X0_LVT U9291 ( .A1(n4003), .A2(n_T_427[1761]), .Y(n7999) );
  NAND2X0_LVT U9292 ( .A1(n3769), .A2(n_T_427[1505]), .Y(n8002) );
  OA21X1_LVT U9293 ( .A1(n4010), .A2(n3335), .A3(n8002), .Y(n8005) );
  NAND2X0_LVT U9294 ( .A1(n3619), .A2(n_T_427[1569]), .Y(n8004) );
  NAND2X0_LVT U9295 ( .A1(n_T_427[1633]), .A2(n3643), .Y(n8003) );
  NAND2X0_LVT U9296 ( .A1(n_T_427[1249]), .A2(n3641), .Y(n8007) );
  NAND2X0_LVT U9297 ( .A1(n3674), .A2(n_T_427[1121]), .Y(n8006) );
  NAND2X0_LVT U9298 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[34]), .Y(n8012) );
  NAND2X0_LVT U9299 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[34]), .Y(n8011)
         );
  NAND2X0_LVT U9300 ( .A1(n2493), .A2(n_T_628[34]), .Y(n8010) );
  NAND2X0_LVT U9301 ( .A1(n9066), .A2(n_T_918[34]), .Y(n8009) );
  NAND4X0_LVT U9302 ( .A1(n8012), .A2(n8011), .A3(n8010), .A4(n8009), .Y(
        io_fpu_fromint_data[34]) );
  NAND2X0_LVT U9303 ( .A1(n3661), .A2(n_T_427[866]), .Y(n8013) );
  OA21X1_LVT U9304 ( .A1(n3400), .A2(n3691), .A3(n8013), .Y(n8022) );
  AO22X1_LVT U9305 ( .A1(n4024), .A2(n_T_427[930]), .A3(n3960), .A4(
        n_T_427[483]), .Y(n8017) );
  AO22X1_LVT U9306 ( .A1(n3967), .A2(n_T_427[291]), .A3(n4037), .A4(
        n_T_427[355]), .Y(n8016) );
  AO22X1_LVT U9307 ( .A1(n3975), .A2(n_T_427[163]), .A3(n4052), .A4(
        n_T_427[35]), .Y(n8015) );
  AO22X1_LVT U9308 ( .A1(n4034), .A2(n_T_427[611]), .A3(n3986), .A4(
        n_T_427[227]), .Y(n8014) );
  NOR4X1_LVT U9309 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .Y(n8019)
         );
  NAND2X0_LVT U9310 ( .A1(n2982), .A2(n4413), .Y(n8018) );
  OA21X1_LVT U9311 ( .A1(n8019), .A2(n3612), .A3(n8018), .Y(n8021) );
  NAND2X0_LVT U9312 ( .A1(n3788), .A2(n_T_427[547]), .Y(n8020) );
  NAND2X0_LVT U9313 ( .A1(n2135), .A2(n4022), .Y(n8996) );
  NAND2X0_LVT U9314 ( .A1(n_T_427[99]), .A2(n3707), .Y(n8023) );
  OA21X1_LVT U9315 ( .A1(n3369), .A2(n8996), .A3(n8023), .Y(n8026) );
  NAND2X0_LVT U9316 ( .A1(n3600), .A2(n_T_427[802]), .Y(n8024) );
  NAND2X0_LVT U9317 ( .A1(n3609), .A2(n_T_427[1378]), .Y(n8027) );
  NAND2X0_LVT U9318 ( .A1(n2966), .A2(n_T_427[1442]), .Y(n8029) );
  NAND2X0_LVT U9319 ( .A1(n2882), .A2(n_T_427[1915]), .Y(n8028) );
  NAND2X0_LVT U9320 ( .A1(n2922), .A2(n_T_427[1698]), .Y(n8031) );
  OA21X1_LVT U9321 ( .A1(n3401), .A2(n3601), .A3(n8031), .Y(n8034) );
  NAND2X0_LVT U9322 ( .A1(n2094), .A2(n_T_427[1314]), .Y(n8033) );
  NAND2X0_LVT U9323 ( .A1(n2092), .A2(n_T_427[1762]), .Y(n8032) );
  NAND2X0_LVT U9324 ( .A1(n3769), .A2(n_T_427[1506]), .Y(n8035) );
  OA21X1_LVT U9325 ( .A1(n2081), .A2(n3299), .A3(n8035), .Y(n8038) );
  NAND2X0_LVT U9326 ( .A1(n3618), .A2(n_T_427[1570]), .Y(n8037) );
  NAND2X0_LVT U9327 ( .A1(n3648), .A2(n_T_427[1634]), .Y(n8036) );
  NAND2X0_LVT U9328 ( .A1(n_T_427[1250]), .A2(n3635), .Y(n8040) );
  NAND2X0_LVT U9329 ( .A1(n3674), .A2(n_T_427[1122]), .Y(n8039) );
  NAND2X0_LVT U9330 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[35]), .Y(n8045) );
  NAND2X0_LVT U9331 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[35]), .Y(n8044)
         );
  NAND2X0_LVT U9332 ( .A1(n2493), .A2(n_T_628[35]), .Y(n8043) );
  NAND2X0_LVT U9333 ( .A1(n9066), .A2(n_T_918[35]), .Y(n8042) );
  NAND4X0_LVT U9334 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .Y(
        io_fpu_fromint_data[35]) );
  NAND2X0_LVT U9335 ( .A1(n2967), .A2(n_T_427[1443]), .Y(n8047) );
  AND3X1_LVT U9336 ( .A1(n8048), .A2(n8047), .A3(n8046), .Y(n8051) );
  NAND2X0_LVT U9337 ( .A1(n3789), .A2(n_T_427[292]), .Y(n8050) );
  NAND2X0_LVT U9338 ( .A1(n3771), .A2(n_T_427[739]), .Y(n8049) );
  NAND2X0_LVT U9339 ( .A1(n3998), .A2(n_T_427[1315]), .Y(n8053) );
  NAND2X0_LVT U9340 ( .A1(n4003), .A2(n_T_427[1763]), .Y(n8052) );
  NAND3X0_LVT U9341 ( .A1(n8053), .A2(n8052), .A3(n8054), .Y(n8060) );
  NAND2X0_LVT U9342 ( .A1(n2922), .A2(n_T_427[1699]), .Y(n8055) );
  OA21X1_LVT U9343 ( .A1(n3753), .A2(n3454), .A3(n8055), .Y(n8058) );
  NAND2X0_LVT U9344 ( .A1(n3620), .A2(n_T_427[1571]), .Y(n8057) );
  NAND2X0_LVT U9345 ( .A1(n_T_427[1635]), .A2(n3650), .Y(n8056) );
  NAND3X0_LVT U9346 ( .A1(n8058), .A2(n8057), .A3(n8056), .Y(n8059) );
  NAND2X0_LVT U9347 ( .A1(n3673), .A2(n_T_427[1123]), .Y(n8062) );
  NAND2X0_LVT U9348 ( .A1(n3759), .A2(n_T_427[995]), .Y(n8061) );
  NAND2X0_LVT U9349 ( .A1(n8062), .A2(n8061), .Y(n8079) );
  NAND2X0_LVT U9350 ( .A1(n3661), .A2(n_T_427[867]), .Y(n8073) );
  AO22X1_LVT U9351 ( .A1(n4039), .A2(n_T_427[356]), .A3(n4041), .A4(
        n_T_427[100]), .Y(n8069) );
  AO22X1_LVT U9352 ( .A1(n3973), .A2(n_T_427[164]), .A3(n3979), .A4(
        n_T_427[803]), .Y(n8068) );
  AOI22X1_LVT U9353 ( .A1(n4025), .A2(n_T_427[931]), .A3(n4031), .A4(
        n_T_427[612]), .Y(n8066) );
  AOI22X1_LVT U9354 ( .A1(n4022), .A2(n_T_427[676]), .A3(n3976), .A4(
        n_T_427[548]), .Y(n8065) );
  AOI22X1_LVT U9355 ( .A1(n3971), .A2(n_T_427[420]), .A3(n3960), .A4(
        n_T_427[484]), .Y(n8064) );
  NAND2X0_LVT U9356 ( .A1(n4052), .A2(n_T_427[36]), .Y(n8063) );
  NAND4X0_LVT U9357 ( .A1(n8066), .A2(n8065), .A3(n8064), .A4(n8063), .Y(n8067) );
  OR3X1_LVT U9358 ( .A1(n8069), .A2(n8068), .A3(n8067), .Y(n8070) );
  NAND2X0_LVT U9359 ( .A1(n4053), .A2(n8070), .Y(n8071) );
  NAND3X0_LVT U9360 ( .A1(n8073), .A2(n8072), .A3(n8071), .Y(n8078) );
  NAND2X0_LVT U9361 ( .A1(n3635), .A2(n_T_427[1251]), .Y(n8074) );
  NAND2X0_LVT U9362 ( .A1(n4014), .A2(n_T_427[1059]), .Y(n8075) );
  NAND2X0_LVT U9363 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[36]), .Y(n8084) );
  NAND2X0_LVT U9364 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[36]), .Y(n8083)
         );
  NAND2X0_LVT U9365 ( .A1(n2497), .A2(n_T_628[36]), .Y(n8082) );
  NAND2X0_LVT U9366 ( .A1(n9066), .A2(n_T_918[36]), .Y(n8081) );
  NAND4X0_LVT U9367 ( .A1(n8084), .A2(n8083), .A3(n8082), .A4(n8081), .Y(
        io_fpu_fromint_data[36]) );
  NAND2X0_LVT U9368 ( .A1(n3789), .A2(n_T_427[293]), .Y(n8094) );
  NAND2X0_LVT U9369 ( .A1(n3060), .A2(n4419), .Y(n8093) );
  AO22X1_LVT U9370 ( .A1(n8980), .A2(n_T_427[549]), .A3(n4043), .A4(
        n_T_427[101]), .Y(n8090) );
  AO22X1_LVT U9371 ( .A1(n4021), .A2(n_T_427[677]), .A3(n4037), .A4(
        n_T_427[357]), .Y(n8089) );
  AO22X1_LVT U9372 ( .A1(n4024), .A2(n_T_427[932]), .A3(n3960), .A4(
        n_T_427[485]), .Y(n8087) );
  AO22X1_LVT U9373 ( .A1(n3982), .A2(n_T_427[804]), .A3(n4047), .A4(
        n_T_427[740]), .Y(n8086) );
  AO22X1_LVT U9374 ( .A1(n4034), .A2(n_T_427[613]), .A3(n4028), .A4(
        n_T_427[868]), .Y(n8085) );
  OR3X1_LVT U9375 ( .A1(n8087), .A2(n8086), .A3(n8085), .Y(n8088) );
  OR3X1_LVT U9376 ( .A1(n8090), .A2(n8089), .A3(n8088), .Y(n8091) );
  NAND2X0_LVT U9377 ( .A1(n4053), .A2(n8091), .Y(n8092) );
  NAND2X0_LVT U9378 ( .A1(n3745), .A2(n_T_427[229]), .Y(n8096) );
  NAND2X0_LVT U9379 ( .A1(n3713), .A2(n_T_427[165]), .Y(n8095) );
  NAND2X0_LVT U9380 ( .A1(n3635), .A2(n_T_427[1252]), .Y(n8098) );
  NAND2X0_LVT U9381 ( .A1(n3670), .A2(n_T_427[1124]), .Y(n8097) );
  NAND2X0_LVT U9382 ( .A1(n3761), .A2(n_T_427[996]), .Y(n8100) );
  NAND2X0_LVT U9383 ( .A1(n3716), .A2(n_T_427[1060]), .Y(n8099) );
  NAND2X0_LVT U9384 ( .A1(n3607), .A2(n_T_427[1380]), .Y(n8101) );
  NAND2X0_LVT U9385 ( .A1(n3630), .A2(n_T_427[1444]), .Y(n8103) );
  NAND2X0_LVT U9386 ( .A1(n2985), .A2(n_T_427[1917]), .Y(n8102) );
  AND3X1_LVT U9387 ( .A1(n8104), .A2(n8103), .A3(n8102), .Y(n8108) );
  NAND2X0_LVT U9388 ( .A1(n3647), .A2(n_T_427[37]), .Y(n8107) );
  NAND2X0_LVT U9389 ( .A1(n3689), .A2(n_T_427[1700]), .Y(n8109) );
  OA21X1_LVT U9390 ( .A1(n3456), .A2(n3601), .A3(n8109), .Y(n8112) );
  NAND2X0_LVT U9391 ( .A1(n4000), .A2(n_T_427[1316]), .Y(n8111) );
  NAND2X0_LVT U9392 ( .A1(n4001), .A2(n_T_427[1764]), .Y(n8110) );
  NAND2X0_LVT U9393 ( .A1(n3769), .A2(n_T_427[1508]), .Y(n8113) );
  NAND2X0_LVT U9394 ( .A1(n3618), .A2(n_T_427[1572]), .Y(n8115) );
  NAND2X0_LVT U9395 ( .A1(n3642), .A2(n_T_427[1636]), .Y(n8114) );
  NAND2X0_LVT U9396 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[37]), .Y(n8120) );
  NAND2X0_LVT U9397 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[37]), .Y(n8119)
         );
  NAND2X0_LVT U9398 ( .A1(n2493), .A2(n_T_628[37]), .Y(n8118) );
  NAND2X0_LVT U9399 ( .A1(n9066), .A2(n_T_918[37]), .Y(n8117) );
  NAND4X0_LVT U9400 ( .A1(n8120), .A2(n8119), .A3(n8118), .A4(n8117), .Y(
        io_fpu_fromint_data[37]) );
  NAND2X0_LVT U9401 ( .A1(n8994), .A2(n_T_427[102]), .Y(n8123) );
  NAND2X0_LVT U9402 ( .A1(n3630), .A2(n_T_427[1445]), .Y(n8122) );
  NAND2X0_LVT U9403 ( .A1(n2985), .A2(n_T_427[1918]), .Y(n8121) );
  AND3X1_LVT U9404 ( .A1(n8123), .A2(n8122), .A3(n8121), .Y(n8126) );
  NAND2X0_LVT U9405 ( .A1(n3771), .A2(n_T_427[741]), .Y(n8124) );
  NAND2X0_LVT U9406 ( .A1(n3606), .A2(n_T_427[1381]), .Y(n8127) );
  OA21X1_LVT U9407 ( .A1(n3481), .A2(n9006), .A3(n8127), .Y(n8130) );
  NAND2X0_LVT U9408 ( .A1(n3999), .A2(n_T_427[1317]), .Y(n8129) );
  NAND2X0_LVT U9409 ( .A1(n4001), .A2(n_T_427[1765]), .Y(n8128) );
  OA21X1_LVT U9410 ( .A1(n3402), .A2(n3753), .A3(n8131), .Y(n8134) );
  NAND2X0_LVT U9411 ( .A1(n3621), .A2(n_T_427[1573]), .Y(n8133) );
  NAND2X0_LVT U9412 ( .A1(n3642), .A2(n_T_427[1637]), .Y(n8132) );
  NAND2X0_LVT U9413 ( .A1(n3670), .A2(n_T_427[1125]), .Y(n8136) );
  NAND2X0_LVT U9414 ( .A1(n3756), .A2(n_T_427[997]), .Y(n8135) );
  NAND2X0_LVT U9415 ( .A1(n3714), .A2(n_T_427[166]), .Y(n8147) );
  NAND2X0_LVT U9416 ( .A1(n2982), .A2(n4421), .Y(n8146) );
  AO22X1_LVT U9417 ( .A1(n3970), .A2(n_T_427[422]), .A3(n4037), .A4(
        n_T_427[358]), .Y(n8143) );
  AO22X1_LVT U9418 ( .A1(n3967), .A2(n_T_427[294]), .A3(n3979), .A4(
        n_T_427[805]), .Y(n8142) );
  AOI22X1_LVT U9419 ( .A1(n4035), .A2(n_T_427[614]), .A3(n4027), .A4(
        n_T_427[869]), .Y(n8140) );
  AOI22X1_LVT U9420 ( .A1(n3978), .A2(n_T_427[550]), .A3(n3983), .A4(
        n_T_427[230]), .Y(n8139) );
  AOI22X1_LVT U9421 ( .A1(n4024), .A2(n_T_427[933]), .A3(n4018), .A4(
        n_T_427[678]), .Y(n8138) );
  NAND2X0_LVT U9422 ( .A1(n4052), .A2(n_T_427[38]), .Y(n8137) );
  NAND4X0_LVT U9423 ( .A1(n8140), .A2(n8139), .A3(n8138), .A4(n8137), .Y(n8141) );
  OR3X1_LVT U9424 ( .A1(n8143), .A2(n8142), .A3(n8141), .Y(n8144) );
  NAND2X0_LVT U9425 ( .A1(n4053), .A2(n8144), .Y(n8145) );
  NAND2X0_LVT U9426 ( .A1(n3635), .A2(n_T_427[1253]), .Y(n8148) );
  NAND2X0_LVT U9427 ( .A1(n2611), .A2(n_T_427[1189]), .Y(n8150) );
  NAND2X0_LVT U9428 ( .A1(n3716), .A2(n_T_427[1061]), .Y(n8149) );
  NAND2X0_LVT U9429 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[38]), .Y(n8154) );
  NAND2X0_LVT U9430 ( .A1(n9065), .A2(io_imem_sfence_bits_addr[38]), .Y(n8153)
         );
  NAND2X0_LVT U9431 ( .A1(n2497), .A2(n_T_628[38]), .Y(n8152) );
  NAND2X0_LVT U9432 ( .A1(n9066), .A2(n_T_918[38]), .Y(n8151) );
  NAND4X0_LVT U9433 ( .A1(n8154), .A2(n8153), .A3(n8152), .A4(n8151), .Y(
        io_fpu_fromint_data[38]) );
  NAND2X0_LVT U9434 ( .A1(n3626), .A2(n_T_427[1446]), .Y(n8156) );
  NAND2X0_LVT U9435 ( .A1(n2986), .A2(n_T_427[1919]), .Y(n8155) );
  AND3X1_LVT U9436 ( .A1(n8157), .A2(n8156), .A3(n8155), .Y(n8160) );
  NAND2X0_LVT U9437 ( .A1(n3789), .A2(n_T_427[295]), .Y(n8159) );
  NAND2X0_LVT U9438 ( .A1(n3647), .A2(n_T_427[39]), .Y(n8158) );
  NAND2X0_LVT U9439 ( .A1(n3606), .A2(n_T_427[1382]), .Y(n8161) );
  OA21X1_LVT U9440 ( .A1(n3457), .A2(n9006), .A3(n8161), .Y(n8164) );
  NAND2X0_LVT U9441 ( .A1(n4000), .A2(n_T_427[1318]), .Y(n8163) );
  NAND2X0_LVT U9442 ( .A1(n2091), .A2(n_T_427[1766]), .Y(n8162) );
  NAND2X0_LVT U9443 ( .A1(n3689), .A2(n_T_427[1702]), .Y(n8165) );
  OA21X1_LVT U9444 ( .A1(n3458), .A2(n3753), .A3(n8165), .Y(n8168) );
  NAND2X0_LVT U9445 ( .A1(n3615), .A2(n_T_427[1574]), .Y(n8167) );
  NAND2X0_LVT U9446 ( .A1(n3649), .A2(n_T_427[1638]), .Y(n8166) );
  NAND2X0_LVT U9447 ( .A1(n3672), .A2(n_T_427[1126]), .Y(n8170) );
  NAND2X0_LVT U9448 ( .A1(n3757), .A2(n_T_427[998]), .Y(n8169) );
  NAND2X0_LVT U9449 ( .A1(n_T_427[167]), .A2(n3713), .Y(n8181) );
  NAND2X0_LVT U9450 ( .A1(n4015), .A2(n4424), .Y(n8180) );
  AO22X1_LVT U9451 ( .A1(n4021), .A2(n_T_427[679]), .A3(n4042), .A4(
        n_T_427[103]), .Y(n8177) );
  AO22X1_LVT U9452 ( .A1(n3982), .A2(n_T_427[806]), .A3(n4037), .A4(
        n_T_427[359]), .Y(n8176) );
  AOI22X1_LVT U9453 ( .A1(n4035), .A2(n_T_427[615]), .A3(n4027), .A4(
        n_T_427[870]), .Y(n8174) );
  AOI22X1_LVT U9454 ( .A1(n3978), .A2(n_T_427[551]), .A3(n3983), .A4(
        n_T_427[231]), .Y(n8173) );
  AOI22X1_LVT U9455 ( .A1(n4026), .A2(n_T_427[934]), .A3(n3960), .A4(
        n_T_427[487]), .Y(n8172) );
  NAND2X0_LVT U9456 ( .A1(n4048), .A2(n_T_427[742]), .Y(n8171) );
  NAND4X0_LVT U9457 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .Y(n8175) );
  OR3X1_LVT U9458 ( .A1(n8177), .A2(n8176), .A3(n8175), .Y(n8178) );
  NAND2X0_LVT U9459 ( .A1(n4053), .A2(n8178), .Y(n8179) );
  NAND2X0_LVT U9460 ( .A1(n3640), .A2(n_T_427[1254]), .Y(n8182) );
  NAND2X0_LVT U9461 ( .A1(n2611), .A2(n_T_427[1190]), .Y(n8184) );
  NAND2X0_LVT U9462 ( .A1(n3717), .A2(n_T_427[1062]), .Y(n8183) );
  NAND2X0_LVT U9463 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[39]), .Y(n8188) );
  NAND2X0_LVT U9464 ( .A1(n9065), .A2(n_T_1165[39]), .Y(n8187) );
  NAND2X0_LVT U9465 ( .A1(n2493), .A2(n_T_628[39]), .Y(n8186) );
  NAND2X0_LVT U9466 ( .A1(n9066), .A2(n_T_918[39]), .Y(n8185) );
  NAND4X0_LVT U9467 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .Y(
        io_fpu_fromint_data[39]) );
  NAND2X0_LVT U9468 ( .A1(n_T_427[1383]), .A2(n3611), .Y(n8189) );
  OA21X1_LVT U9469 ( .A1(n3147), .A2(n3988), .A3(n8189), .Y(n8192) );
  NAND2X0_LVT U9470 ( .A1(n2967), .A2(n_T_427[1447]), .Y(n8191) );
  NAND2X0_LVT U9471 ( .A1(n3992), .A2(n_T_427[1920]), .Y(n8190) );
  NAND3X0_LVT U9472 ( .A1(n8192), .A2(n8191), .A3(n8190), .Y(n8197) );
  NAND2X0_LVT U9473 ( .A1(n3657), .A2(n_T_427[1703]), .Y(n8193) );
  NAND2X0_LVT U9474 ( .A1(n3998), .A2(n_T_427[1319]), .Y(n8195) );
  NAND2X0_LVT U9475 ( .A1(n4003), .A2(n_T_427[1767]), .Y(n8194) );
  NAND2X0_LVT U9476 ( .A1(n3769), .A2(n_T_427[1511]), .Y(n8198) );
  OA21X1_LVT U9477 ( .A1(n4008), .A2(n3337), .A3(n8198), .Y(n8201) );
  NAND2X0_LVT U9478 ( .A1(n3621), .A2(n_T_427[1575]), .Y(n8200) );
  NAND2X0_LVT U9479 ( .A1(n3642), .A2(n_T_427[1639]), .Y(n8199) );
  NAND3X0_LVT U9480 ( .A1(n8201), .A2(n8200), .A3(n8199), .Y(n8206) );
  NAND2X0_LVT U9481 ( .A1(n3760), .A2(n_T_427[999]), .Y(n8202) );
  NAND2X0_LVT U9482 ( .A1(n_T_427[1255]), .A2(n3638), .Y(n8204) );
  NAND2X0_LVT U9483 ( .A1(n3668), .A2(n_T_427[1127]), .Y(n8203) );
  NAND2X0_LVT U9484 ( .A1(n3786), .A2(n_T_427[552]), .Y(n8214) );
  NAND2X0_LVT U9485 ( .A1(n3060), .A2(n4427), .Y(n8213) );
  AO22X1_LVT U9486 ( .A1(n4024), .A2(n_T_427[935]), .A3(n3960), .A4(
        n_T_427[488]), .Y(n8210) );
  AO22X1_LVT U9487 ( .A1(n4021), .A2(n_T_427[680]), .A3(n2836), .A4(
        n_T_427[104]), .Y(n8209) );
  AO22X1_LVT U9488 ( .A1(n3982), .A2(n_T_427[807]), .A3(n4037), .A4(
        n_T_427[360]), .Y(n8208) );
  AO22X1_LVT U9489 ( .A1(n4034), .A2(n_T_427[616]), .A3(n3986), .A4(
        n_T_427[232]), .Y(n8207) );
  NOR4X1_LVT U9490 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .Y(n8211)
         );
  OR2X1_LVT U9491 ( .A1(n8211), .A2(n3656), .Y(n8212) );
  NAND3X0_LVT U9492 ( .A1(n8214), .A2(n8213), .A3(n8212), .Y(n8222) );
  NAND2X0_LVT U9493 ( .A1(n3661), .A2(n_T_427[871]), .Y(n8216) );
  NAND2X0_LVT U9494 ( .A1(n3790), .A2(n_T_427[296]), .Y(n8215) );
  NAND2X0_LVT U9495 ( .A1(n8216), .A2(n8215), .Y(n8221) );
  NAND2X0_LVT U9496 ( .A1(n_T_427[168]), .A2(n3791), .Y(n8217) );
  OA21X1_LVT U9497 ( .A1(n3461), .A2(n3708), .A3(n8217), .Y(n8220) );
  NAND2X0_LVT U9498 ( .A1(n8944), .A2(n_T_427[40]), .Y(n8218) );
  NAND2X0_LVT U9499 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[40]), .Y(n8226) );
  NAND2X0_LVT U9500 ( .A1(n9065), .A2(n_T_1165[40]), .Y(n8225) );
  NAND2X0_LVT U9501 ( .A1(n2493), .A2(n_T_628[40]), .Y(n8224) );
  NAND2X0_LVT U9502 ( .A1(n9066), .A2(n_T_918[40]), .Y(n8223) );
  NAND4X0_LVT U9503 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8223), .Y(
        io_fpu_fromint_data[40]) );
  NAND2X0_LVT U9504 ( .A1(n_T_427[489]), .A2(n9052), .Y(n8228) );
  NAND2X0_LVT U9505 ( .A1(n3790), .A2(n_T_427[297]), .Y(n8227) );
  AND2X1_LVT U9506 ( .A1(n8228), .A2(n8227), .Y(n8237) );
  AO22X1_LVT U9507 ( .A1(n3970), .A2(n_T_427[425]), .A3(n4023), .A4(
        n_T_427[936]), .Y(n8232) );
  AO22X1_LVT U9508 ( .A1(n3982), .A2(n_T_427[808]), .A3(n4048), .A4(
        n_T_427[744]), .Y(n8231) );
  AO22X1_LVT U9509 ( .A1(n4034), .A2(n_T_427[617]), .A3(n3986), .A4(
        n_T_427[233]), .Y(n8230) );
  AO22X1_LVT U9510 ( .A1(n2836), .A2(n_T_427[105]), .A3(n4037), .A4(
        n_T_427[361]), .Y(n8229) );
  NOR4X1_LVT U9511 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8229), .Y(n8234)
         );
  NAND2X0_LVT U9512 ( .A1(n3060), .A2(n4430), .Y(n8233) );
  OA21X1_LVT U9513 ( .A1(n8234), .A2(n3612), .A3(n8233), .Y(n8236) );
  NAND2X0_LVT U9514 ( .A1(n3786), .A2(n_T_427[553]), .Y(n8235) );
  NAND2X0_LVT U9515 ( .A1(n8944), .A2(n_T_427[41]), .Y(n8238) );
  OA21X1_LVT U9516 ( .A1(n3404), .A2(n8996), .A3(n8238), .Y(n8241) );
  NAND2X0_LVT U9517 ( .A1(n3714), .A2(n_T_427[169]), .Y(n8240) );
  NAND2X0_LVT U9518 ( .A1(n8991), .A2(n_T_427[872]), .Y(n8239) );
  NAND2X0_LVT U9519 ( .A1(n3605), .A2(n_T_427[1384]), .Y(n8242) );
  NAND2X0_LVT U9520 ( .A1(n3627), .A2(n_T_427[1448]), .Y(n8244) );
  NAND2X0_LVT U9521 ( .A1(n2986), .A2(n_T_427[1921]), .Y(n8243) );
  NAND2X0_LVT U9522 ( .A1(n2093), .A2(n_T_427[1320]), .Y(n8248) );
  NAND2X0_LVT U9523 ( .A1(n4004), .A2(n_T_427[1768]), .Y(n8247) );
  NAND2X0_LVT U9524 ( .A1(n3770), .A2(n_T_427[1512]), .Y(n8250) );
  NAND2X0_LVT U9525 ( .A1(n_T_427[1576]), .A2(n3617), .Y(n8252) );
  NAND2X0_LVT U9526 ( .A1(n3650), .A2(n_T_427[1640]), .Y(n8251) );
  NAND2X0_LVT U9527 ( .A1(n_T_427[1256]), .A2(n3640), .Y(n8255) );
  NAND2X0_LVT U9528 ( .A1(n3668), .A2(n_T_427[1128]), .Y(n8254) );
  NAND2X0_LVT U9529 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[41]), .Y(n8260) );
  NAND2X0_LVT U9530 ( .A1(n9065), .A2(n_T_1165[41]), .Y(n8259) );
  NAND2X0_LVT U9531 ( .A1(n2497), .A2(n_T_628[41]), .Y(n8258) );
  NAND2X0_LVT U9532 ( .A1(n9066), .A2(n_T_918[41]), .Y(n8257) );
  NAND4X0_LVT U9533 ( .A1(n8260), .A2(n8259), .A3(n8258), .A4(n8257), .Y(
        io_fpu_fromint_data[41]) );
  NAND2X0_LVT U9534 ( .A1(n3771), .A2(n_T_427[745]), .Y(n8263) );
  NAND2X0_LVT U9535 ( .A1(n2966), .A2(n_T_427[1449]), .Y(n8262) );
  NAND2X0_LVT U9536 ( .A1(n2998), .A2(n_T_427[1922]), .Y(n8261) );
  AND3X1_LVT U9537 ( .A1(n8263), .A2(n8262), .A3(n8261), .Y(n8266) );
  NAND2X0_LVT U9538 ( .A1(n3787), .A2(n_T_427[554]), .Y(n8265) );
  NAND2X0_LVT U9539 ( .A1(n_T_427[1385]), .A2(n3611), .Y(n8267) );
  OA21X1_LVT U9540 ( .A1(n3149), .A2(n3989), .A3(n8267), .Y(n8270) );
  NAND2X0_LVT U9541 ( .A1(n3998), .A2(n_T_427[1321]), .Y(n8269) );
  NAND2X0_LVT U9542 ( .A1(n4003), .A2(n_T_427[1769]), .Y(n8268) );
  NAND3X0_LVT U9543 ( .A1(n8268), .A2(n8269), .A3(n8270), .Y(n8276) );
  NAND2X0_LVT U9544 ( .A1(n_T_427[1705]), .A2(n3689), .Y(n8271) );
  OA21X1_LVT U9545 ( .A1(n3462), .A2(n3753), .A3(n8271), .Y(n8274) );
  NAND2X0_LVT U9546 ( .A1(n3621), .A2(n_T_427[1577]), .Y(n8273) );
  NAND3X0_LVT U9547 ( .A1(n8274), .A2(n8273), .A3(n8272), .Y(n8275) );
  NAND2X0_LVT U9548 ( .A1(n3671), .A2(n_T_427[1129]), .Y(n8278) );
  NAND2X0_LVT U9549 ( .A1(n3712), .A2(n_T_427[1001]), .Y(n8277) );
  NAND2X0_LVT U9550 ( .A1(n4015), .A2(n4433), .Y(n8288) );
  AO22X1_LVT U9551 ( .A1(n4039), .A2(n_T_427[362]), .A3(n4044), .A4(
        n_T_427[106]), .Y(n8285) );
  AO22X1_LVT U9552 ( .A1(n2859), .A2(n_T_427[170]), .A3(n3979), .A4(
        n_T_427[809]), .Y(n8284) );
  AOI22X1_LVT U9553 ( .A1(n4035), .A2(n_T_427[618]), .A3(n4027), .A4(
        n_T_427[873]), .Y(n8282) );
  AOI22X1_LVT U9554 ( .A1(n4022), .A2(n_T_427[682]), .A3(n3983), .A4(
        n_T_427[234]), .Y(n8281) );
  AOI22X1_LVT U9555 ( .A1(n3971), .A2(n_T_427[426]), .A3(n4023), .A4(
        n_T_427[937]), .Y(n8280) );
  NAND2X0_LVT U9556 ( .A1(n4052), .A2(n_T_427[42]), .Y(n8279) );
  NAND4X0_LVT U9557 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8279), .Y(n8283) );
  OR3X1_LVT U9558 ( .A1(n8285), .A2(n8284), .A3(n8283), .Y(n8286) );
  NAND2X0_LVT U9559 ( .A1(n4053), .A2(n8286), .Y(n8287) );
  NAND2X0_LVT U9560 ( .A1(n_T_427[1257]), .A2(n3640), .Y(n8290) );
  OA21X1_LVT U9561 ( .A1(n3463), .A2(n2897), .A3(n8290), .Y(n8293) );
  NAND2X0_LVT U9562 ( .A1(n2611), .A2(n_T_427[1193]), .Y(n8292) );
  NAND2X0_LVT U9563 ( .A1(n4014), .A2(n_T_427[1065]), .Y(n8291) );
  NAND2X0_LVT U9564 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[42]), .Y(n8297) );
  NAND2X0_LVT U9565 ( .A1(n9065), .A2(n_T_1165[42]), .Y(n8296) );
  NAND2X0_LVT U9566 ( .A1(n2497), .A2(n_T_628[42]), .Y(n8295) );
  NAND2X0_LVT U9567 ( .A1(n9066), .A2(n_T_918[42]), .Y(n8294) );
  NAND4X0_LVT U9568 ( .A1(n8297), .A2(n8296), .A3(n8295), .A4(n8294), .Y(
        io_fpu_fromint_data[42]) );
  NAND2X0_LVT U9569 ( .A1(n3609), .A2(n_T_427[1386]), .Y(n8298) );
  OA21X1_LVT U9570 ( .A1(n3150), .A2(n3989), .A3(n8298), .Y(n8301) );
  NAND2X0_LVT U9571 ( .A1(n2967), .A2(n_T_427[1450]), .Y(n8300) );
  NAND2X0_LVT U9572 ( .A1(n3991), .A2(n_T_427[1923]), .Y(n8299) );
  NAND2X0_LVT U9573 ( .A1(n3689), .A2(n_T_427[1706]), .Y(n8302) );
  OA21X1_LVT U9574 ( .A1(n3464), .A2(n3994), .A3(n8302), .Y(n8305) );
  NAND2X0_LVT U9575 ( .A1(n3998), .A2(n_T_427[1322]), .Y(n8304) );
  NAND2X0_LVT U9576 ( .A1(n2091), .A2(n_T_427[1770]), .Y(n8303) );
  NAND2X0_LVT U9577 ( .A1(n3769), .A2(n_T_427[1514]), .Y(n8306) );
  OA21X1_LVT U9578 ( .A1(n4008), .A2(n3340), .A3(n8306), .Y(n8309) );
  NAND2X0_LVT U9579 ( .A1(n3616), .A2(n_T_427[1578]), .Y(n8308) );
  NAND2X0_LVT U9580 ( .A1(n_T_427[1642]), .A2(n3648), .Y(n8307) );
  NAND3X0_LVT U9581 ( .A1(n8307), .A2(n8308), .A3(n8309), .Y(n8314) );
  NAND2X0_LVT U9582 ( .A1(n3757), .A2(n_T_427[1002]), .Y(n8310) );
  NAND2X0_LVT U9583 ( .A1(n3637), .A2(n_T_427[1258]), .Y(n8312) );
  NAND2X0_LVT U9584 ( .A1(n3670), .A2(n_T_427[1130]), .Y(n8311) );
  NAND2X0_LVT U9585 ( .A1(n_T_427[938]), .A2(n8873), .Y(n8322) );
  AO22X1_LVT U9586 ( .A1(n3970), .A2(n_T_427[427]), .A3(n4021), .A4(
        n_T_427[683]), .Y(n8318) );
  AO22X1_LVT U9587 ( .A1(n3967), .A2(n_T_427[299]), .A3(n4052), .A4(
        n_T_427[43]), .Y(n8317) );
  AO22X1_LVT U9588 ( .A1(n4034), .A2(n_T_427[619]), .A3(n4027), .A4(
        n_T_427[874]), .Y(n8316) );
  AO22X1_LVT U9589 ( .A1(n2837), .A2(n_T_427[107]), .A3(n4037), .A4(
        n_T_427[363]), .Y(n8315) );
  NOR4X1_LVT U9590 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .Y(n8319)
         );
  NAND3X0_LVT U9591 ( .A1(n8321), .A2(n8322), .A3(n8320), .Y(n8329) );
  NAND2X0_LVT U9592 ( .A1(n_T_427[491]), .A2(n9052), .Y(n8325) );
  NAND2X0_LVT U9593 ( .A1(n_T_427[235]), .A2(n3624), .Y(n8324) );
  NAND3X0_LVT U9594 ( .A1(n8326), .A2(n8325), .A3(n8324), .Y(n8327) );
  NAND2X0_LVT U9595 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[43]), .Y(n8333) );
  NAND2X0_LVT U9596 ( .A1(n9065), .A2(n_T_1165[43]), .Y(n8332) );
  NAND2X0_LVT U9597 ( .A1(n2497), .A2(n_T_628[43]), .Y(n8331) );
  NAND2X0_LVT U9598 ( .A1(n9066), .A2(n_T_918[43]), .Y(n8330) );
  NAND4X0_LVT U9599 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .Y(
        io_fpu_fromint_data[43]) );
  NAND2X0_LVT U9600 ( .A1(n3787), .A2(n_T_427[556]), .Y(n8343) );
  NAND2X0_LVT U9601 ( .A1(n2982), .A2(n4439), .Y(n8342) );
  AO22X1_LVT U9602 ( .A1(n3963), .A2(n_T_427[492]), .A3(n4037), .A4(
        n_T_427[364]), .Y(n8339) );
  AO22X1_LVT U9603 ( .A1(n3970), .A2(n_T_427[428]), .A3(n3966), .A4(
        n_T_427[300]), .Y(n8338) );
  AO22X1_LVT U9604 ( .A1(n4024), .A2(n_T_427[939]), .A3(n4020), .A4(
        n_T_427[684]), .Y(n8336) );
  AO22X1_LVT U9605 ( .A1(n3974), .A2(n_T_427[172]), .A3(n4048), .A4(
        n_T_427[747]), .Y(n8335) );
  AO22X1_LVT U9606 ( .A1(n4034), .A2(n_T_427[620]), .A3(n4027), .A4(
        n_T_427[875]), .Y(n8334) );
  OR3X1_LVT U9607 ( .A1(n8336), .A2(n8335), .A3(n8334), .Y(n8337) );
  OR3X1_LVT U9608 ( .A1(n8339), .A2(n8338), .A3(n8337), .Y(n8340) );
  NAND2X0_LVT U9609 ( .A1(n4053), .A2(n8340), .Y(n8341) );
  NAND2X0_LVT U9610 ( .A1(n8944), .A2(n_T_427[44]), .Y(n8345) );
  NAND2X0_LVT U9611 ( .A1(n3745), .A2(n_T_427[236]), .Y(n8344) );
  NAND2X0_LVT U9612 ( .A1(n3635), .A2(n_T_427[1259]), .Y(n8347) );
  NAND2X0_LVT U9613 ( .A1(n3669), .A2(n_T_427[1131]), .Y(n8346) );
  AND2X1_LVT U9614 ( .A1(n8347), .A2(n8346), .Y(n8350) );
  NAND2X0_LVT U9615 ( .A1(n3761), .A2(n_T_427[1003]), .Y(n8349) );
  NAND2X0_LVT U9616 ( .A1(n3716), .A2(n_T_427[1067]), .Y(n8348) );
  NAND2X0_LVT U9617 ( .A1(n3602), .A2(n_T_427[1387]), .Y(n8351) );
  OA21X1_LVT U9618 ( .A1(n3465), .A2(n3988), .A3(n8351), .Y(n8354) );
  NAND2X0_LVT U9619 ( .A1(n3626), .A2(n_T_427[1451]), .Y(n8353) );
  AND3X1_LVT U9620 ( .A1(n8354), .A2(n8353), .A3(n8352), .Y(n8357) );
  NAND2X0_LVT U9621 ( .A1(n3600), .A2(n_T_427[811]), .Y(n8356) );
  NAND2X0_LVT U9622 ( .A1(n3707), .A2(n_T_427[108]), .Y(n8355) );
  NAND2X0_LVT U9623 ( .A1(n3657), .A2(n_T_427[1707]), .Y(n8358) );
  NAND2X0_LVT U9624 ( .A1(n2093), .A2(n_T_427[1323]), .Y(n8360) );
  NAND2X0_LVT U9625 ( .A1(n2092), .A2(n_T_427[1771]), .Y(n8359) );
  NAND2X0_LVT U9626 ( .A1(n3770), .A2(n_T_427[1515]), .Y(n8362) );
  NAND2X0_LVT U9627 ( .A1(n3619), .A2(n_T_427[1579]), .Y(n8364) );
  NAND2X0_LVT U9628 ( .A1(n3648), .A2(n_T_427[1643]), .Y(n8363) );
  NAND2X0_LVT U9629 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[44]), .Y(n8369) );
  NAND2X0_LVT U9630 ( .A1(n9065), .A2(n_T_1165[44]), .Y(n8368) );
  NAND2X0_LVT U9631 ( .A1(n2493), .A2(n_T_628[44]), .Y(n8367) );
  NAND2X0_LVT U9632 ( .A1(n9066), .A2(n_T_918[44]), .Y(n8366) );
  NAND4X0_LVT U9633 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), .Y(
        io_fpu_fromint_data[44]) );
  NAND2X0_LVT U9634 ( .A1(n_T_427[1388]), .A2(n3611), .Y(n8370) );
  OA21X1_LVT U9635 ( .A1(n3151), .A2(n3987), .A3(n8370), .Y(n8373) );
  NAND2X0_LVT U9636 ( .A1(n3628), .A2(n_T_427[1452]), .Y(n8372) );
  NAND2X0_LVT U9637 ( .A1(n2998), .A2(n_T_427[1925]), .Y(n8371) );
  NAND2X0_LVT U9638 ( .A1(n2922), .A2(n_T_427[1708]), .Y(n8374) );
  NAND2X0_LVT U9639 ( .A1(n3997), .A2(n_T_427[1324]), .Y(n8376) );
  NAND2X0_LVT U9640 ( .A1(n4004), .A2(n_T_427[1772]), .Y(n8375) );
  NAND2X0_LVT U9641 ( .A1(n3770), .A2(n_T_427[1516]), .Y(n8378) );
  OA21X1_LVT U9642 ( .A1(n3664), .A2(n3343), .A3(n8378), .Y(n8381) );
  NAND2X0_LVT U9643 ( .A1(n3615), .A2(n_T_427[1580]), .Y(n8380) );
  NAND2X0_LVT U9644 ( .A1(n3651), .A2(n_T_427[1644]), .Y(n8379) );
  NAND2X0_LVT U9645 ( .A1(n3761), .A2(n_T_427[1004]), .Y(n8382) );
  NAND2X0_LVT U9646 ( .A1(n3639), .A2(n_T_427[1260]), .Y(n8384) );
  NAND2X0_LVT U9647 ( .A1(n3671), .A2(n_T_427[1132]), .Y(n8383) );
  NAND2X0_LVT U9648 ( .A1(n8873), .A2(n_T_427[940]), .Y(n8390) );
  AO22X1_LVT U9649 ( .A1(n4021), .A2(n_T_427[685]), .A3(n3960), .A4(
        n_T_427[493]), .Y(n8387) );
  AO22X1_LVT U9650 ( .A1(n3978), .A2(n_T_427[557]), .A3(n4031), .A4(
        n_T_427[621]), .Y(n8386) );
  AO22X1_LVT U9651 ( .A1(n3967), .A2(n_T_427[301]), .A3(n4036), .A4(
        n_T_427[365]), .Y(n8385) );
  NAND3X0_LVT U9652 ( .A1(n8390), .A2(n8388), .A3(n8389), .Y(n8400) );
  NAND2X0_LVT U9653 ( .A1(n3661), .A2(n_T_427[876]), .Y(n8392) );
  NAND2X0_LVT U9654 ( .A1(n3624), .A2(n_T_427[237]), .Y(n8391) );
  NAND2X0_LVT U9655 ( .A1(n8392), .A2(n8391), .Y(n8399) );
  NAND2X0_LVT U9656 ( .A1(n8944), .A2(n_T_427[45]), .Y(n8394) );
  NAND2X0_LVT U9657 ( .A1(n8994), .A2(n_T_427[109]), .Y(n8393) );
  AND2X1_LVT U9658 ( .A1(n8394), .A2(n8393), .Y(n8397) );
  NAND2X0_LVT U9659 ( .A1(n3714), .A2(n_T_427[173]), .Y(n8396) );
  NAND3X0_LVT U9660 ( .A1(n8397), .A2(n8396), .A3(n8395), .Y(n8398) );
  NAND2X0_LVT U9661 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[45]), .Y(n8404) );
  NAND2X0_LVT U9662 ( .A1(n9065), .A2(n_T_1165[45]), .Y(n8403) );
  NAND2X0_LVT U9663 ( .A1(n2493), .A2(n_T_628[45]), .Y(n8402) );
  NAND2X0_LVT U9664 ( .A1(n9066), .A2(n_T_918[45]), .Y(n8401) );
  NAND4X0_LVT U9665 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .Y(
        io_fpu_fromint_data[45]) );
  NAND2X0_LVT U9666 ( .A1(n3610), .A2(n_T_427[1389]), .Y(n8405) );
  OA21X1_LVT U9667 ( .A1(n3466), .A2(n2969), .A3(n8405), .Y(n8408) );
  NAND2X0_LVT U9668 ( .A1(n2966), .A2(n_T_427[1453]), .Y(n8407) );
  NAND2X0_LVT U9669 ( .A1(n3991), .A2(n_T_427[1926]), .Y(n8406) );
  NAND2X0_LVT U9670 ( .A1(n3689), .A2(n_T_427[1709]), .Y(n8409) );
  OA21X1_LVT U9671 ( .A1(n3467), .A2(n3753), .A3(n8409), .Y(n8412) );
  NAND2X0_LVT U9672 ( .A1(n3996), .A2(n_T_427[1325]), .Y(n8411) );
  NAND2X0_LVT U9673 ( .A1(n4005), .A2(n_T_427[1773]), .Y(n8410) );
  NAND2X0_LVT U9674 ( .A1(n3770), .A2(n_T_427[1517]), .Y(n8413) );
  OA21X1_LVT U9675 ( .A1(n4008), .A2(n3345), .A3(n8413), .Y(n8416) );
  NAND2X0_LVT U9676 ( .A1(n3617), .A2(n_T_427[1581]), .Y(n8415) );
  NAND2X0_LVT U9677 ( .A1(n3650), .A2(n_T_427[1645]), .Y(n8414) );
  NAND2X0_LVT U9678 ( .A1(n3760), .A2(n_T_427[1005]), .Y(n8417) );
  NAND2X0_LVT U9679 ( .A1(n3640), .A2(n_T_427[1261]), .Y(n8419) );
  NAND2X0_LVT U9680 ( .A1(n3667), .A2(n_T_427[1133]), .Y(n8418) );
  NAND2X0_LVT U9681 ( .A1(n8939), .A2(n_T_427[366]), .Y(n8427) );
  AO22X1_LVT U9682 ( .A1(n4024), .A2(n_T_427[941]), .A3(n4021), .A4(
        n_T_427[686]), .Y(n8423) );
  AO22X1_LVT U9683 ( .A1(n3974), .A2(n_T_427[174]), .A3(n3966), .A4(
        n_T_427[302]), .Y(n8422) );
  AO22X1_LVT U9684 ( .A1(n3971), .A2(n_T_427[430]), .A3(n4041), .A4(
        n_T_427[110]), .Y(n8421) );
  AO22X1_LVT U9685 ( .A1(n4034), .A2(n_T_427[622]), .A3(n3986), .A4(
        n_T_427[238]), .Y(n8420) );
  NOR4X1_LVT U9686 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .Y(n8424)
         );
  NAND2X0_LVT U9687 ( .A1(n3786), .A2(n_T_427[558]), .Y(n8429) );
  NAND2X0_LVT U9688 ( .A1(n8991), .A2(n_T_427[877]), .Y(n8428) );
  NAND2X0_LVT U9689 ( .A1(n9056), .A2(n_T_427[813]), .Y(n8430) );
  OA21X1_LVT U9690 ( .A1(n3406), .A2(n3691), .A3(n8430), .Y(n8433) );
  NAND2X0_LVT U9691 ( .A1(n_T_427[494]), .A2(n9052), .Y(n8432) );
  NAND2X0_LVT U9692 ( .A1(n8944), .A2(n_T_427[46]), .Y(n8431) );
  NAND2X0_LVT U9693 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[46]), .Y(n8437) );
  NAND2X0_LVT U9694 ( .A1(n9065), .A2(n_T_1165[46]), .Y(n8436) );
  NAND2X0_LVT U9695 ( .A1(n2493), .A2(n_T_628[46]), .Y(n8435) );
  NAND2X0_LVT U9696 ( .A1(n9066), .A2(n_T_918[46]), .Y(n8434) );
  NAND4X0_LVT U9697 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .Y(
        io_fpu_fromint_data[46]) );
  NAND2X0_LVT U9698 ( .A1(n3610), .A2(n_T_427[1390]), .Y(n8438) );
  OA21X1_LVT U9699 ( .A1(n3152), .A2(n3989), .A3(n8438), .Y(n8441) );
  NAND2X0_LVT U9700 ( .A1(n3626), .A2(n_T_427[1454]), .Y(n8440) );
  NAND2X0_LVT U9701 ( .A1(n3992), .A2(n_T_427[1927]), .Y(n8439) );
  NAND2X0_LVT U9702 ( .A1(n3689), .A2(n_T_427[1710]), .Y(n8442) );
  NAND2X0_LVT U9703 ( .A1(n2094), .A2(n_T_427[1326]), .Y(n8444) );
  NAND2X0_LVT U9704 ( .A1(n2091), .A2(n_T_427[1774]), .Y(n8443) );
  NAND2X0_LVT U9705 ( .A1(n3770), .A2(n_T_427[1518]), .Y(n8446) );
  NAND2X0_LVT U9706 ( .A1(n3618), .A2(n_T_427[1582]), .Y(n8448) );
  NAND2X0_LVT U9707 ( .A1(n3642), .A2(n_T_427[1646]), .Y(n8447) );
  NAND2X0_LVT U9708 ( .A1(n3758), .A2(n_T_427[1006]), .Y(n8450) );
  NAND2X0_LVT U9709 ( .A1(n3639), .A2(n_T_427[1262]), .Y(n8452) );
  NAND2X0_LVT U9710 ( .A1(n3675), .A2(n_T_427[1134]), .Y(n8451) );
  NAND2X0_LVT U9711 ( .A1(n2982), .A2(n4448), .Y(n8459) );
  AO22X1_LVT U9712 ( .A1(n4024), .A2(n_T_427[942]), .A3(n4031), .A4(
        n_T_427[623]), .Y(n8456) );
  AO22X1_LVT U9713 ( .A1(n3978), .A2(n_T_427[559]), .A3(n3960), .A4(
        n_T_427[495]), .Y(n8455) );
  AO22X1_LVT U9714 ( .A1(n3971), .A2(n_T_427[431]), .A3(n4036), .A4(
        n_T_427[367]), .Y(n8454) );
  AO22X1_LVT U9715 ( .A1(n4052), .A2(n_T_427[47]), .A3(n4047), .A4(
        n_T_427[750]), .Y(n8453) );
  NOR4X1_LVT U9716 ( .A1(n8456), .A2(n8455), .A3(n8454), .A4(n8453), .Y(n8457)
         );
  NAND2X0_LVT U9717 ( .A1(n3714), .A2(n_T_427[175]), .Y(n8461) );
  NAND2X0_LVT U9718 ( .A1(n8991), .A2(n_T_427[878]), .Y(n8460) );
  NAND2X0_LVT U9719 ( .A1(n_T_427[111]), .A2(n8994), .Y(n8462) );
  OA21X1_LVT U9720 ( .A1(n3482), .A2(n8996), .A3(n8462), .Y(n8465) );
  NAND2X0_LVT U9721 ( .A1(n9056), .A2(n_T_427[814]), .Y(n8464) );
  NAND2X0_LVT U9722 ( .A1(n3624), .A2(n_T_427[239]), .Y(n8463) );
  NAND2X0_LVT U9723 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[47]), .Y(n8469) );
  NAND2X0_LVT U9724 ( .A1(n9065), .A2(n_T_1165[47]), .Y(n8468) );
  NAND2X0_LVT U9725 ( .A1(n2493), .A2(n_T_628[47]), .Y(n8467) );
  NAND2X0_LVT U9726 ( .A1(n9066), .A2(n_T_918[47]), .Y(n8466) );
  NAND4X0_LVT U9727 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), .Y(
        io_fpu_fromint_data[47]) );
  NAND2X0_LVT U9728 ( .A1(n3787), .A2(n_T_427[560]), .Y(n8476) );
  NAND2X0_LVT U9729 ( .A1(n3060), .A2(n4451), .Y(n8475) );
  AO22X1_LVT U9730 ( .A1(n4024), .A2(n_T_427[943]), .A3(n3966), .A4(
        n_T_427[304]), .Y(n8472) );
  AO22X1_LVT U9731 ( .A1(n4038), .A2(n_T_427[368]), .A3(n4048), .A4(
        n_T_427[751]), .Y(n8471) );
  OR3X1_LVT U9732 ( .A1(n8472), .A2(n8471), .A3(n8470), .Y(n8473) );
  NAND2X0_LVT U9733 ( .A1(n4053), .A2(n8473), .Y(n8474) );
  NAND2X0_LVT U9734 ( .A1(n_T_427[496]), .A2(n9052), .Y(n8478) );
  NAND2X0_LVT U9735 ( .A1(n9056), .A2(n_T_427[815]), .Y(n8477) );
  NAND2X0_LVT U9736 ( .A1(n3759), .A2(n_T_427[1007]), .Y(n8480) );
  NAND2X0_LVT U9737 ( .A1(n4014), .A2(n_T_427[1071]), .Y(n8479) );
  NAND2X0_LVT U9738 ( .A1(n3604), .A2(n_T_427[1391]), .Y(n8481) );
  OA21X1_LVT U9739 ( .A1(n3153), .A2(n3987), .A3(n8481), .Y(n8484) );
  NAND2X0_LVT U9740 ( .A1(n2966), .A2(n_T_427[1455]), .Y(n8483) );
  NAND2X0_LVT U9741 ( .A1(n3991), .A2(n_T_427[1928]), .Y(n8482) );
  AND3X1_LVT U9742 ( .A1(n8484), .A2(n8483), .A3(n8482), .Y(n8487) );
  NAND2X0_LVT U9743 ( .A1(n3707), .A2(n_T_427[112]), .Y(n8485) );
  NAND2X0_LVT U9744 ( .A1(n3689), .A2(n_T_427[1711]), .Y(n8488) );
  NAND2X0_LVT U9745 ( .A1(n3997), .A2(n_T_427[1327]), .Y(n8490) );
  NAND2X0_LVT U9746 ( .A1(n2091), .A2(n_T_427[1775]), .Y(n8489) );
  NAND3X0_LVT U9747 ( .A1(n8490), .A2(n8491), .A3(n8489), .Y(n8497) );
  OA21X1_LVT U9748 ( .A1(n4009), .A2(n3348), .A3(n8492), .Y(n8495) );
  NAND2X0_LVT U9749 ( .A1(n3620), .A2(n_T_427[1583]), .Y(n8494) );
  NAND3X0_LVT U9750 ( .A1(n8493), .A2(n8494), .A3(n8495), .Y(n8496) );
  NAND2X0_LVT U9751 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[48]), .Y(n8501) );
  NAND2X0_LVT U9752 ( .A1(n9065), .A2(n_T_1165[48]), .Y(n8500) );
  NAND2X0_LVT U9753 ( .A1(n2497), .A2(n_T_628[48]), .Y(n8499) );
  NAND2X0_LVT U9754 ( .A1(n9066), .A2(n_T_918[48]), .Y(n8498) );
  NAND4X0_LVT U9755 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .Y(
        io_fpu_fromint_data[48]) );
  NAND2X0_LVT U9756 ( .A1(n_T_427[1392]), .A2(n3611), .Y(n8502) );
  OA21X1_LVT U9757 ( .A1(n3154), .A2(n3988), .A3(n8502), .Y(n8505) );
  NAND2X0_LVT U9758 ( .A1(n3626), .A2(n_T_427[1456]), .Y(n8504) );
  NAND2X0_LVT U9759 ( .A1(n2986), .A2(n_T_427[1929]), .Y(n8503) );
  NAND2X0_LVT U9760 ( .A1(n3657), .A2(n_T_427[1712]), .Y(n8506) );
  OA21X1_LVT U9761 ( .A1(n3468), .A2(n3994), .A3(n8506), .Y(n8509) );
  NAND2X0_LVT U9762 ( .A1(n3997), .A2(n_T_427[1328]), .Y(n8508) );
  NAND2X0_LVT U9763 ( .A1(n4004), .A2(n_T_427[1776]), .Y(n8507) );
  NAND2X0_LVT U9764 ( .A1(n3769), .A2(n_T_427[1520]), .Y(n8510) );
  NAND2X0_LVT U9765 ( .A1(n3619), .A2(n_T_427[1584]), .Y(n8512) );
  NAND2X0_LVT U9766 ( .A1(n3648), .A2(n_T_427[1648]), .Y(n8511) );
  NAND2X0_LVT U9767 ( .A1(n3756), .A2(n_T_427[1008]), .Y(n8514) );
  NAND2X0_LVT U9768 ( .A1(n_T_427[1264]), .A2(n3636), .Y(n8516) );
  NAND2X0_LVT U9769 ( .A1(n3673), .A2(n_T_427[1136]), .Y(n8515) );
  NAND2X0_LVT U9770 ( .A1(n8837), .A2(n_T_427[625]), .Y(n8524) );
  NAND2X0_LVT U9771 ( .A1(n2982), .A2(n4454), .Y(n8523) );
  AO22X1_LVT U9772 ( .A1(n4021), .A2(n_T_427[689]), .A3(n3976), .A4(
        n_T_427[561]), .Y(n8520) );
  AO22X1_LVT U9773 ( .A1(n3971), .A2(n_T_427[433]), .A3(n4036), .A4(
        n_T_427[369]), .Y(n8519) );
  AO22X1_LVT U9774 ( .A1(n4023), .A2(n_T_427[944]), .A3(n3986), .A4(
        n_T_427[241]), .Y(n8518) );
  AO22X1_LVT U9775 ( .A1(n3967), .A2(n_T_427[305]), .A3(n4048), .A4(
        n_T_427[752]), .Y(n8517) );
  NOR4X1_LVT U9776 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .Y(n8521)
         );
  NAND2X0_LVT U9777 ( .A1(n_T_427[497]), .A2(n9052), .Y(n8526) );
  NAND2X0_LVT U9778 ( .A1(n_T_427[177]), .A2(n3713), .Y(n8525) );
  NAND2X0_LVT U9779 ( .A1(n8991), .A2(n_T_427[880]), .Y(n8528) );
  NAND2X0_LVT U9780 ( .A1(n9056), .A2(n_T_427[816]), .Y(n8527) );
  AND2X1_LVT U9781 ( .A1(n8528), .A2(n8527), .Y(n8531) );
  NAND2X0_LVT U9782 ( .A1(n8944), .A2(n_T_427[49]), .Y(n8530) );
  NAND2X0_LVT U9783 ( .A1(n8994), .A2(n_T_427[113]), .Y(n8529) );
  NAND2X0_LVT U9784 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[49]), .Y(n8535) );
  NAND2X0_LVT U9785 ( .A1(n9065), .A2(n_T_1165[49]), .Y(n8534) );
  NAND2X0_LVT U9786 ( .A1(n2493), .A2(n_T_628[49]), .Y(n8533) );
  NAND2X0_LVT U9787 ( .A1(n9066), .A2(n_T_918[49]), .Y(n8532) );
  NAND4X0_LVT U9788 ( .A1(n8535), .A2(n8534), .A3(n8533), .A4(n8532), .Y(
        io_fpu_fromint_data[49]) );
  NAND2X0_LVT U9789 ( .A1(n3759), .A2(n_T_427[1009]), .Y(n8536) );
  OA21X1_LVT U9790 ( .A1(n4012), .A2(n3351), .A3(n8536), .Y(n8539) );
  NAND2X0_LVT U9791 ( .A1(n3637), .A2(n_T_427[1265]), .Y(n8538) );
  NAND2X0_LVT U9792 ( .A1(n3670), .A2(n_T_427[1137]), .Y(n8537) );
  NAND2X0_LVT U9793 ( .A1(n3788), .A2(n_T_427[562]), .Y(n8549) );
  NAND2X0_LVT U9794 ( .A1(n2982), .A2(n4457), .Y(n8548) );
  AO22X1_LVT U9795 ( .A1(n3971), .A2(n_T_427[434]), .A3(n3966), .A4(
        n_T_427[306]), .Y(n8545) );
  AO22X1_LVT U9796 ( .A1(n3975), .A2(n_T_427[178]), .A3(n4036), .A4(
        n_T_427[370]), .Y(n8544) );
  AO22X1_LVT U9797 ( .A1(n4023), .A2(n_T_427[945]), .A3(n4031), .A4(
        n_T_427[626]), .Y(n8542) );
  AO22X1_LVT U9798 ( .A1(n4021), .A2(n_T_427[690]), .A3(n4043), .A4(
        n_T_427[114]), .Y(n8541) );
  AO22X1_LVT U9799 ( .A1(n3982), .A2(n_T_427[817]), .A3(n4052), .A4(
        n_T_427[50]), .Y(n8540) );
  OR3X1_LVT U9800 ( .A1(n8542), .A2(n8541), .A3(n8540), .Y(n8543) );
  OR3X1_LVT U9801 ( .A1(n8545), .A2(n8544), .A3(n8543), .Y(n8546) );
  NAND2X0_LVT U9802 ( .A1(n4053), .A2(n8546), .Y(n8547) );
  AND3X1_LVT U9803 ( .A1(n8549), .A2(n8548), .A3(n8547), .Y(n8552) );
  NAND2X0_LVT U9804 ( .A1(n8991), .A2(n_T_427[881]), .Y(n8551) );
  NAND2X0_LVT U9805 ( .A1(n2922), .A2(n_T_427[1713]), .Y(n8553) );
  NAND2X0_LVT U9806 ( .A1(n3996), .A2(n_T_427[1329]), .Y(n8555) );
  NAND2X0_LVT U9807 ( .A1(n4002), .A2(n_T_427[1777]), .Y(n8554) );
  NAND2X0_LVT U9808 ( .A1(n3770), .A2(n_T_427[1521]), .Y(n8557) );
  OA21X1_LVT U9809 ( .A1(n2081), .A2(n3352), .A3(n8557), .Y(n8560) );
  NAND2X0_LVT U9810 ( .A1(n3615), .A2(n_T_427[1585]), .Y(n8559) );
  NAND2X0_LVT U9811 ( .A1(n3650), .A2(n_T_427[1649]), .Y(n8558) );
  NAND2X0_LVT U9812 ( .A1(n_T_427[242]), .A2(n9058), .Y(n8561) );
  NAND2X0_LVT U9813 ( .A1(n3606), .A2(n_T_427[1393]), .Y(n8563) );
  OA21X1_LVT U9814 ( .A1(n3155), .A2(n2969), .A3(n8563), .Y(n8564) );
  NAND2X0_LVT U9815 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[50]), .Y(n8568) );
  NAND2X0_LVT U9816 ( .A1(n9065), .A2(n_T_1165[50]), .Y(n8567) );
  NAND2X0_LVT U9817 ( .A1(n2493), .A2(n_T_628[50]), .Y(n8566) );
  NAND2X0_LVT U9818 ( .A1(n9066), .A2(n_T_918[50]), .Y(n8565) );
  NAND4X0_LVT U9819 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .Y(
        io_fpu_fromint_data[50]) );
  NAND2X0_LVT U9820 ( .A1(n3608), .A2(n_T_427[1394]), .Y(n8569) );
  OA21X1_LVT U9821 ( .A1(n3156), .A2(n3988), .A3(n8569), .Y(n8572) );
  NAND2X0_LVT U9822 ( .A1(n3627), .A2(n_T_427[1458]), .Y(n8571) );
  NAND2X0_LVT U9823 ( .A1(n2985), .A2(n_T_427[1930]), .Y(n8570) );
  AND3X1_LVT U9824 ( .A1(n8572), .A2(n8571), .A3(n8570), .Y(n8575) );
  NAND2X0_LVT U9825 ( .A1(n3661), .A2(n_T_427[882]), .Y(n8574) );
  NAND2X0_LVT U9826 ( .A1(n3647), .A2(n_T_427[51]), .Y(n8573) );
  NAND2X0_LVT U9827 ( .A1(n3788), .A2(n_T_427[563]), .Y(n8586) );
  NAND2X0_LVT U9828 ( .A1(n3060), .A2(n4460), .Y(n8585) );
  AO22X1_LVT U9829 ( .A1(n4022), .A2(n_T_427[691]), .A3(n4036), .A4(
        n_T_427[371]), .Y(n8582) );
  AO22X1_LVT U9830 ( .A1(n4043), .A2(n_T_427[115]), .A3(n4048), .A4(
        n_T_427[754]), .Y(n8581) );
  AOI22X1_LVT U9831 ( .A1(n2859), .A2(n_T_427[179]), .A3(n3979), .A4(
        n_T_427[818]), .Y(n8579) );
  AOI22X1_LVT U9832 ( .A1(n3971), .A2(n_T_427[435]), .A3(n4023), .A4(
        n_T_427[946]), .Y(n8578) );
  NAND2X0_LVT U9833 ( .A1(n4031), .A2(n_T_427[627]), .Y(n8577) );
  NAND2X0_LVT U9834 ( .A1(n3986), .A2(n_T_427[243]), .Y(n8576) );
  NAND4X0_LVT U9835 ( .A1(n8579), .A2(n8578), .A3(n8577), .A4(n8576), .Y(n8580) );
  OR3X1_LVT U9836 ( .A1(n8582), .A2(n8581), .A3(n8580), .Y(n8583) );
  NAND2X0_LVT U9837 ( .A1(n4053), .A2(n8583), .Y(n8584) );
  NAND2X0_LVT U9838 ( .A1(n_T_427[499]), .A2(n9052), .Y(n8588) );
  NAND2X0_LVT U9839 ( .A1(n3789), .A2(n_T_427[307]), .Y(n8587) );
  NAND2X0_LVT U9840 ( .A1(n3641), .A2(n_T_427[1266]), .Y(n8590) );
  NAND2X0_LVT U9841 ( .A1(n3668), .A2(n_T_427[1138]), .Y(n8589) );
  NAND2X0_LVT U9842 ( .A1(n3689), .A2(n_T_427[1714]), .Y(n8591) );
  NAND2X0_LVT U9843 ( .A1(n3996), .A2(n_T_427[1330]), .Y(n8593) );
  NAND2X0_LVT U9844 ( .A1(n4005), .A2(n_T_427[1778]), .Y(n8592) );
  NAND3X0_LVT U9845 ( .A1(n8593), .A2(n8594), .A3(n8592), .Y(n8600) );
  NAND2X0_LVT U9846 ( .A1(n3769), .A2(n_T_427[1522]), .Y(n8595) );
  NAND2X0_LVT U9847 ( .A1(n3620), .A2(n_T_427[1586]), .Y(n8597) );
  NAND3X0_LVT U9848 ( .A1(n8598), .A2(n8597), .A3(n8596), .Y(n8599) );
  NAND2X0_LVT U9849 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[51]), .Y(n8604) );
  NAND2X0_LVT U9850 ( .A1(n9065), .A2(n_T_1165[51]), .Y(n8603) );
  NAND2X0_LVT U9851 ( .A1(n_T_628[51]), .A2(n2497), .Y(n8602) );
  NAND2X0_LVT U9852 ( .A1(n9066), .A2(n_T_918[51]), .Y(n8601) );
  NAND4X0_LVT U9853 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .Y(
        io_fpu_fromint_data[51]) );
  NAND2X0_LVT U9854 ( .A1(n3603), .A2(n_T_427[1395]), .Y(n8605) );
  OA21X1_LVT U9855 ( .A1(n3157), .A2(n3987), .A3(n8605), .Y(n8608) );
  NAND2X0_LVT U9856 ( .A1(n3627), .A2(n_T_427[1459]), .Y(n8607) );
  NAND2X0_LVT U9857 ( .A1(n3991), .A2(n_T_427[1931]), .Y(n8606) );
  NAND2X0_LVT U9858 ( .A1(n2922), .A2(n_T_427[1715]), .Y(n8609) );
  OA21X1_LVT U9859 ( .A1(n3469), .A2(n3994), .A3(n8609), .Y(n8612) );
  NAND2X0_LVT U9860 ( .A1(n3996), .A2(n_T_427[1331]), .Y(n8611) );
  NAND2X0_LVT U9861 ( .A1(n4002), .A2(n_T_427[1779]), .Y(n8610) );
  NAND2X0_LVT U9862 ( .A1(n3770), .A2(n_T_427[1523]), .Y(n8613) );
  OA21X1_LVT U9863 ( .A1(n4010), .A2(n3355), .A3(n8613), .Y(n8616) );
  NAND2X0_LVT U9864 ( .A1(n3617), .A2(n_T_427[1587]), .Y(n8615) );
  NAND2X0_LVT U9865 ( .A1(n3652), .A2(n_T_427[1651]), .Y(n8614) );
  NAND2X0_LVT U9866 ( .A1(n3761), .A2(n_T_427[1011]), .Y(n8617) );
  NAND2X0_LVT U9867 ( .A1(n3641), .A2(n_T_427[1267]), .Y(n8619) );
  NAND2X0_LVT U9868 ( .A1(n3673), .A2(n_T_427[1139]), .Y(n8618) );
  NAND2X0_LVT U9869 ( .A1(n3786), .A2(n_T_427[564]), .Y(n8627) );
  NAND2X0_LVT U9870 ( .A1(n3060), .A2(n4463), .Y(n8626) );
  AO22X1_LVT U9871 ( .A1(n4022), .A2(n_T_427[692]), .A3(n4036), .A4(
        n_T_427[372]), .Y(n8623) );
  AO22X1_LVT U9872 ( .A1(n4023), .A2(n_T_427[947]), .A3(n3986), .A4(
        n_T_427[244]), .Y(n8622) );
  AO22X1_LVT U9873 ( .A1(n4034), .A2(n_T_427[628]), .A3(n4027), .A4(
        n_T_427[883]), .Y(n8621) );
  AO22X1_LVT U9874 ( .A1(n3982), .A2(n_T_427[819]), .A3(n4052), .A4(
        n_T_427[52]), .Y(n8620) );
  NOR4X1_LVT U9875 ( .A1(n8623), .A2(n8622), .A3(n8621), .A4(n8620), .Y(n8624)
         );
  NAND2X0_LVT U9876 ( .A1(n_T_427[500]), .A2(n9052), .Y(n8629) );
  NAND2X0_LVT U9877 ( .A1(n3789), .A2(n_T_427[308]), .Y(n8628) );
  NAND2X0_LVT U9878 ( .A1(n_T_427[180]), .A2(n3791), .Y(n8630) );
  OA21X1_LVT U9879 ( .A1(n3408), .A2(n3691), .A3(n8630), .Y(n8632) );
  NAND2X0_LVT U9880 ( .A1(n_T_427[116]), .A2(n8994), .Y(n8631) );
  NAND2X0_LVT U9881 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[52]), .Y(n8636) );
  NAND2X0_LVT U9882 ( .A1(n9065), .A2(n_T_1165[52]), .Y(n8635) );
  NAND2X0_LVT U9883 ( .A1(n2497), .A2(n_T_628[52]), .Y(n8634) );
  NAND2X0_LVT U9884 ( .A1(n9066), .A2(n_T_918[52]), .Y(n8633) );
  NAND4X0_LVT U9885 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .Y(
        io_fpu_fromint_data[52]) );
  NAND2X0_LVT U9886 ( .A1(n3607), .A2(n_T_427[1396]), .Y(n8637) );
  OA21X1_LVT U9887 ( .A1(n3158), .A2(n3989), .A3(n8637), .Y(n8640) );
  NAND2X0_LVT U9888 ( .A1(n3627), .A2(n_T_427[1460]), .Y(n8639) );
  NAND2X0_LVT U9889 ( .A1(n3991), .A2(n_T_427[1932]), .Y(n8638) );
  AND3X1_LVT U9890 ( .A1(n8638), .A2(n8639), .A3(n8640), .Y(n8643) );
  NAND2X0_LVT U9891 ( .A1(n3647), .A2(n_T_427[53]), .Y(n8642) );
  NAND2X0_LVT U9892 ( .A1(n3786), .A2(n_T_427[565]), .Y(n8654) );
  NAND2X0_LVT U9893 ( .A1(n3665), .A2(n4466), .Y(n8653) );
  AO22X1_LVT U9894 ( .A1(n3963), .A2(n_T_427[501]), .A3(n4036), .A4(
        n_T_427[373]), .Y(n8650) );
  AO22X1_LVT U9895 ( .A1(n4042), .A2(n_T_427[117]), .A3(n4048), .A4(
        n_T_427[756]), .Y(n8649) );
  AOI22X1_LVT U9896 ( .A1(n3974), .A2(n_T_427[181]), .A3(n3979), .A4(
        n_T_427[820]), .Y(n8647) );
  AOI22X1_LVT U9897 ( .A1(n4023), .A2(n_T_427[948]), .A3(n4018), .A4(
        n_T_427[693]), .Y(n8646) );
  NAND2X0_LVT U9898 ( .A1(n4031), .A2(n_T_427[629]), .Y(n8645) );
  NAND2X0_LVT U9899 ( .A1(n3986), .A2(n_T_427[245]), .Y(n8644) );
  NAND4X0_LVT U9900 ( .A1(n8647), .A2(n8646), .A3(n8645), .A4(n8644), .Y(n8648) );
  OR3X1_LVT U9901 ( .A1(n8650), .A2(n8649), .A3(n8648), .Y(n8651) );
  NAND2X0_LVT U9902 ( .A1(n4053), .A2(n8651), .Y(n8652) );
  NAND2X0_LVT U9903 ( .A1(n8991), .A2(n_T_427[884]), .Y(n8656) );
  NAND2X0_LVT U9904 ( .A1(n3789), .A2(n_T_427[309]), .Y(n8655) );
  NAND2X0_LVT U9905 ( .A1(n3755), .A2(n_T_427[1012]), .Y(n8657) );
  OA21X1_LVT U9906 ( .A1(n4013), .A2(n3357), .A3(n8657), .Y(n8660) );
  NAND2X0_LVT U9907 ( .A1(n3637), .A2(n_T_427[1268]), .Y(n8659) );
  NAND2X0_LVT U9908 ( .A1(n3667), .A2(n_T_427[1140]), .Y(n8658) );
  NAND2X0_LVT U9909 ( .A1(n3689), .A2(n_T_427[1716]), .Y(n8661) );
  OA21X1_LVT U9910 ( .A1(n3470), .A2(n3601), .A3(n8661), .Y(n8664) );
  NAND2X0_LVT U9911 ( .A1(n2094), .A2(n_T_427[1332]), .Y(n8663) );
  NAND2X0_LVT U9912 ( .A1(n4002), .A2(n_T_427[1780]), .Y(n8662) );
  NAND3X0_LVT U9913 ( .A1(n8663), .A2(n8664), .A3(n8662), .Y(n8670) );
  NAND2X0_LVT U9914 ( .A1(n3770), .A2(n_T_427[1524]), .Y(n8665) );
  OA21X1_LVT U9915 ( .A1(n3663), .A2(n3358), .A3(n8665), .Y(n8668) );
  NAND2X0_LVT U9916 ( .A1(n3615), .A2(n_T_427[1588]), .Y(n8667) );
  NAND2X0_LVT U9917 ( .A1(n3650), .A2(n_T_427[1652]), .Y(n8666) );
  NAND3X0_LVT U9918 ( .A1(n8668), .A2(n8667), .A3(n8666), .Y(n8669) );
  NAND2X0_LVT U9919 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[53]), .Y(n8674) );
  NAND2X0_LVT U9920 ( .A1(n9065), .A2(n_T_1165[53]), .Y(n8673) );
  NAND2X0_LVT U9921 ( .A1(n_T_628[53]), .A2(n2493), .Y(n8672) );
  NAND2X0_LVT U9922 ( .A1(n9066), .A2(n_T_918[53]), .Y(n8671) );
  NAND4X0_LVT U9923 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .Y(
        io_fpu_fromint_data[53]) );
  NAND2X0_LVT U9924 ( .A1(n3607), .A2(n_T_427[1397]), .Y(n8675) );
  NAND2X0_LVT U9925 ( .A1(n3627), .A2(n_T_427[1461]), .Y(n8677) );
  NAND2X0_LVT U9926 ( .A1(n2882), .A2(n_T_427[1933]), .Y(n8676) );
  AND3X1_LVT U9927 ( .A1(n8678), .A2(n8677), .A3(n8676), .Y(n8681) );
  NAND2X0_LVT U9928 ( .A1(n3647), .A2(n_T_427[54]), .Y(n8680) );
  NAND2X0_LVT U9929 ( .A1(n3789), .A2(n_T_427[310]), .Y(n8692) );
  NAND2X0_LVT U9930 ( .A1(n2982), .A2(n4469), .Y(n8691) );
  AO22X1_LVT U9931 ( .A1(n3976), .A2(n_T_427[566]), .A3(n4042), .A4(
        n_T_427[118]), .Y(n8688) );
  AO22X1_LVT U9932 ( .A1(n4022), .A2(n_T_427[694]), .A3(n4036), .A4(
        n_T_427[374]), .Y(n8687) );
  AOI22X1_LVT U9933 ( .A1(n4023), .A2(n_T_427[949]), .A3(n3960), .A4(
        n_T_427[502]), .Y(n8685) );
  AOI22X1_LVT U9934 ( .A1(n3975), .A2(n_T_427[182]), .A3(n3979), .A4(
        n_T_427[821]), .Y(n8684) );
  NAND2X0_LVT U9935 ( .A1(n4031), .A2(n_T_427[630]), .Y(n8683) );
  NAND2X0_LVT U9936 ( .A1(n4030), .A2(n_T_427[885]), .Y(n8682) );
  NAND4X0_LVT U9937 ( .A1(n8685), .A2(n8684), .A3(n8683), .A4(n8682), .Y(n8686) );
  OR3X1_LVT U9938 ( .A1(n8688), .A2(n8687), .A3(n8686), .Y(n8689) );
  NAND2X0_LVT U9939 ( .A1(n4053), .A2(n8689), .Y(n8690) );
  NAND2X0_LVT U9940 ( .A1(n3712), .A2(n_T_427[1013]), .Y(n8693) );
  OA21X1_LVT U9941 ( .A1(n4012), .A2(n3359), .A3(n8693), .Y(n8696) );
  NAND2X0_LVT U9942 ( .A1(n3636), .A2(n_T_427[1269]), .Y(n8695) );
  NAND2X0_LVT U9943 ( .A1(n3668), .A2(n_T_427[1141]), .Y(n8694) );
  OA21X1_LVT U9944 ( .A1(n3471), .A2(n3601), .A3(n8697), .Y(n8700) );
  NAND2X0_LVT U9945 ( .A1(n3999), .A2(n_T_427[1333]), .Y(n8699) );
  NAND2X0_LVT U9946 ( .A1(n4004), .A2(n_T_427[1781]), .Y(n8698) );
  NAND3X0_LVT U9947 ( .A1(n8700), .A2(n8699), .A3(n8698), .Y(n8706) );
  NAND2X0_LVT U9948 ( .A1(n3770), .A2(n_T_427[1525]), .Y(n8701) );
  OA21X1_LVT U9949 ( .A1(n4009), .A2(n3360), .A3(n8701), .Y(n8704) );
  NAND2X0_LVT U9950 ( .A1(n3616), .A2(n_T_427[1589]), .Y(n8703) );
  NAND2X0_LVT U9951 ( .A1(n_T_427[1653]), .A2(n3651), .Y(n8702) );
  NAND3X0_LVT U9952 ( .A1(n8704), .A2(n8703), .A3(n8702), .Y(n8705) );
  NAND2X0_LVT U9953 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[54]), .Y(n8710) );
  NAND2X0_LVT U9954 ( .A1(n9065), .A2(n_T_1165[54]), .Y(n8709) );
  NAND2X0_LVT U9955 ( .A1(n2493), .A2(n_T_628[54]), .Y(n8708) );
  NAND2X0_LVT U9956 ( .A1(n9066), .A2(n_T_918[54]), .Y(n8707) );
  NAND4X0_LVT U9957 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .Y(
        io_fpu_fromint_data[54]) );
  NAND2X0_LVT U9958 ( .A1(n_T_427[503]), .A2(n9052), .Y(n8711) );
  OA21X1_LVT U9959 ( .A1(n3691), .A2(n3301), .A3(n8711), .Y(n8720) );
  AO22X1_LVT U9960 ( .A1(n4024), .A2(n_T_427[950]), .A3(n3976), .A4(
        n_T_427[567]), .Y(n8715) );
  AO22X1_LVT U9961 ( .A1(n3971), .A2(n_T_427[439]), .A3(n4021), .A4(
        n_T_427[695]), .Y(n8714) );
  AO22X1_LVT U9962 ( .A1(n3967), .A2(n_T_427[311]), .A3(n3979), .A4(
        n_T_427[822]), .Y(n8713) );
  AO22X1_LVT U9963 ( .A1(n4034), .A2(n_T_427[631]), .A3(n4027), .A4(
        n_T_427[886]), .Y(n8712) );
  NOR4X1_LVT U9964 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .Y(n8717)
         );
  NAND2X0_LVT U9965 ( .A1(n2982), .A2(n4472), .Y(n8716) );
  OA21X1_LVT U9966 ( .A1(n8717), .A2(n3612), .A3(n8716), .Y(n8719) );
  NAND2X0_LVT U9967 ( .A1(n8939), .A2(n_T_427[375]), .Y(n8718) );
  NAND2X0_LVT U9968 ( .A1(n3624), .A2(n_T_427[247]), .Y(n8722) );
  NAND2X0_LVT U9969 ( .A1(n8994), .A2(n_T_427[119]), .Y(n8721) );
  AND2X1_LVT U9970 ( .A1(n8722), .A2(n8721), .Y(n8725) );
  NAND2X0_LVT U9971 ( .A1(n_T_427[183]), .A2(n3714), .Y(n8724) );
  NAND2X0_LVT U9972 ( .A1(n3647), .A2(n_T_427[55]), .Y(n8723) );
  NAND2X0_LVT U9973 ( .A1(n3608), .A2(n_T_427[1398]), .Y(n8726) );
  OA21X1_LVT U9974 ( .A1(n3160), .A2(n2969), .A3(n8726), .Y(n8729) );
  NAND2X0_LVT U9975 ( .A1(n2967), .A2(n_T_427[1462]), .Y(n8728) );
  NAND2X0_LVT U9976 ( .A1(n2986), .A2(n_T_427[1934]), .Y(n8727) );
  NAND2X0_LVT U9977 ( .A1(n3657), .A2(n_T_427[1718]), .Y(n8730) );
  OA21X1_LVT U9978 ( .A1(n3161), .A2(n3751), .A3(n8730), .Y(n8733) );
  NAND2X0_LVT U9979 ( .A1(n2094), .A2(n_T_427[1334]), .Y(n8732) );
  NAND2X0_LVT U9980 ( .A1(n4001), .A2(n_T_427[1782]), .Y(n8731) );
  NAND2X0_LVT U9981 ( .A1(n3769), .A2(n_T_427[1526]), .Y(n8734) );
  OA21X1_LVT U9982 ( .A1(n4009), .A2(n3361), .A3(n8734), .Y(n8737) );
  NAND2X0_LVT U9983 ( .A1(n3616), .A2(n_T_427[1590]), .Y(n8736) );
  NAND2X0_LVT U9984 ( .A1(n3643), .A2(n_T_427[1654]), .Y(n8735) );
  NAND2X0_LVT U9985 ( .A1(n_T_427[1270]), .A2(n3636), .Y(n8739) );
  NAND2X0_LVT U9986 ( .A1(n3669), .A2(n_T_427[1142]), .Y(n8738) );
  NAND2X0_LVT U9987 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[55]), .Y(n8744) );
  NAND2X0_LVT U9988 ( .A1(n9065), .A2(n_T_1165[55]), .Y(n8743) );
  NAND2X0_LVT U9989 ( .A1(n2493), .A2(n_T_628[55]), .Y(n8742) );
  NAND2X0_LVT U9990 ( .A1(n9066), .A2(n_T_918[55]), .Y(n8741) );
  NAND4X0_LVT U9991 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .Y(
        io_fpu_fromint_data[55]) );
  AO22X1_LVT U9992 ( .A1(n4022), .A2(n_T_427[696]), .A3(n4036), .A4(
        n_T_427[376]), .Y(n8750) );
  AO22X1_LVT U9993 ( .A1(n4044), .A2(n_T_427[120]), .A3(n4048), .A4(
        n_T_427[759]), .Y(n8749) );
  AO22X1_LVT U9994 ( .A1(n3975), .A2(n_T_427[184]), .A3(n3979), .A4(
        n_T_427[823]), .Y(n8747) );
  AO22X1_LVT U9995 ( .A1(n4023), .A2(n_T_427[951]), .A3(n4031), .A4(
        n_T_427[632]), .Y(n8746) );
  AO22X1_LVT U9996 ( .A1(n3971), .A2(n_T_427[440]), .A3(n3976), .A4(
        n_T_427[568]), .Y(n8745) );
  OR3X1_LVT U9997 ( .A1(n8747), .A2(n8746), .A3(n8745), .Y(n8748) );
  OR3X1_LVT U9998 ( .A1(n8750), .A2(n8749), .A3(n8748), .Y(n8751) );
  NAND2X0_LVT U9999 ( .A1(n4053), .A2(n8751), .Y(n8752) );
  NAND2X0_LVT U10000 ( .A1(n3661), .A2(n_T_427[887]), .Y(n8755) );
  NAND2X0_LVT U10001 ( .A1(n_T_427[504]), .A2(n9052), .Y(n8754) );
  NAND2X0_LVT U10002 ( .A1(n3675), .A2(n_T_427[1143]), .Y(n8756) );
  NAND2X0_LVT U10003 ( .A1(n3758), .A2(n_T_427[1015]), .Y(n8758) );
  NAND2X0_LVT U10004 ( .A1(n3716), .A2(n_T_427[1079]), .Y(n8757) );
  NAND2X0_LVT U10005 ( .A1(n_T_427[1399]), .A2(n3609), .Y(n8759) );
  OA21X1_LVT U10006 ( .A1(n3162), .A2(n3989), .A3(n8759), .Y(n8762) );
  NAND2X0_LVT U10007 ( .A1(n3627), .A2(n_T_427[1463]), .Y(n8761) );
  NAND2X0_LVT U10008 ( .A1(n2998), .A2(n_T_427[1935]), .Y(n8760) );
  AND3X1_LVT U10009 ( .A1(n8762), .A2(n8761), .A3(n8760), .Y(n8765) );
  NAND2X0_LVT U10010 ( .A1(n3745), .A2(n_T_427[248]), .Y(n8764) );
  NAND2X0_LVT U10011 ( .A1(n3647), .A2(n_T_427[56]), .Y(n8763) );
  NAND3X0_LVT U10012 ( .A1(n8765), .A2(n8764), .A3(n8763), .Y(n8775) );
  NAND2X0_LVT U10013 ( .A1(n3689), .A2(n_T_427[1719]), .Y(n8766) );
  OA21X1_LVT U10014 ( .A1(n3472), .A2(n3994), .A3(n8766), .Y(n8769) );
  NAND2X0_LVT U10015 ( .A1(n3999), .A2(n_T_427[1335]), .Y(n8768) );
  NAND2X0_LVT U10016 ( .A1(n4004), .A2(n_T_427[1783]), .Y(n8767) );
  NAND2X0_LVT U10017 ( .A1(n3770), .A2(n_T_427[1527]), .Y(n8770) );
  OA21X1_LVT U10018 ( .A1(n3664), .A2(n3362), .A3(n8770), .Y(n8773) );
  NAND2X0_LVT U10019 ( .A1(n3617), .A2(n_T_427[1591]), .Y(n8772) );
  NAND2X0_LVT U10020 ( .A1(n3642), .A2(n_T_427[1655]), .Y(n8771) );
  OR3X1_LVT U10021 ( .A1(n8776), .A2(n8775), .A3(n8774), .Y(N736) );
  NAND2X0_LVT U10022 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[56]), .Y(n8780)
         );
  NAND2X0_LVT U10023 ( .A1(n9065), .A2(n_T_1165[56]), .Y(n8779) );
  NAND2X0_LVT U10024 ( .A1(n2497), .A2(n_T_628[56]), .Y(n8778) );
  NAND2X0_LVT U10025 ( .A1(n9066), .A2(n_T_918[56]), .Y(n8777) );
  NAND4X0_LVT U10026 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .Y(
        io_fpu_fromint_data[56]) );
  NAND2X0_LVT U10027 ( .A1(n3629), .A2(n_T_427[1464]), .Y(n8783) );
  NAND2X0_LVT U10028 ( .A1(n3992), .A2(n_T_427[1936]), .Y(n8782) );
  NAND3X0_LVT U10029 ( .A1(n8784), .A2(n8783), .A3(n8782), .Y(n8790) );
  NAND2X0_LVT U10030 ( .A1(n3689), .A2(n_T_427[1720]), .Y(n8785) );
  OA21X1_LVT U10031 ( .A1(n3751), .A2(n3473), .A3(n8785), .Y(n8788) );
  NAND2X0_LVT U10032 ( .A1(n3997), .A2(n_T_427[1336]), .Y(n8787) );
  NAND2X0_LVT U10033 ( .A1(n4005), .A2(n_T_427[1784]), .Y(n8786) );
  NAND3X0_LVT U10034 ( .A1(n8788), .A2(n8787), .A3(n8786), .Y(n8789) );
  NAND2X0_LVT U10035 ( .A1(n3770), .A2(n_T_427[1528]), .Y(n8791) );
  OA21X1_LVT U10036 ( .A1(n4009), .A2(n3363), .A3(n8791), .Y(n8794) );
  NAND2X0_LVT U10037 ( .A1(n3616), .A2(n_T_427[1592]), .Y(n8793) );
  NAND2X0_LVT U10038 ( .A1(n3649), .A2(n_T_427[1656]), .Y(n8792) );
  NAND3X0_LVT U10039 ( .A1(n8794), .A2(n8793), .A3(n8792), .Y(n8798) );
  NAND2X0_LVT U10040 ( .A1(n_T_427[1272]), .A2(n3638), .Y(n8796) );
  NAND2X0_LVT U10041 ( .A1(n3674), .A2(n_T_427[1144]), .Y(n8795) );
  NAND2X0_LVT U10042 ( .A1(n3787), .A2(n_T_427[569]), .Y(n8806) );
  NAND2X0_LVT U10043 ( .A1(n3665), .A2(n4478), .Y(n8805) );
  AO22X1_LVT U10044 ( .A1(n4023), .A2(n_T_427[952]), .A3(n3960), .A4(
        n_T_427[505]), .Y(n8802) );
  AO22X1_LVT U10045 ( .A1(n4022), .A2(n_T_427[697]), .A3(n4043), .A4(
        n_T_427[121]), .Y(n8801) );
  AO22X1_LVT U10046 ( .A1(n4035), .A2(n_T_427[633]), .A3(n4027), .A4(
        n_T_427[888]), .Y(n8800) );
  AO22X1_LVT U10047 ( .A1(n4039), .A2(n_T_427[377]), .A3(n4052), .A4(
        n_T_427[57]), .Y(n8799) );
  NOR4X1_LVT U10048 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .Y(n8803) );
  NAND3X0_LVT U10049 ( .A1(n8806), .A2(n8805), .A3(n8804), .Y(n8815) );
  NAND2X0_LVT U10050 ( .A1(n3713), .A2(n_T_427[185]), .Y(n8808) );
  NAND2X0_LVT U10051 ( .A1(n3790), .A2(n_T_427[313]), .Y(n8807) );
  NAND2X0_LVT U10052 ( .A1(n8808), .A2(n8807), .Y(n8814) );
  NAND2X0_LVT U10053 ( .A1(n9058), .A2(n_T_427[249]), .Y(n8809) );
  OA21X1_LVT U10054 ( .A1(n3708), .A2(n3302), .A3(n8809), .Y(n8812) );
  NAND2X0_LVT U10055 ( .A1(n9056), .A2(n_T_427[824]), .Y(n8810) );
  NAND3X0_LVT U10056 ( .A1(n8811), .A2(n8812), .A3(n8810), .Y(n8813) );
  NAND2X0_LVT U10057 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[57]), .Y(n8819)
         );
  NAND2X0_LVT U10058 ( .A1(n9065), .A2(n_T_1165[57]), .Y(n8818) );
  NAND2X0_LVT U10059 ( .A1(n2497), .A2(n_T_628[57]), .Y(n8817) );
  NAND2X0_LVT U10060 ( .A1(n9066), .A2(n_T_918[57]), .Y(n8816) );
  NAND4X0_LVT U10061 ( .A1(n8819), .A2(n8818), .A3(n8817), .A4(n8816), .Y(
        io_fpu_fromint_data[57]) );
  NAND2X0_LVT U10062 ( .A1(n3610), .A2(n_T_427[1401]), .Y(n8820) );
  OA21X1_LVT U10063 ( .A1(n3164), .A2(n2969), .A3(n8820), .Y(n8823) );
  NAND2X0_LVT U10064 ( .A1(n3630), .A2(n_T_427[1465]), .Y(n8822) );
  NAND2X0_LVT U10065 ( .A1(n2882), .A2(n_T_427[1937]), .Y(n8821) );
  NAND2X0_LVT U10066 ( .A1(n3689), .A2(n_T_427[1721]), .Y(n8824) );
  OA21X1_LVT U10067 ( .A1(n3474), .A2(n3994), .A3(n8824), .Y(n8827) );
  NAND2X0_LVT U10068 ( .A1(n3999), .A2(n_T_427[1337]), .Y(n8826) );
  NAND2X0_LVT U10069 ( .A1(n4001), .A2(n_T_427[1785]), .Y(n8825) );
  NAND2X0_LVT U10070 ( .A1(n3769), .A2(n_T_427[1529]), .Y(n8828) );
  NAND2X0_LVT U10071 ( .A1(n3619), .A2(n_T_427[1593]), .Y(n8830) );
  NAND3X0_LVT U10072 ( .A1(n8831), .A2(n8830), .A3(n8829), .Y(n8836) );
  NAND2X0_LVT U10073 ( .A1(n3759), .A2(n_T_427[1017]), .Y(n8832) );
  NAND2X0_LVT U10074 ( .A1(n_T_427[1273]), .A2(n3640), .Y(n8834) );
  NAND2X0_LVT U10075 ( .A1(n3675), .A2(n_T_427[1145]), .Y(n8833) );
  NAND2X0_LVT U10076 ( .A1(n8837), .A2(n_T_427[634]), .Y(n8845) );
  NAND2X0_LVT U10077 ( .A1(n3060), .A2(n4481), .Y(n8844) );
  AO22X1_LVT U10078 ( .A1(n4023), .A2(n_T_427[953]), .A3(n4021), .A4(
        n_T_427[698]), .Y(n8841) );
  AO22X1_LVT U10079 ( .A1(n3971), .A2(n_T_427[442]), .A3(n4036), .A4(
        n_T_427[378]), .Y(n8840) );
  AO22X1_LVT U10080 ( .A1(n3986), .A2(n_T_427[250]), .A3(n4028), .A4(
        n_T_427[889]), .Y(n8839) );
  AO22X1_LVT U10081 ( .A1(n4052), .A2(n_T_427[58]), .A3(n4048), .A4(
        n_T_427[761]), .Y(n8838) );
  NOR4X1_LVT U10082 ( .A1(n8841), .A2(n8840), .A3(n8839), .A4(n8838), .Y(n8842) );
  NAND3X0_LVT U10083 ( .A1(n8845), .A2(n8844), .A3(n8843), .Y(n8851) );
  NAND2X0_LVT U10084 ( .A1(n3788), .A2(n_T_427[570]), .Y(n8847) );
  NAND2X0_LVT U10085 ( .A1(n_T_427[506]), .A2(n9052), .Y(n8846) );
  NAND2X0_LVT U10086 ( .A1(n8847), .A2(n8846), .Y(n8850) );
  NAND2X0_LVT U10087 ( .A1(n_T_427[314]), .A2(n9053), .Y(n8848) );
  NAND2X0_LVT U10088 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[58]), .Y(n8855)
         );
  NAND2X0_LVT U10089 ( .A1(n9065), .A2(n_T_1165[58]), .Y(n8854) );
  NAND2X0_LVT U10090 ( .A1(n2497), .A2(n_T_628[58]), .Y(n8853) );
  NAND2X0_LVT U10091 ( .A1(n9066), .A2(n_T_918[58]), .Y(n8852) );
  NAND4X0_LVT U10092 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .Y(
        io_fpu_fromint_data[58]) );
  NAND2X0_LVT U10093 ( .A1(n3609), .A2(n_T_427[1402]), .Y(n8856) );
  OA21X1_LVT U10094 ( .A1(n3165), .A2(n3988), .A3(n8856), .Y(n8859) );
  NAND2X0_LVT U10095 ( .A1(n3628), .A2(n_T_427[1466]), .Y(n8858) );
  NAND2X0_LVT U10096 ( .A1(n2998), .A2(n_T_427[1938]), .Y(n8857) );
  NAND2X0_LVT U10097 ( .A1(n3689), .A2(n_T_427[1722]), .Y(n8860) );
  OA21X1_LVT U10098 ( .A1(n3166), .A2(n3994), .A3(n8860), .Y(n8863) );
  NAND2X0_LVT U10099 ( .A1(n4000), .A2(n_T_427[1338]), .Y(n8862) );
  NAND2X0_LVT U10100 ( .A1(n2092), .A2(n_T_427[1786]), .Y(n8861) );
  NAND2X0_LVT U10101 ( .A1(n3769), .A2(n_T_427[1530]), .Y(n8864) );
  OA21X1_LVT U10102 ( .A1(n3663), .A2(n3367), .A3(n8864), .Y(n8867) );
  NAND2X0_LVT U10103 ( .A1(n3617), .A2(n_T_427[1594]), .Y(n8866) );
  NAND2X0_LVT U10104 ( .A1(n3643), .A2(n_T_427[1658]), .Y(n8865) );
  NAND3X0_LVT U10105 ( .A1(n8867), .A2(n8866), .A3(n8865), .Y(n8872) );
  NAND2X0_LVT U10106 ( .A1(n3757), .A2(n_T_427[1018]), .Y(n8868) );
  NAND2X0_LVT U10107 ( .A1(n3637), .A2(n_T_427[1274]), .Y(n8870) );
  NAND2X0_LVT U10108 ( .A1(n_T_427[1146]), .A2(n3669), .Y(n8869) );
  NAND2X0_LVT U10109 ( .A1(n8873), .A2(n_T_427[954]), .Y(n8881) );
  NAND2X0_LVT U10110 ( .A1(n3060), .A2(n4484), .Y(n8880) );
  AO22X1_LVT U10111 ( .A1(n3971), .A2(n_T_427[443]), .A3(n4021), .A4(
        n_T_427[699]), .Y(n8877) );
  AO22X1_LVT U10112 ( .A1(n2858), .A2(n_T_427[187]), .A3(n4048), .A4(
        n_T_427[762]), .Y(n8876) );
  AO22X1_LVT U10113 ( .A1(n3963), .A2(n_T_427[507]), .A3(n4031), .A4(
        n_T_427[635]), .Y(n8875) );
  AO22X1_LVT U10114 ( .A1(n4041), .A2(n_T_427[123]), .A3(n4036), .A4(
        n_T_427[379]), .Y(n8874) );
  NOR4X1_LVT U10115 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .Y(n8878) );
  NAND3X0_LVT U10116 ( .A1(n8881), .A2(n8880), .A3(n8879), .Y(n8889) );
  NAND2X0_LVT U10117 ( .A1(n3787), .A2(n_T_427[571]), .Y(n8883) );
  NAND2X0_LVT U10118 ( .A1(n3661), .A2(n_T_427[890]), .Y(n8882) );
  NAND2X0_LVT U10119 ( .A1(n8883), .A2(n8882), .Y(n8888) );
  NAND2X0_LVT U10120 ( .A1(n_T_427[251]), .A2(n9058), .Y(n8885) );
  AND2X1_LVT U10121 ( .A1(n8885), .A2(n8884), .Y(n8887) );
  NAND2X0_LVT U10122 ( .A1(n_T_427[315]), .A2(n3790), .Y(n8886) );
  NAND2X0_LVT U10123 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[59]), .Y(n8893)
         );
  NAND2X0_LVT U10124 ( .A1(n9065), .A2(n_T_1165[59]), .Y(n8892) );
  NAND2X0_LVT U10125 ( .A1(n2497), .A2(n_T_628[59]), .Y(n8891) );
  NAND2X0_LVT U10126 ( .A1(n9066), .A2(n_T_918[59]), .Y(n8890) );
  NAND4X0_LVT U10127 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .Y(
        io_fpu_fromint_data[59]) );
  NAND2X0_LVT U10128 ( .A1(n3610), .A2(n_T_427[1403]), .Y(n8894) );
  NAND2X0_LVT U10129 ( .A1(n3628), .A2(n_T_427[1467]), .Y(n8896) );
  NAND2X0_LVT U10130 ( .A1(n2882), .A2(n_T_427[1939]), .Y(n8895) );
  NAND2X0_LVT U10131 ( .A1(n3600), .A2(n_T_427[827]), .Y(n8898) );
  NAND2X0_LVT U10132 ( .A1(n3707), .A2(n_T_427[124]), .Y(n8897) );
  NAND3X0_LVT U10133 ( .A1(n8899), .A2(n8898), .A3(n8897), .Y(n8925) );
  NAND2X0_LVT U10134 ( .A1(n3786), .A2(n_T_427[572]), .Y(n8908) );
  NAND2X0_LVT U10135 ( .A1(n3060), .A2(n4487), .Y(n8907) );
  AO22X1_LVT U10136 ( .A1(n3960), .A2(n_T_427[508]), .A3(n4036), .A4(
        n_T_427[380]), .Y(n8904) );
  AO22X1_LVT U10137 ( .A1(n3970), .A2(n_T_427[444]), .A3(n3964), .A4(
        n_T_427[316]), .Y(n8903) );
  OR3X1_LVT U10138 ( .A1(n8904), .A2(n8903), .A3(n8902), .Y(n8905) );
  NAND2X0_LVT U10139 ( .A1(n4053), .A2(n8905), .Y(n8906) );
  NAND2X0_LVT U10140 ( .A1(n8991), .A2(n_T_427[891]), .Y(n8909) );
  NAND2X0_LVT U10141 ( .A1(n_T_427[1019]), .A2(n3755), .Y(n8911) );
  OA21X1_LVT U10142 ( .A1(n4011), .A2(n3303), .A3(n8911), .Y(n8914) );
  NAND2X0_LVT U10143 ( .A1(n_T_427[1275]), .A2(n3638), .Y(n8913) );
  NAND2X0_LVT U10144 ( .A1(n3668), .A2(n_T_427[1147]), .Y(n8912) );
  NAND2X0_LVT U10145 ( .A1(n3689), .A2(n_T_427[1723]), .Y(n8915) );
  OA21X1_LVT U10146 ( .A1(n3410), .A2(n3747), .A3(n8915), .Y(n8918) );
  NAND2X0_LVT U10147 ( .A1(n3996), .A2(n_T_427[1339]), .Y(n8917) );
  NAND2X0_LVT U10148 ( .A1(n4002), .A2(n_T_427[1787]), .Y(n8916) );
  NAND2X0_LVT U10149 ( .A1(n3769), .A2(n_T_427[1531]), .Y(n8919) );
  OA21X1_LVT U10150 ( .A1(n4009), .A2(n3304), .A3(n8919), .Y(n8922) );
  NAND2X0_LVT U10151 ( .A1(n3618), .A2(n_T_427[1595]), .Y(n8921) );
  NAND2X0_LVT U10152 ( .A1(n3649), .A2(n_T_427[1659]), .Y(n8920) );
  OR3X1_LVT U10153 ( .A1(n8924), .A2(n8925), .A3(n8923), .Y(N740) );
  NAND2X0_LVT U10154 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[60]), .Y(n8929)
         );
  NAND2X0_LVT U10155 ( .A1(n9065), .A2(n_T_1165[60]), .Y(n8928) );
  NAND2X0_LVT U10156 ( .A1(n2493), .A2(n_T_628[60]), .Y(n8927) );
  NAND2X0_LVT U10157 ( .A1(n9066), .A2(n_T_918[60]), .Y(n8926) );
  NAND4X0_LVT U10158 ( .A1(n8929), .A2(n8928), .A3(n8927), .A4(n8926), .Y(
        io_fpu_fromint_data[60]) );
  NAND2X0_LVT U10159 ( .A1(n3789), .A2(n_T_427[317]), .Y(n8930) );
  OA21X1_LVT U10160 ( .A1(n3691), .A2(n3280), .A3(n8930), .Y(n8942) );
  AO22X1_LVT U10161 ( .A1(n4023), .A2(n_T_427[956]), .A3(n3976), .A4(
        n_T_427[573]), .Y(n8936) );
  AO22X1_LVT U10162 ( .A1(n3968), .A2(n_T_427[445]), .A3(n4020), .A4(
        n_T_427[701]), .Y(n8935) );
  AO22X1_LVT U10163 ( .A1(n2858), .A2(n_T_427[189]), .A3(n3979), .A4(
        n_T_427[828]), .Y(n8934) );
  AO22X1_LVT U10164 ( .A1(n4035), .A2(n_T_427[637]), .A3(n4027), .A4(
        n_T_427[892]), .Y(n8933) );
  NOR4X1_LVT U10165 ( .A1(n8936), .A2(n8935), .A3(n8934), .A4(n8933), .Y(n8938) );
  NAND2X0_LVT U10166 ( .A1(n2982), .A2(n4490), .Y(n8937) );
  OA21X1_LVT U10167 ( .A1(n8938), .A2(n3612), .A3(n8937), .Y(n8941) );
  NAND2X0_LVT U10168 ( .A1(n8939), .A2(n_T_427[381]), .Y(n8940) );
  NAND2X0_LVT U10169 ( .A1(n3745), .A2(n_T_427[253]), .Y(n8943) );
  NAND2X0_LVT U10170 ( .A1(n_T_427[509]), .A2(n3614), .Y(n8946) );
  NAND2X0_LVT U10171 ( .A1(n8944), .A2(n_T_427[61]), .Y(n8945) );
  NAND2X0_LVT U10172 ( .A1(n3605), .A2(n_T_427[1404]), .Y(n8947) );
  OA21X1_LVT U10173 ( .A1(n3167), .A2(n3987), .A3(n8947), .Y(n8950) );
  NAND2X0_LVT U10174 ( .A1(n2966), .A2(n_T_427[1468]), .Y(n8949) );
  NAND2X0_LVT U10175 ( .A1(n3991), .A2(n_T_427[1940]), .Y(n8948) );
  NAND2X0_LVT U10176 ( .A1(n3657), .A2(n_T_427[1724]), .Y(n8951) );
  OA21X1_LVT U10177 ( .A1(n3168), .A2(n3751), .A3(n8951), .Y(n8954) );
  NAND2X0_LVT U10178 ( .A1(n2094), .A2(n_T_427[1340]), .Y(n8953) );
  NAND2X0_LVT U10179 ( .A1(n4005), .A2(n_T_427[1788]), .Y(n8952) );
  NAND2X0_LVT U10180 ( .A1(n3770), .A2(n_T_427[1532]), .Y(n8955) );
  NAND2X0_LVT U10181 ( .A1(n3615), .A2(n_T_427[1596]), .Y(n8957) );
  NAND2X0_LVT U10182 ( .A1(n_T_427[1660]), .A2(n3650), .Y(n8956) );
  NAND2X0_LVT U10183 ( .A1(n3712), .A2(n_T_427[1020]), .Y(n8959) );
  OA21X1_LVT U10184 ( .A1(n4011), .A2(n3281), .A3(n8959), .Y(n8962) );
  NAND2X0_LVT U10185 ( .A1(n_T_427[1276]), .A2(n3638), .Y(n8961) );
  NAND2X0_LVT U10186 ( .A1(n3667), .A2(n_T_427[1148]), .Y(n8960) );
  NAND2X0_LVT U10187 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[61]), .Y(n8966)
         );
  NAND2X0_LVT U10188 ( .A1(n9065), .A2(n_T_1165[61]), .Y(n8965) );
  NAND2X0_LVT U10189 ( .A1(n2493), .A2(n_T_628[61]), .Y(n8964) );
  NAND2X0_LVT U10190 ( .A1(n9066), .A2(n_T_918[61]), .Y(n8963) );
  NAND4X0_LVT U10191 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .Y(
        io_fpu_fromint_data[61]) );
  NAND2X0_LVT U10192 ( .A1(n_T_427[1405]), .A2(n3608), .Y(n8967) );
  OA21X1_LVT U10193 ( .A1(n3169), .A2(n3989), .A3(n8967), .Y(n8970) );
  NAND2X0_LVT U10194 ( .A1(n3626), .A2(n_T_427[1469]), .Y(n8969) );
  NAND2X0_LVT U10195 ( .A1(n2986), .A2(n_T_427[1941]), .Y(n8968) );
  NAND2X0_LVT U10196 ( .A1(n3657), .A2(n_T_427[1725]), .Y(n8971) );
  OA21X1_LVT U10197 ( .A1(n3411), .A2(n3751), .A3(n8971), .Y(n8974) );
  NAND2X0_LVT U10198 ( .A1(n3998), .A2(n_T_427[1341]), .Y(n8973) );
  NAND2X0_LVT U10199 ( .A1(n4003), .A2(n_T_427[1789]), .Y(n8972) );
  NAND2X0_LVT U10200 ( .A1(n3770), .A2(n_T_427[1533]), .Y(n8975) );
  NAND2X0_LVT U10201 ( .A1(n3620), .A2(n_T_427[1597]), .Y(n8977) );
  NAND2X0_LVT U10202 ( .A1(n3650), .A2(n_T_427[1661]), .Y(n8976) );
  NAND2X0_LVT U10203 ( .A1(n3756), .A2(n_T_427[1021]), .Y(n8979) );
  NAND2X0_LVT U10204 ( .A1(n_T_427[318]), .A2(n3790), .Y(n8990) );
  NAND2X0_LVT U10205 ( .A1(n3665), .A2(n4493), .Y(n8989) );
  AO22X1_LVT U10206 ( .A1(n4023), .A2(n_T_427[957]), .A3(n3976), .A4(
        n_T_427[574]), .Y(n8986) );
  AO22X1_LVT U10207 ( .A1(n3979), .A2(n_T_427[829]), .A3(n4052), .A4(
        n_T_427[62]), .Y(n8985) );
  AO22X1_LVT U10208 ( .A1(n4034), .A2(n_T_427[638]), .A3(n3983), .A4(
        n_T_427[254]), .Y(n8984) );
  AO22X1_LVT U10209 ( .A1(n4039), .A2(n_T_427[382]), .A3(n4048), .A4(
        n_T_427[765]), .Y(n8983) );
  NOR4X1_LVT U10210 ( .A1(n8986), .A2(n8985), .A3(n8984), .A4(n8983), .Y(n8987) );
  NAND2X0_LVT U10211 ( .A1(n8991), .A2(n_T_427[893]), .Y(n8993) );
  NAND2X0_LVT U10212 ( .A1(n_T_427[510]), .A2(n9052), .Y(n8992) );
  NAND2X0_LVT U10213 ( .A1(n8994), .A2(n_T_427[126]), .Y(n8995) );
  OA21X1_LVT U10214 ( .A1(n3478), .A2(n8996), .A3(n8995), .Y(n8999) );
  NAND2X0_LVT U10215 ( .A1(n3713), .A2(n_T_427[190]), .Y(n8997) );
  NAND2X0_LVT U10216 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[62]), .Y(n9003)
         );
  NAND2X0_LVT U10217 ( .A1(n9065), .A2(n_T_1165[62]), .Y(n9002) );
  NAND2X0_LVT U10218 ( .A1(n2493), .A2(n_T_628[62]), .Y(n9001) );
  NAND2X0_LVT U10219 ( .A1(n9066), .A2(n_T_918[62]), .Y(n9000) );
  NAND4X0_LVT U10220 ( .A1(n9003), .A2(n9002), .A3(n9001), .A4(n9000), .Y(
        io_fpu_fromint_data[62]) );
  NAND2X0_LVT U10221 ( .A1(n3604), .A2(n_T_427[1406]), .Y(n9005) );
  NAND2X0_LVT U10222 ( .A1(n3626), .A2(n_T_427[1470]), .Y(n9010) );
  NAND2X0_LVT U10223 ( .A1(n3992), .A2(n_T_427[1942]), .Y(n9009) );
  NAND2X0_LVT U10224 ( .A1(n2922), .A2(n_T_427[1726]), .Y(n9013) );
  OA21X1_LVT U10225 ( .A1(n3171), .A2(n3747), .A3(n9013), .Y(n9019) );
  NAND2X0_LVT U10226 ( .A1(n3997), .A2(n_T_427[1342]), .Y(n9018) );
  NAND2X0_LVT U10227 ( .A1(n4003), .A2(n_T_427[1790]), .Y(n9017) );
  NAND2X0_LVT U10228 ( .A1(n3769), .A2(n_T_427[1534]), .Y(n9020) );
  OA21X1_LVT U10229 ( .A1(n3663), .A2(n3308), .A3(n9020), .Y(n9025) );
  NAND2X0_LVT U10230 ( .A1(n3620), .A2(n_T_427[1598]), .Y(n9024) );
  NAND3X0_LVT U10231 ( .A1(n9025), .A2(n9024), .A3(n9023), .Y(n9034) );
  NAND2X0_LVT U10232 ( .A1(n_T_427[1022]), .A2(n3761), .Y(n9027) );
  NAND2X0_LVT U10233 ( .A1(n3639), .A2(n_T_427[1278]), .Y(n9032) );
  NAND2X0_LVT U10234 ( .A1(n3674), .A2(n_T_427[1150]), .Y(n9031) );
  NAND2X0_LVT U10235 ( .A1(n3787), .A2(n_T_427[575]), .Y(n9051) );
  NAND2X0_LVT U10236 ( .A1(n3665), .A2(n4496), .Y(n9050) );
  AO22X1_LVT U10237 ( .A1(n4025), .A2(n_T_427[958]), .A3(n4018), .A4(
        n_T_427[703]), .Y(n9046) );
  AO22X1_LVT U10238 ( .A1(n4031), .A2(n_T_427[639]), .A3(n4028), .A4(
        n_T_427[894]), .Y(n9045) );
  AO22X1_LVT U10239 ( .A1(n4044), .A2(n_T_427[127]), .A3(n4038), .A4(
        n_T_427[383]), .Y(n9044) );
  AO22X1_LVT U10240 ( .A1(n4052), .A2(n_T_427[63]), .A3(n4045), .A4(
        n_T_427[766]), .Y(n9043) );
  NOR4X1_LVT U10241 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .Y(n9048) );
  NAND3X0_LVT U10242 ( .A1(n9051), .A2(n9050), .A3(n9049), .Y(n9063) );
  NAND2X0_LVT U10243 ( .A1(n_T_427[511]), .A2(n9052), .Y(n9055) );
  NAND2X0_LVT U10244 ( .A1(n3790), .A2(n_T_427[319]), .Y(n9054) );
  NAND2X0_LVT U10245 ( .A1(n9055), .A2(n9054), .Y(n9062) );
  NAND2X0_LVT U10246 ( .A1(n9056), .A2(n_T_427[830]), .Y(n9057) );
  NAND2X0_LVT U10247 ( .A1(n_T_427[255]), .A2(n3624), .Y(n9061) );
  NAND2X0_LVT U10248 ( .A1(n3714), .A2(n_T_427[191]), .Y(n9060) );
  NAND2X0_LVT U10249 ( .A1(n9064), .A2(io_fpu_dmem_resp_data[63]), .Y(n9070)
         );
  NAND2X0_LVT U10250 ( .A1(n9065), .A2(n_T_1165[63]), .Y(n9069) );
  NAND2X0_LVT U10251 ( .A1(n2493), .A2(n_T_628[63]), .Y(n9068) );
  NAND2X0_LVT U10252 ( .A1(n9066), .A2(n_T_918[63]), .Y(n9067) );
  NAND4X0_LVT U10253 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .Y(
        io_fpu_fromint_data[63]) );
  MUX21X1_LVT U10254 ( .A1(n2553), .A2(io_fpu_inst[14]), .S0(io_fpu_inst[13]), 
        .Y(n9072) );
  NAND2X0_LVT U10255 ( .A1(n9107), .A2(n1891), .Y(n9071) );
  NAND2X0_LVT U10256 ( .A1(n9071), .A2(n9413), .Y(n9078) );
  AO21X1_LVT U10257 ( .A1(n9073), .A2(n9072), .A3(n9078), .Y(n9074) );
  AND2X1_LVT U10258 ( .A1(n2677), .A2(n9074), .Y(n1589) );
  NAND2X0_LVT U10259 ( .A1(n9087), .A2(io_fpu_inst[13]), .Y(n9085) );
  NAND2X0_LVT U10260 ( .A1(n9078), .A2(io_fpu_inst[13]), .Y(n9082) );
  NAND3X0_LVT U10261 ( .A1(n9082), .A2(n9081), .A3(n9080), .Y(n9083) );
  NAND2X0_LVT U10262 ( .A1(n2677), .A2(n9083), .Y(n9084) );
  NAND3X0_LVT U10263 ( .A1(n9084), .A2(n9228), .A3(n9085), .Y(N282) );
  NAND2X0_LVT U10264 ( .A1(n3079), .A2(n2618), .Y(n9086) );
  NAND2X0_LVT U10265 ( .A1(n9086), .A2(n9087), .Y(n9093) );
  NAND3X0_LVT U10266 ( .A1(n9093), .A2(n9233), .A3(n9229), .Y(N283) );
  INVX1_LVT U10267 ( .A(bpu_io_debug_if), .Y(n9242) );
  AO22X1_LVT U10268 ( .A1(io_fpu_inst[6]), .A2(io_fpu_inst[3]), .A3(n9097), 
        .A4(n1863), .Y(n9098) );
  NAND2X0_LVT U10269 ( .A1(n9116), .A2(n9098), .Y(n9100) );
  AO21X1_LVT U10270 ( .A1(n9103), .A2(io_fpu_fromint_data[40]), .A3(n9102), 
        .Y(alu_io_in1[40]) );
  AO21X1_LVT U10271 ( .A1(n9103), .A2(io_fpu_fromint_data[42]), .A3(n9102), 
        .Y(alu_io_in1[42]) );
  AO21X1_LVT U10272 ( .A1(n9103), .A2(io_fpu_fromint_data[44]), .A3(n9102), 
        .Y(alu_io_in1[44]) );
  AO21X1_LVT U10273 ( .A1(n9103), .A2(io_fpu_fromint_data[45]), .A3(n9102), 
        .Y(alu_io_in1[45]) );
  AO21X1_LVT U10274 ( .A1(n9103), .A2(io_fpu_fromint_data[46]), .A3(n9102), 
        .Y(alu_io_in1[46]) );
  AO21X1_LVT U10275 ( .A1(n9103), .A2(io_fpu_fromint_data[47]), .A3(n9102), 
        .Y(alu_io_in1[47]) );
  AO21X1_LVT U10276 ( .A1(n9103), .A2(io_fpu_fromint_data[48]), .A3(n9102), 
        .Y(alu_io_in1[48]) );
  AO21X1_LVT U10277 ( .A1(n9103), .A2(io_fpu_fromint_data[50]), .A3(n9102), 
        .Y(alu_io_in1[50]) );
  AO21X1_LVT U10278 ( .A1(n9103), .A2(io_fpu_fromint_data[52]), .A3(n9102), 
        .Y(alu_io_in1[52]) );
  AO21X1_LVT U10279 ( .A1(n9103), .A2(io_fpu_fromint_data[53]), .A3(n9102), 
        .Y(alu_io_in1[53]) );
  AO21X1_LVT U10280 ( .A1(n9103), .A2(io_fpu_fromint_data[54]), .A3(n9102), 
        .Y(alu_io_in1[54]) );
  AO21X1_LVT U10281 ( .A1(n9103), .A2(io_fpu_fromint_data[56]), .A3(n9102), 
        .Y(alu_io_in1[56]) );
  AO21X1_LVT U10282 ( .A1(n9103), .A2(io_fpu_fromint_data[57]), .A3(n9102), 
        .Y(alu_io_in1[57]) );
  AO21X1_LVT U10283 ( .A1(n9103), .A2(io_fpu_fromint_data[58]), .A3(n9102), 
        .Y(alu_io_in1[58]) );
  AO21X1_LVT U10284 ( .A1(n9103), .A2(io_fpu_fromint_data[59]), .A3(n9102), 
        .Y(alu_io_in1[59]) );
  AO21X1_LVT U10285 ( .A1(n9103), .A2(io_fpu_fromint_data[60]), .A3(n9102), 
        .Y(alu_io_in1[60]) );
  AO21X1_LVT U10286 ( .A1(n9103), .A2(io_fpu_fromint_data[61]), .A3(n9102), 
        .Y(alu_io_in1[61]) );
  AO21X1_LVT U10287 ( .A1(n9103), .A2(io_fpu_fromint_data[62]), .A3(n9102), 
        .Y(alu_io_in1[62]) );
  MUX21X1_LVT U10288 ( .A1(n9105), .A2(n1867), .S0(n1863), .Y(n9106) );
  AO21X1_LVT U10289 ( .A1(n9108), .A2(n9107), .A3(n9106), .Y(
        id_ctrl_sel_imm[2]) );
  NAND2X0_LVT U10290 ( .A1(n9110), .A2(io_fpu_inst[2]), .Y(n9114) );
  NAND2X0_LVT U10291 ( .A1(n9116), .A2(n9115), .Y(n9117) );
  NAND2X0_LVT U10292 ( .A1(n9117), .A2(n9430), .Y(n9119) );
  AND3X1_LVT U10293 ( .A1(n9119), .A2(n9118), .A3(n9244), .Y(N274) );
  AND2X1_LVT U10294 ( .A1(ex_ctrl_sel_alu2[1]), .A2(ex_ctrl_sel_alu2[0]), .Y(
        n9179) );
  NAND3X0_LVT U10295 ( .A1(n546), .A2(ex_ctrl_sel_imm[0]), .A3(
        ex_ctrl_sel_imm[2]), .Y(n9173) );
  AND2X1_LVT U10296 ( .A1(n9120), .A2(n9227), .Y(n9130) );
  AOI22X1_LVT U10297 ( .A1(n9144), .A2(n_T_648[3]), .A3(
        io_fpu_dmem_resp_data[0]), .A4(n9130), .Y(n9129) );
  NAND3X0_LVT U10298 ( .A1(n546), .A2(ex_ctrl_sel_imm[2]), .A3(n_T_642[0]), 
        .Y(n9121) );
  NAND2X0_LVT U10299 ( .A1(n3231), .A2(n546), .Y(n9172) );
  OA22X1_LVT U10300 ( .A1(n9121), .A2(n9201), .A3(n592), .A4(n9163), .Y(n9122)
         );
  OR2X1_LVT U10301 ( .A1(ex_ctrl_sel_imm[0]), .A2(n9122), .Y(n9128) );
  NAND3X0_LVT U10302 ( .A1(n9125), .A2(n9124), .A3(n9123), .Y(n9126) );
  NAND2X0_LVT U10303 ( .A1(n9227), .A2(n9126), .Y(n9127) );
  NAND3X0_LVT U10304 ( .A1(n9129), .A2(n9128), .A3(n9127), .Y(alu_io_in2[0])
         );
  OR2X1_LVT U10305 ( .A1(ex_ctrl_sel_imm[0]), .A2(n9178), .Y(n9200) );
  AND2X1_LVT U10306 ( .A1(n9199), .A2(n9172), .Y(n9158) );
  NAND2X0_LVT U10307 ( .A1(n9158), .A2(n_T_642[1]), .Y(n9141) );
  NAND2X0_LVT U10308 ( .A1(io_fpu_dmem_resp_data[1]), .A2(n9130), .Y(n9134) );
  NAND2X0_LVT U10309 ( .A1(ex_ctrl_sel_alu2[0]), .A2(n3278), .Y(n9142) );
  OR2X1_LVT U10310 ( .A1(n3215), .A2(n9142), .Y(n9131) );
  OA21X1_LVT U10311 ( .A1(n591), .A2(n9163), .A3(n9131), .Y(n9133) );
  NAND2X0_LVT U10312 ( .A1(n_T_648[4]), .A2(n9144), .Y(n9132) );
  AND3X1_LVT U10313 ( .A1(n9134), .A2(n9133), .A3(n9132), .Y(n9140) );
  NAND3X0_LVT U10314 ( .A1(n9137), .A2(n9136), .A3(n9135), .Y(n9138) );
  NAND2X0_LVT U10315 ( .A1(n9227), .A2(n9138), .Y(n9139) );
  NAND3X0_LVT U10316 ( .A1(n9141), .A2(n9140), .A3(n9139), .Y(alu_io_in2[1])
         );
  NAND2X0_LVT U10317 ( .A1(n_T_642[2]), .A2(n9158), .Y(n9154) );
  OR2X1_LVT U10318 ( .A1(ex_reg_rvc), .A2(n9142), .Y(n9143) );
  OA21X1_LVT U10319 ( .A1(n590), .A2(n9163), .A3(n9143), .Y(n9147) );
  NAND3X0_LVT U10320 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[2]), .A3(n9227), 
        .Y(n9146) );
  NAND2X0_LVT U10321 ( .A1(n9144), .A2(n_T_648[5]), .Y(n9145) );
  AND3X1_LVT U10322 ( .A1(n9147), .A2(n9146), .A3(n9145), .Y(n9153) );
  NAND3X0_LVT U10323 ( .A1(n9150), .A2(n9149), .A3(n9148), .Y(n9151) );
  NAND2X0_LVT U10324 ( .A1(n9227), .A2(n9151), .Y(n9152) );
  NAND3X0_LVT U10325 ( .A1(n9154), .A2(n9153), .A3(n9152), .Y(alu_io_in2[2])
         );
  NAND2X0_LVT U10326 ( .A1(n_T_642[4]), .A2(n9158), .Y(n9169) );
  NAND3X0_LVT U10327 ( .A1(n9161), .A2(n9160), .A3(n9159), .Y(n9162) );
  NAND2X0_LVT U10328 ( .A1(n9227), .A2(n9162), .Y(n9168) );
  OA22X1_LVT U10329 ( .A1(n160), .A2(n9164), .A3(n588), .A4(n9163), .Y(n9167)
         );
  NAND3X0_LVT U10330 ( .A1(n9165), .A2(io_fpu_dmem_resp_data[4]), .A3(n9227), 
        .Y(n9166) );
  NAND4X0_LVT U10331 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .Y(
        alu_io_in2[4]) );
  AO22X1_LVT U10332 ( .A1(n_T_642[5]), .A2(n9199), .A3(n_T_702[5]), .A4(n9227), 
        .Y(alu_io_in2[5]) );
  AO22X1_LVT U10333 ( .A1(n_T_642[6]), .A2(n9199), .A3(n_T_702[6]), .A4(n9227), 
        .Y(alu_io_in2[6]) );
  AO22X1_LVT U10334 ( .A1(n_T_642[7]), .A2(n9199), .A3(n_T_702[7]), .A4(n9227), 
        .Y(alu_io_in2[7]) );
  AO22X1_LVT U10335 ( .A1(n_T_642[8]), .A2(n9199), .A3(n_T_702[8]), .A4(n9227), 
        .Y(alu_io_in2[8]) );
  AO22X1_LVT U10336 ( .A1(n_T_642[9]), .A2(n9199), .A3(n_T_702[9]), .A4(n9227), 
        .Y(alu_io_in2[9]) );
  AO22X1_LVT U10337 ( .A1(n_T_642[10]), .A2(n9199), .A3(n_T_702[10]), .A4(
        n9227), .Y(alu_io_in2[10]) );
  NAND2X0_LVT U10338 ( .A1(n9227), .A2(n_T_702[11]), .Y(n9177) );
  AND2X1_LVT U10339 ( .A1(io_dmem_req_bits_tag[1]), .A2(ex_ctrl_sel_imm[0]), 
        .Y(n9170) );
  MUX21X1_LVT U10340 ( .A1(n_T_642[0]), .A2(n9170), .S0(n546), .Y(n9171) );
  NAND3X0_LVT U10341 ( .A1(n9199), .A2(n3231), .A3(n9171), .Y(n9176) );
  NAND2X0_LVT U10342 ( .A1(n9178), .A2(n9226), .Y(n9197) );
  AO21X1_LVT U10343 ( .A1(n9174), .A2(ex_ctrl_sel_imm[0]), .A3(n9197), .Y(
        n9175) );
  NAND3X0_LVT U10344 ( .A1(n9177), .A2(n9176), .A3(n9175), .Y(alu_io_in2[11])
         );
  NAND2X0_LVT U10345 ( .A1(n9227), .A2(n_T_702[12]), .Y(n9182) );
  AND2X1_LVT U10346 ( .A1(n9180), .A2(n9179), .Y(n9195) );
  NAND2X0_LVT U10347 ( .A1(n9195), .A2(n_T_648[0]), .Y(n9181) );
  NAND3X0_LVT U10348 ( .A1(n9182), .A2(n9197), .A3(n9181), .Y(alu_io_in2[12])
         );
  NAND2X0_LVT U10349 ( .A1(n9227), .A2(n_T_702[13]), .Y(n9184) );
  NAND2X0_LVT U10350 ( .A1(n9195), .A2(n_T_648[1]), .Y(n9183) );
  NAND3X0_LVT U10351 ( .A1(n9184), .A2(n9197), .A3(n9183), .Y(alu_io_in2[13])
         );
  NAND2X0_LVT U10352 ( .A1(n9227), .A2(n_T_702[14]), .Y(n9186) );
  NAND2X0_LVT U10353 ( .A1(n9195), .A2(n_T_648[2]), .Y(n9185) );
  NAND3X0_LVT U10354 ( .A1(n9186), .A2(n9197), .A3(n9185), .Y(alu_io_in2[14])
         );
  NAND2X0_LVT U10355 ( .A1(n9227), .A2(n_T_702[15]), .Y(n9188) );
  NAND2X0_LVT U10356 ( .A1(n9195), .A2(n_T_648[3]), .Y(n9187) );
  NAND3X0_LVT U10357 ( .A1(n9188), .A2(n9197), .A3(n9187), .Y(alu_io_in2[15])
         );
  NAND2X0_LVT U10358 ( .A1(n9227), .A2(n_T_702[16]), .Y(n9190) );
  NAND2X0_LVT U10359 ( .A1(n9195), .A2(n_T_648[4]), .Y(n9189) );
  NAND3X0_LVT U10360 ( .A1(n9190), .A2(n9197), .A3(n9189), .Y(alu_io_in2[16])
         );
  NAND2X0_LVT U10361 ( .A1(n9227), .A2(n_T_702[17]), .Y(n9192) );
  NAND2X0_LVT U10362 ( .A1(n9195), .A2(n_T_648[5]), .Y(n9191) );
  NAND3X0_LVT U10363 ( .A1(n9192), .A2(n9197), .A3(n9191), .Y(alu_io_in2[17])
         );
  NAND2X0_LVT U10364 ( .A1(n9227), .A2(n_T_702[18]), .Y(n9194) );
  NAND2X0_LVT U10365 ( .A1(n9195), .A2(n_T_648[6]), .Y(n9193) );
  NAND3X0_LVT U10366 ( .A1(n9194), .A2(n9197), .A3(n9193), .Y(alu_io_in2[18])
         );
  NAND2X0_LVT U10367 ( .A1(n9227), .A2(n_T_702[19]), .Y(n9198) );
  NAND2X0_LVT U10368 ( .A1(n9195), .A2(n_T_648[7]), .Y(n9196) );
  NAND3X0_LVT U10369 ( .A1(n9198), .A2(n9197), .A3(n9196), .Y(alu_io_in2[19])
         );
  NAND2X0_LVT U10370 ( .A1(n9227), .A2(n_T_702[20]), .Y(n9203) );
  NAND2X0_LVT U10371 ( .A1(n9199), .A2(ex_reg_inst_31_), .Y(n9224) );
  NAND2X0_LVT U10372 ( .A1(n9222), .A2(n_T_642[0]), .Y(n9202) );
  NAND3X0_LVT U10373 ( .A1(n9203), .A2(n9224), .A3(n9202), .Y(alu_io_in2[20])
         );
  NAND2X0_LVT U10374 ( .A1(n9227), .A2(n_T_702[21]), .Y(n9205) );
  NAND2X0_LVT U10375 ( .A1(n9222), .A2(n_T_642[1]), .Y(n9204) );
  NAND3X0_LVT U10376 ( .A1(n9205), .A2(n9224), .A3(n9204), .Y(alu_io_in2[21])
         );
  NAND2X0_LVT U10377 ( .A1(n9227), .A2(n_T_702[22]), .Y(n9207) );
  NAND2X0_LVT U10378 ( .A1(n9222), .A2(n_T_642[2]), .Y(n9206) );
  NAND3X0_LVT U10379 ( .A1(n9207), .A2(n9224), .A3(n9206), .Y(alu_io_in2[22])
         );
  NAND2X0_LVT U10380 ( .A1(n9227), .A2(n_T_702[23]), .Y(n9209) );
  NAND2X0_LVT U10381 ( .A1(n9222), .A2(n_T_642[3]), .Y(n9208) );
  NAND3X0_LVT U10382 ( .A1(n9209), .A2(n9224), .A3(n9208), .Y(alu_io_in2[23])
         );
  NAND2X0_LVT U10383 ( .A1(n9227), .A2(n_T_702[24]), .Y(n9211) );
  NAND2X0_LVT U10384 ( .A1(n9222), .A2(n_T_642[4]), .Y(n9210) );
  NAND3X0_LVT U10385 ( .A1(n9211), .A2(n9224), .A3(n9210), .Y(alu_io_in2[24])
         );
  NAND2X0_LVT U10386 ( .A1(n9227), .A2(n_T_702[25]), .Y(n9213) );
  NAND2X0_LVT U10387 ( .A1(n9222), .A2(n_T_642[5]), .Y(n9212) );
  NAND3X0_LVT U10388 ( .A1(n9213), .A2(n9224), .A3(n9212), .Y(alu_io_in2[25])
         );
  NAND2X0_LVT U10389 ( .A1(n9227), .A2(n_T_702[26]), .Y(n9215) );
  NAND2X0_LVT U10390 ( .A1(n9222), .A2(n_T_642[6]), .Y(n9214) );
  NAND3X0_LVT U10391 ( .A1(n9215), .A2(n9224), .A3(n9214), .Y(alu_io_in2[26])
         );
  NAND2X0_LVT U10392 ( .A1(n9227), .A2(n_T_702[27]), .Y(n9217) );
  NAND2X0_LVT U10393 ( .A1(n9222), .A2(n_T_642[7]), .Y(n9216) );
  NAND3X0_LVT U10394 ( .A1(n9217), .A2(n9224), .A3(n9216), .Y(alu_io_in2[27])
         );
  NAND2X0_LVT U10395 ( .A1(n9227), .A2(n_T_702[28]), .Y(n9219) );
  NAND2X0_LVT U10396 ( .A1(n9222), .A2(n_T_642[8]), .Y(n9218) );
  NAND3X0_LVT U10397 ( .A1(n9219), .A2(n9224), .A3(n9218), .Y(alu_io_in2[28])
         );
  NAND2X0_LVT U10398 ( .A1(n9227), .A2(n_T_702[29]), .Y(n9221) );
  NAND2X0_LVT U10399 ( .A1(n9222), .A2(n_T_642[9]), .Y(n9220) );
  NAND3X0_LVT U10400 ( .A1(n9221), .A2(n9224), .A3(n9220), .Y(alu_io_in2[29])
         );
  NAND2X0_LVT U10401 ( .A1(n9227), .A2(n_T_702[30]), .Y(n9225) );
  NAND2X0_LVT U10402 ( .A1(n9222), .A2(n_T_642[10]), .Y(n9223) );
  NAND3X0_LVT U10403 ( .A1(n9225), .A2(n9224), .A3(n9223), .Y(alu_io_in2[30])
         );
  AO21X1_LVT U10404 ( .A1(n9227), .A2(n_T_702[31]), .A3(n9226), .Y(
        alu_io_in2[31]) );
  AO21X1_LVT U10405 ( .A1(n9227), .A2(n_T_702[32]), .A3(n9226), .Y(
        alu_io_in2[32]) );
  AO21X1_LVT U10406 ( .A1(n9227), .A2(n_T_702[33]), .A3(n9226), .Y(
        alu_io_in2[33]) );
  AO21X1_LVT U10407 ( .A1(n9227), .A2(n_T_702[34]), .A3(n9226), .Y(
        alu_io_in2[34]) );
  AO21X1_LVT U10408 ( .A1(n9227), .A2(n_T_702[35]), .A3(n9226), .Y(
        alu_io_in2[35]) );
  AO21X1_LVT U10409 ( .A1(n9227), .A2(n_T_702[36]), .A3(n9226), .Y(
        alu_io_in2[36]) );
  AO21X1_LVT U10410 ( .A1(n9227), .A2(n_T_702[37]), .A3(n9226), .Y(
        alu_io_in2[37]) );
  AO21X1_LVT U10411 ( .A1(n9227), .A2(n_T_702[38]), .A3(n9226), .Y(
        alu_io_in2[38]) );
  AO21X1_LVT U10412 ( .A1(n9227), .A2(n_T_702[39]), .A3(n9226), .Y(
        alu_io_in2[39]) );
  AO21X1_LVT U10413 ( .A1(n9227), .A2(n_T_702[40]), .A3(n9226), .Y(
        alu_io_in2[40]) );
  AO21X1_LVT U10414 ( .A1(n9227), .A2(n_T_702[41]), .A3(n9226), .Y(
        alu_io_in2[41]) );
  AO21X1_LVT U10415 ( .A1(n9227), .A2(n_T_702[42]), .A3(n9226), .Y(
        alu_io_in2[42]) );
  AO21X1_LVT U10416 ( .A1(n9227), .A2(n_T_702[43]), .A3(n9226), .Y(
        alu_io_in2[43]) );
  AO21X1_LVT U10417 ( .A1(n9227), .A2(n_T_702[44]), .A3(n9226), .Y(
        alu_io_in2[44]) );
  AO21X1_LVT U10418 ( .A1(n9227), .A2(n_T_702[45]), .A3(n9226), .Y(
        alu_io_in2[45]) );
  AO21X1_LVT U10419 ( .A1(n9227), .A2(n_T_702[46]), .A3(n9226), .Y(
        alu_io_in2[46]) );
  AO21X1_LVT U10420 ( .A1(n9227), .A2(n_T_702[47]), .A3(n9226), .Y(
        alu_io_in2[47]) );
  AO21X1_LVT U10421 ( .A1(n9227), .A2(n_T_702[48]), .A3(n9226), .Y(
        alu_io_in2[48]) );
  AO21X1_LVT U10422 ( .A1(n9227), .A2(n_T_702[49]), .A3(n9226), .Y(
        alu_io_in2[49]) );
  AO21X1_LVT U10423 ( .A1(n9227), .A2(n_T_702[50]), .A3(n9226), .Y(
        alu_io_in2[50]) );
  AO21X1_LVT U10424 ( .A1(n9227), .A2(n_T_702[51]), .A3(n9226), .Y(
        alu_io_in2[51]) );
  AO21X1_LVT U10425 ( .A1(n9227), .A2(n_T_702[52]), .A3(n9226), .Y(
        alu_io_in2[52]) );
  AO21X1_LVT U10426 ( .A1(n9227), .A2(n_T_702[53]), .A3(n9226), .Y(
        alu_io_in2[53]) );
  AO21X1_LVT U10427 ( .A1(n9227), .A2(n_T_702[54]), .A3(n9226), .Y(
        alu_io_in2[54]) );
  AO21X1_LVT U10428 ( .A1(n9227), .A2(n_T_702[55]), .A3(n9226), .Y(
        alu_io_in2[55]) );
  AO21X1_LVT U10429 ( .A1(n9227), .A2(n_T_702[56]), .A3(n9226), .Y(
        alu_io_in2[56]) );
  AO21X1_LVT U10430 ( .A1(n9227), .A2(n_T_702[57]), .A3(n9226), .Y(
        alu_io_in2[57]) );
  AO21X1_LVT U10431 ( .A1(n9227), .A2(n_T_702[58]), .A3(n9226), .Y(
        alu_io_in2[58]) );
  AO21X1_LVT U10432 ( .A1(n9227), .A2(n_T_702[59]), .A3(n9226), .Y(
        alu_io_in2[59]) );
  AO21X1_LVT U10433 ( .A1(n9227), .A2(n_T_702[60]), .A3(n9226), .Y(
        alu_io_in2[60]) );
  AO21X1_LVT U10434 ( .A1(n9227), .A2(n_T_702[61]), .A3(n9226), .Y(
        alu_io_in2[61]) );
  AO21X1_LVT U10435 ( .A1(n9227), .A2(n_T_702[62]), .A3(n9226), .Y(
        alu_io_in2[62]) );
  AO21X1_LVT U10436 ( .A1(n9227), .A2(n_T_702[63]), .A3(n9226), .Y(
        alu_io_in2[63]) );
  OA21X1_LVT U10437 ( .A1(io_fpu_inst[14]), .A2(n9229), .A3(n9228), .Y(n9234)
         );
  NAND3X0_LVT U10438 ( .A1(n9234), .A2(n9233), .A3(n9232), .Y(N284) );
  INVX1_LVT U10439 ( .A(n9237), .Y(n9235) );
  AO22X1_LVT U10440 ( .A1(n9235), .A2(n9425), .A3(mem_reg_cause[0]), .A4(n1279), .Y(N533) );
  NAND2X0_LVT U10441 ( .A1(n3262), .A2(wb_reg_cause[0]), .Y(n9236) );
  NAND2X0_LVT U10442 ( .A1(n9240), .A2(n9236), .Y(wb_cause[0]) );
  AND2X1_LVT U10443 ( .A1(n9425), .A2(n9237), .Y(n9238) );
  AO21X1_LVT U10444 ( .A1(mem_reg_cause[2]), .A2(n1279), .A3(n9238), .Y(N535)
         );
  OR2X1_LVT U10445 ( .A1(wb_reg_cause[2]), .A2(n576), .Y(wb_cause[2]) );
  AO21X1_LVT U10446 ( .A1(mem_reg_cause[3]), .A2(n1279), .A3(n9238), .Y(N536)
         );
  NAND2X0_LVT U10447 ( .A1(n9249), .A2(n9239), .Y(n9241) );
  OAI22X1_LVT U10448 ( .A1(n576), .A2(n3565), .A3(n9241), .A4(n9240), .Y(
        wb_cause[3]) );
  MUX21X1_LVT U10449 ( .A1(csr_io_interrupt_cause[1]), .A2(n9245), .S0(n9448), 
        .Y(N304) );
  AND2X1_LVT U10450 ( .A1(io_dmem_s2_xcpt_ae_st), .A2(n9246), .Y(n9248) );
  OA21X1_LVT U10451 ( .A1(io_dmem_s2_xcpt_pf_st), .A2(n9248), .A3(n9247), .Y(
        n9250) );
  OA21X1_LVT U10452 ( .A1(io_dmem_s2_xcpt_ma_st), .A2(n9250), .A3(n9249), .Y(
        n9251) );
  INVX1_LVT U10453 ( .A(wb_cause[2]), .Y(n9252) );
  AND2X1_LVT U10454 ( .A1(n3262), .A2(wb_reg_cause[63]), .Y(wb_cause[63]) );
  AND2X1_LVT U10455 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[0]), .Y(
        csr_io_tval[0]) );
  AND2X1_LVT U10456 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[1]), .Y(
        csr_io_tval[1]) );
  AND2X1_LVT U10457 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[2]), .Y(
        csr_io_tval[2]) );
  AND2X1_LVT U10458 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[3]), .Y(
        csr_io_tval[3]) );
  AND2X1_LVT U10459 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[4]), .Y(
        csr_io_tval[4]) );
  AND2X1_LVT U10460 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[5]), .Y(
        csr_io_tval[5]) );
  AND2X1_LVT U10461 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[6]), .Y(
        csr_io_tval[6]) );
  AND2X1_LVT U10462 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[7]), .Y(
        csr_io_tval[7]) );
  AND2X1_LVT U10463 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[8]), .Y(
        csr_io_tval[8]) );
  AND2X1_LVT U10464 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[9]), .Y(
        csr_io_tval[9]) );
  AND2X1_LVT U10465 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[10]), .Y(
        csr_io_tval[10]) );
  AND2X1_LVT U10466 ( .A1(n4055), .A2(io_imem_sfence_bits_addr[11]), .Y(
        csr_io_tval[11]) );
  AND2X1_LVT U10467 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[12]), .Y(
        csr_io_tval[12]) );
  AND2X1_LVT U10468 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[13]), .Y(
        csr_io_tval[13]) );
  AND2X1_LVT U10469 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[14]), .Y(
        csr_io_tval[14]) );
  AND2X1_LVT U10470 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[15]), .Y(
        csr_io_tval[15]) );
  AND2X1_LVT U10471 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[16]), .Y(
        csr_io_tval[16]) );
  AND2X1_LVT U10472 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[17]), .Y(
        csr_io_tval[17]) );
  AND2X1_LVT U10473 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[18]), .Y(
        csr_io_tval[18]) );
  AND2X1_LVT U10474 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[19]), .Y(
        csr_io_tval[19]) );
  AND2X1_LVT U10475 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[20]), .Y(
        csr_io_tval[20]) );
  AND2X1_LVT U10476 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[21]), .Y(
        csr_io_tval[21]) );
  AND2X1_LVT U10477 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[22]), .Y(
        csr_io_tval[22]) );
  AND2X1_LVT U10478 ( .A1(n4056), .A2(io_imem_sfence_bits_addr[23]), .Y(
        csr_io_tval[23]) );
  AND2X1_LVT U10479 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[24]), .Y(
        csr_io_tval[24]) );
  AND2X1_LVT U10480 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[25]), .Y(
        csr_io_tval[25]) );
  AND2X1_LVT U10481 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[26]), .Y(
        csr_io_tval[26]) );
  AND2X1_LVT U10482 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[27]), .Y(
        csr_io_tval[27]) );
  AND2X1_LVT U10483 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[28]), .Y(
        csr_io_tval[28]) );
  AND2X1_LVT U10484 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[29]), .Y(
        csr_io_tval[29]) );
  AND2X1_LVT U10485 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[30]), .Y(
        csr_io_tval[30]) );
  AND2X1_LVT U10486 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[31]), .Y(
        csr_io_tval[31]) );
  AND2X1_LVT U10487 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[32]), .Y(
        csr_io_tval[32]) );
  AND2X1_LVT U10488 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[33]), .Y(
        csr_io_tval[33]) );
  AND2X1_LVT U10489 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[34]), .Y(
        csr_io_tval[34]) );
  AND2X1_LVT U10490 ( .A1(n4057), .A2(io_imem_sfence_bits_addr[35]), .Y(
        csr_io_tval[35]) );
  AND2X1_LVT U10491 ( .A1(n9276), .A2(io_imem_sfence_bits_addr[36]), .Y(
        csr_io_tval[36]) );
  AND2X1_LVT U10492 ( .A1(n9276), .A2(io_imem_sfence_bits_addr[37]), .Y(
        csr_io_tval[37]) );
  AND2X1_LVT U10493 ( .A1(n9276), .A2(io_imem_sfence_bits_addr[38]), .Y(
        csr_io_tval[38]) );
  NOR4X1_LVT U10494 ( .A1(n_T_1165[45]), .A2(n_T_1165[44]), .A3(n_T_1165[46]), 
        .A4(n_T_1165[47]), .Y(n9258) );
  NOR4X1_LVT U10495 ( .A1(n_T_1165[40]), .A2(n_T_1165[42]), .A3(n_T_1165[41]), 
        .A4(n_T_1165[43]), .Y(n9257) );
  NAND2X0_LVT U10496 ( .A1(n9258), .A2(n9257), .Y(n9264) );
  NOR4X1_LVT U10497 ( .A1(n_T_1165[57]), .A2(n_T_1165[56]), .A3(n_T_1165[58]), 
        .A4(n_T_1165[60]), .Y(n9262) );
  NOR4X1_LVT U10498 ( .A1(n_T_1165[52]), .A2(n_T_1165[54]), .A3(n_T_1165[53]), 
        .A4(n_T_1165[55]), .Y(n9261) );
  NOR4X1_LVT U10499 ( .A1(n_T_1165[48]), .A2(n_T_1165[49]), .A3(n_T_1165[51]), 
        .A4(n_T_1165[50]), .Y(n9260) );
  NOR4X1_LVT U10500 ( .A1(n_T_1165[59]), .A2(n_T_1165[61]), .A3(n_T_1165[63]), 
        .A4(n_T_1165[62]), .Y(n9259) );
  NAND4X0_LVT U10501 ( .A1(n9262), .A2(n9261), .A3(n9260), .A4(n9259), .Y(
        n9263) );
  OR2X1_LVT U10502 ( .A1(n9264), .A2(n9263), .Y(n9273) );
  NAND4X0_LVT U10503 ( .A1(n_T_1165[61]), .A2(n_T_1165[63]), .A3(n_T_1165[62]), 
        .A4(n_T_1165[59]), .Y(n9268) );
  NAND4X0_LVT U10504 ( .A1(n_T_1165[57]), .A2(n_T_1165[56]), .A3(n_T_1165[58]), 
        .A4(n_T_1165[60]), .Y(n9267) );
  NAND4X0_LVT U10505 ( .A1(n_T_1165[52]), .A2(n_T_1165[54]), .A3(n_T_1165[53]), 
        .A4(n_T_1165[55]), .Y(n9266) );
  NAND4X0_LVT U10506 ( .A1(n_T_1165[48]), .A2(n_T_1165[49]), .A3(n_T_1165[51]), 
        .A4(n_T_1165[50]), .Y(n9265) );
  NOR4X1_LVT U10507 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .Y(n9271) );
  AND4X1_LVT U10508 ( .A1(n_T_1165[45]), .A2(n_T_1165[44]), .A3(n_T_1165[46]), 
        .A4(n_T_1165[47]), .Y(n9270) );
  AND4X1_LVT U10509 ( .A1(n_T_1165[40]), .A2(n_T_1165[42]), .A3(n_T_1165[41]), 
        .A4(n_T_1165[43]), .Y(n9269) );
  NAND3X0_LVT U10510 ( .A1(n9271), .A2(n9270), .A3(n9269), .Y(n9272) );
  MUX21X1_LVT U10511 ( .A1(n9273), .A2(n9272), .S0(n_T_1165[39]), .Y(n9274) );
  MUX21X1_LVT U10512 ( .A1(n_T_1165[39]), .A2(n3228), .S0(n9274), .Y(n9275) );
  AND2X1_LVT U10513 ( .A1(n9276), .A2(n9275), .Y(csr_io_tval[39]) );
  AND2X1_LVT U10514 ( .A1(wb_reg_valid), .A2(wb_ctrl_csr[2]), .Y(
        csr_io_rw_cmd_2_) );
  NAND3X0_LVT U10515 ( .A1(n9279), .A2(n9278), .A3(n9277), .Y(n9284) );
  NOR3X0_LVT U10516 ( .A1(mem_reg_valid), .A2(mem_reg_xcpt_interrupt), .A3(
        mem_reg_replay), .Y(n9449) );
  INVX1_LVT U10517 ( .A(n9449), .Y(mem_pc_valid) );
  AND2X1_LVT U10518 ( .A1(wb_reg_valid), .A2(wb_reg_sfence), .Y(
        io_imem_sfence_valid) );
  MUX21X1_LVT U10519 ( .A1(mem_reg_rs2[0]), .A2(io_fpu_store_data[0]), .S0(
        n2498), .Y(io_dmem_s1_data_data[0]) );
  MUX21X1_LVT U10520 ( .A1(mem_reg_rs2[1]), .A2(io_fpu_store_data[1]), .S0(
        n2498), .Y(io_dmem_s1_data_data[1]) );
  MUX21X1_LVT U10521 ( .A1(mem_reg_rs2[2]), .A2(io_fpu_store_data[2]), .S0(
        n2498), .Y(io_dmem_s1_data_data[2]) );
  MUX21X1_LVT U10522 ( .A1(mem_reg_rs2[3]), .A2(io_fpu_store_data[3]), .S0(
        n2498), .Y(io_dmem_s1_data_data[3]) );
  MUX21X1_LVT U10523 ( .A1(mem_reg_rs2[4]), .A2(io_fpu_store_data[4]), .S0(
        n2492), .Y(io_dmem_s1_data_data[4]) );
  MUX21X1_LVT U10524 ( .A1(mem_reg_rs2[5]), .A2(io_fpu_store_data[5]), .S0(
        n2498), .Y(io_dmem_s1_data_data[5]) );
  MUX21X1_LVT U10525 ( .A1(mem_reg_rs2[6]), .A2(io_fpu_store_data[6]), .S0(
        n2498), .Y(io_dmem_s1_data_data[6]) );
  MUX21X1_LVT U10526 ( .A1(mem_reg_rs2[7]), .A2(io_fpu_store_data[7]), .S0(
        n2498), .Y(io_dmem_s1_data_data[7]) );
  NAND2X0_LVT U10527 ( .A1(n313), .A2(io_dmem_req_bits_size[1]), .Y(n9292) );
  NAND2X0_LVT U10528 ( .A1(n586), .A2(io_dmem_req_bits_size[0]), .Y(n9289) );
  NAND2X0_LVT U10529 ( .A1(n9292), .A2(n9289), .Y(n9290) );
  AO22X1_LVT U10530 ( .A1(n_T_702[8]), .A2(n9290), .A3(n9291), .A4(n_T_702[0]), 
        .Y(n9293) );
  AO21X1_LVT U10531 ( .A1(n4058), .A2(n_T_702[8]), .A3(n9293), .Y(N469) );
  MUX21X1_LVT U10532 ( .A1(mem_reg_rs2[8]), .A2(io_fpu_store_data[8]), .S0(
        n2492), .Y(io_dmem_s1_data_data[8]) );
  AO22X1_LVT U10533 ( .A1(n_T_702[9]), .A2(n9290), .A3(n9291), .A4(n_T_702[1]), 
        .Y(n9295) );
  AO21X1_LVT U10534 ( .A1(n4058), .A2(n_T_702[9]), .A3(n9295), .Y(N470) );
  MUX21X1_LVT U10535 ( .A1(mem_reg_rs2[9]), .A2(io_fpu_store_data[9]), .S0(
        n2498), .Y(io_dmem_s1_data_data[9]) );
  AO22X1_LVT U10536 ( .A1(n_T_702[10]), .A2(n9290), .A3(n9291), .A4(n_T_702[2]), .Y(n9296) );
  AO21X1_LVT U10537 ( .A1(n4058), .A2(n_T_702[10]), .A3(n9296), .Y(N471) );
  MUX21X1_LVT U10538 ( .A1(mem_reg_rs2[10]), .A2(io_fpu_store_data[10]), .S0(
        n2498), .Y(io_dmem_s1_data_data[10]) );
  AO22X1_LVT U10539 ( .A1(n_T_702[11]), .A2(n9290), .A3(n9291), .A4(n_T_702[3]), .Y(n9297) );
  AO21X1_LVT U10540 ( .A1(n4058), .A2(n_T_702[11]), .A3(n9297), .Y(N472) );
  MUX21X1_LVT U10541 ( .A1(mem_reg_rs2[11]), .A2(io_fpu_store_data[11]), .S0(
        n2498), .Y(io_dmem_s1_data_data[11]) );
  AO22X1_LVT U10542 ( .A1(n_T_702[12]), .A2(n9290), .A3(n9291), .A4(n_T_702[4]), .Y(n9298) );
  AO21X1_LVT U10543 ( .A1(n4058), .A2(n_T_702[12]), .A3(n9298), .Y(N473) );
  MUX21X1_LVT U10544 ( .A1(mem_reg_rs2[12]), .A2(io_fpu_store_data[12]), .S0(
        n2498), .Y(io_dmem_s1_data_data[12]) );
  AO22X1_LVT U10545 ( .A1(n_T_702[5]), .A2(n9291), .A3(n9290), .A4(n_T_702[13]), .Y(n9299) );
  AO21X1_LVT U10546 ( .A1(n4058), .A2(n_T_702[13]), .A3(n9299), .Y(N474) );
  MUX21X1_LVT U10547 ( .A1(mem_reg_rs2[13]), .A2(io_fpu_store_data[13]), .S0(
        n2498), .Y(io_dmem_s1_data_data[13]) );
  AO22X1_LVT U10548 ( .A1(n_T_702[6]), .A2(n9291), .A3(n9290), .A4(n_T_702[14]), .Y(n9300) );
  AO21X1_LVT U10549 ( .A1(n4058), .A2(n_T_702[14]), .A3(n9300), .Y(N475) );
  MUX21X1_LVT U10550 ( .A1(mem_reg_rs2[14]), .A2(io_fpu_store_data[14]), .S0(
        n2498), .Y(io_dmem_s1_data_data[14]) );
  AO22X1_LVT U10551 ( .A1(n_T_702[7]), .A2(n9291), .A3(n9290), .A4(n_T_702[15]), .Y(n9302) );
  AO21X1_LVT U10552 ( .A1(n4058), .A2(n_T_702[15]), .A3(n9302), .Y(N476) );
  MUX21X1_LVT U10553 ( .A1(mem_reg_rs2[15]), .A2(io_fpu_store_data[15]), .S0(
        n2498), .Y(io_dmem_s1_data_data[15]) );
  MUX21X1_LVT U10554 ( .A1(n_T_702[16]), .A2(n_T_702[0]), .S0(n586), .Y(N477)
         );
  MUX21X1_LVT U10555 ( .A1(mem_reg_rs2[16]), .A2(io_fpu_store_data[16]), .S0(
        n2492), .Y(io_dmem_s1_data_data[16]) );
  MUX21X1_LVT U10556 ( .A1(n_T_702[17]), .A2(n_T_702[1]), .S0(n2515), .Y(N478)
         );
  MUX21X1_LVT U10557 ( .A1(mem_reg_rs2[17]), .A2(io_fpu_store_data[17]), .S0(
        n2498), .Y(io_dmem_s1_data_data[17]) );
  MUX21X1_LVT U10558 ( .A1(n_T_702[18]), .A2(n_T_702[2]), .S0(n586), .Y(N479)
         );
  MUX21X1_LVT U10559 ( .A1(mem_reg_rs2[18]), .A2(io_fpu_store_data[18]), .S0(
        n2498), .Y(io_dmem_s1_data_data[18]) );
  MUX21X1_LVT U10560 ( .A1(n_T_702[19]), .A2(n_T_702[3]), .S0(n2515), .Y(N480)
         );
  MUX21X1_LVT U10561 ( .A1(mem_reg_rs2[19]), .A2(io_fpu_store_data[19]), .S0(
        n2498), .Y(io_dmem_s1_data_data[19]) );
  MUX21X1_LVT U10562 ( .A1(n_T_702[20]), .A2(n_T_702[4]), .S0(n586), .Y(N481)
         );
  MUX21X1_LVT U10563 ( .A1(mem_reg_rs2[20]), .A2(io_fpu_store_data[20]), .S0(
        n2498), .Y(io_dmem_s1_data_data[20]) );
  MUX21X1_LVT U10564 ( .A1(n_T_702[5]), .A2(n_T_702[21]), .S0(
        io_dmem_req_bits_size[1]), .Y(N482) );
  MUX21X1_LVT U10565 ( .A1(mem_reg_rs2[21]), .A2(io_fpu_store_data[21]), .S0(
        n2498), .Y(io_dmem_s1_data_data[21]) );
  MUX21X1_LVT U10566 ( .A1(n_T_702[6]), .A2(n_T_702[22]), .S0(
        io_dmem_req_bits_size[1]), .Y(N483) );
  MUX21X1_LVT U10567 ( .A1(mem_reg_rs2[22]), .A2(io_fpu_store_data[22]), .S0(
        n2498), .Y(io_dmem_s1_data_data[22]) );
  MUX21X1_LVT U10568 ( .A1(n_T_702[7]), .A2(n_T_702[23]), .S0(
        io_dmem_req_bits_size[1]), .Y(N484) );
  MUX21X1_LVT U10569 ( .A1(mem_reg_rs2[23]), .A2(io_fpu_store_data[23]), .S0(
        n2498), .Y(io_dmem_s1_data_data[23]) );
  MUX21X1_LVT U10570 ( .A1(n_T_702[24]), .A2(n9293), .S0(n586), .Y(N485) );
  MUX21X1_LVT U10571 ( .A1(mem_reg_rs2[24]), .A2(io_fpu_store_data[24]), .S0(
        n2498), .Y(io_dmem_s1_data_data[24]) );
  MUX21X1_LVT U10572 ( .A1(n_T_702[25]), .A2(n9295), .S0(n586), .Y(N486) );
  MUX21X1_LVT U10573 ( .A1(mem_reg_rs2[25]), .A2(io_fpu_store_data[25]), .S0(
        n2498), .Y(io_dmem_s1_data_data[25]) );
  MUX21X1_LVT U10574 ( .A1(n_T_702[26]), .A2(n9296), .S0(n586), .Y(N487) );
  MUX21X1_LVT U10575 ( .A1(mem_reg_rs2[26]), .A2(io_fpu_store_data[26]), .S0(
        n2498), .Y(io_dmem_s1_data_data[26]) );
  MUX21X1_LVT U10576 ( .A1(n_T_702[27]), .A2(n9297), .S0(n586), .Y(N488) );
  MUX21X1_LVT U10577 ( .A1(mem_reg_rs2[27]), .A2(io_fpu_store_data[27]), .S0(
        n2498), .Y(io_dmem_s1_data_data[27]) );
  MUX21X1_LVT U10578 ( .A1(n_T_702[28]), .A2(n9298), .S0(n586), .Y(N489) );
  MUX21X1_LVT U10579 ( .A1(mem_reg_rs2[28]), .A2(io_fpu_store_data[28]), .S0(
        n2498), .Y(io_dmem_s1_data_data[28]) );
  MUX21X1_LVT U10580 ( .A1(n_T_702[29]), .A2(n9299), .S0(n586), .Y(N490) );
  MUX21X1_LVT U10581 ( .A1(mem_reg_rs2[29]), .A2(io_fpu_store_data[29]), .S0(
        n2498), .Y(io_dmem_s1_data_data[29]) );
  MUX21X1_LVT U10582 ( .A1(n_T_702[30]), .A2(n9300), .S0(n586), .Y(N491) );
  MUX21X1_LVT U10583 ( .A1(mem_reg_rs2[30]), .A2(io_fpu_store_data[30]), .S0(
        n2498), .Y(io_dmem_s1_data_data[30]) );
  MUX21X1_LVT U10584 ( .A1(n_T_702[31]), .A2(n9302), .S0(n2515), .Y(N492) );
  MUX21X1_LVT U10585 ( .A1(mem_reg_rs2[31]), .A2(io_fpu_store_data[31]), .S0(
        n2492), .Y(io_dmem_s1_data_data[31]) );
  MUX21X1_LVT U10586 ( .A1(n_T_702[32]), .A2(n_T_702[0]), .S0(n3234), .Y(N493)
         );
  MUX21X1_LVT U10587 ( .A1(mem_reg_rs2[32]), .A2(io_fpu_store_data[32]), .S0(
        n2498), .Y(io_dmem_s1_data_data[32]) );
  MUX21X1_LVT U10588 ( .A1(n_T_702[33]), .A2(n_T_702[1]), .S0(n3234), .Y(N494)
         );
  MUX21X1_LVT U10589 ( .A1(mem_reg_rs2[33]), .A2(io_fpu_store_data[33]), .S0(
        n2498), .Y(io_dmem_s1_data_data[33]) );
  MUX21X1_LVT U10590 ( .A1(n_T_702[34]), .A2(n_T_702[2]), .S0(n3234), .Y(N495)
         );
  MUX21X1_LVT U10591 ( .A1(mem_reg_rs2[34]), .A2(io_fpu_store_data[34]), .S0(
        n2498), .Y(io_dmem_s1_data_data[34]) );
  MUX21X1_LVT U10592 ( .A1(n_T_702[35]), .A2(n_T_702[3]), .S0(n3234), .Y(N496)
         );
  MUX21X1_LVT U10593 ( .A1(mem_reg_rs2[35]), .A2(io_fpu_store_data[35]), .S0(
        n2492), .Y(io_dmem_s1_data_data[35]) );
  MUX21X1_LVT U10594 ( .A1(n_T_702[36]), .A2(n_T_702[4]), .S0(n3234), .Y(N497)
         );
  MUX21X1_LVT U10595 ( .A1(mem_reg_rs2[36]), .A2(io_fpu_store_data[36]), .S0(
        n2498), .Y(io_dmem_s1_data_data[36]) );
  MUX21X1_LVT U10596 ( .A1(n_T_702[37]), .A2(n_T_702[5]), .S0(n3234), .Y(N498)
         );
  MUX21X1_LVT U10597 ( .A1(mem_reg_rs2[37]), .A2(io_fpu_store_data[37]), .S0(
        n2498), .Y(io_dmem_s1_data_data[37]) );
  MUX21X1_LVT U10598 ( .A1(n_T_702[38]), .A2(n_T_702[6]), .S0(n3234), .Y(N499)
         );
  MUX21X1_LVT U10599 ( .A1(mem_reg_rs2[38]), .A2(io_fpu_store_data[38]), .S0(
        n2498), .Y(io_dmem_s1_data_data[38]) );
  MUX21X1_LVT U10600 ( .A1(n_T_702[39]), .A2(n_T_702[7]), .S0(n3234), .Y(N500)
         );
  MUX21X1_LVT U10601 ( .A1(mem_reg_rs2[39]), .A2(io_fpu_store_data[39]), .S0(
        n2492), .Y(io_dmem_s1_data_data[39]) );
  AO21X1_LVT U10602 ( .A1(n4058), .A2(n_T_702[40]), .A3(n9293), .Y(N501) );
  MUX21X1_LVT U10603 ( .A1(mem_reg_rs2[40]), .A2(io_fpu_store_data[40]), .S0(
        n2498), .Y(io_dmem_s1_data_data[40]) );
  AO21X1_LVT U10604 ( .A1(n4058), .A2(n_T_702[41]), .A3(n9295), .Y(N502) );
  MUX21X1_LVT U10605 ( .A1(mem_reg_rs2[41]), .A2(io_fpu_store_data[41]), .S0(
        n2498), .Y(io_dmem_s1_data_data[41]) );
  AO21X1_LVT U10606 ( .A1(n4058), .A2(n_T_702[42]), .A3(n9296), .Y(N503) );
  MUX21X1_LVT U10607 ( .A1(mem_reg_rs2[42]), .A2(io_fpu_store_data[42]), .S0(
        n2498), .Y(io_dmem_s1_data_data[42]) );
  AO21X1_LVT U10608 ( .A1(n4058), .A2(n_T_702[43]), .A3(n9297), .Y(N504) );
  MUX21X1_LVT U10609 ( .A1(mem_reg_rs2[43]), .A2(io_fpu_store_data[43]), .S0(
        n2492), .Y(io_dmem_s1_data_data[43]) );
  AO21X1_LVT U10610 ( .A1(n4058), .A2(n_T_702[44]), .A3(n9298), .Y(N505) );
  MUX21X1_LVT U10611 ( .A1(mem_reg_rs2[44]), .A2(io_fpu_store_data[44]), .S0(
        n2498), .Y(io_dmem_s1_data_data[44]) );
  AO21X1_LVT U10612 ( .A1(n4058), .A2(n_T_702[45]), .A3(n9299), .Y(N506) );
  MUX21X1_LVT U10613 ( .A1(mem_reg_rs2[45]), .A2(io_fpu_store_data[45]), .S0(
        n2498), .Y(io_dmem_s1_data_data[45]) );
  AO21X1_LVT U10614 ( .A1(n4058), .A2(n_T_702[46]), .A3(n9300), .Y(N507) );
  MUX21X1_LVT U10615 ( .A1(mem_reg_rs2[46]), .A2(io_fpu_store_data[46]), .S0(
        n2498), .Y(io_dmem_s1_data_data[46]) );
  AO21X1_LVT U10616 ( .A1(n4058), .A2(n_T_702[47]), .A3(n9302), .Y(N508) );
  MUX21X1_LVT U10617 ( .A1(mem_reg_rs2[47]), .A2(io_fpu_store_data[47]), .S0(
        n2492), .Y(io_dmem_s1_data_data[47]) );
  MUX21X1_LVT U10618 ( .A1(mem_reg_rs2[48]), .A2(io_fpu_store_data[48]), .S0(
        n2498), .Y(io_dmem_s1_data_data[48]) );
  MUX21X1_LVT U10619 ( .A1(mem_reg_rs2[49]), .A2(io_fpu_store_data[49]), .S0(
        n2498), .Y(io_dmem_s1_data_data[49]) );
  MUX21X1_LVT U10620 ( .A1(mem_reg_rs2[50]), .A2(io_fpu_store_data[50]), .S0(
        n2498), .Y(io_dmem_s1_data_data[50]) );
  MUX21X1_LVT U10621 ( .A1(mem_reg_rs2[51]), .A2(io_fpu_store_data[51]), .S0(
        n2492), .Y(io_dmem_s1_data_data[51]) );
  MUX21X1_LVT U10622 ( .A1(mem_reg_rs2[52]), .A2(io_fpu_store_data[52]), .S0(
        n2492), .Y(io_dmem_s1_data_data[52]) );
  MUX21X1_LVT U10623 ( .A1(mem_reg_rs2[53]), .A2(io_fpu_store_data[53]), .S0(
        n2498), .Y(io_dmem_s1_data_data[53]) );
  MUX21X1_LVT U10624 ( .A1(mem_reg_rs2[54]), .A2(io_fpu_store_data[54]), .S0(
        n2498), .Y(io_dmem_s1_data_data[54]) );
  MUX21X1_LVT U10625 ( .A1(mem_reg_rs2[55]), .A2(io_fpu_store_data[55]), .S0(
        n2498), .Y(io_dmem_s1_data_data[55]) );
  MUX21X1_LVT U10626 ( .A1(mem_reg_rs2[56]), .A2(io_fpu_store_data[56]), .S0(
        n2492), .Y(io_dmem_s1_data_data[56]) );
  AO22X1_LVT U10627 ( .A1(n_T_702[57]), .A2(n4058), .A3(n9301), .A4(
        n_T_702[25]), .Y(n9294) );
  AO21X1_LVT U10628 ( .A1(n2515), .A2(n9295), .A3(n9294), .Y(N518) );
  MUX21X1_LVT U10629 ( .A1(mem_reg_rs2[57]), .A2(io_fpu_store_data[57]), .S0(
        n2498), .Y(io_dmem_s1_data_data[57]) );
  MUX21X1_LVT U10630 ( .A1(mem_reg_rs2[58]), .A2(io_fpu_store_data[58]), .S0(
        n2498), .Y(io_dmem_s1_data_data[58]) );
  MUX21X1_LVT U10631 ( .A1(mem_reg_rs2[59]), .A2(io_fpu_store_data[59]), .S0(
        n2498), .Y(io_dmem_s1_data_data[59]) );
  MUX21X1_LVT U10632 ( .A1(mem_reg_rs2[60]), .A2(io_fpu_store_data[60]), .S0(
        n2492), .Y(io_dmem_s1_data_data[60]) );
  MUX21X1_LVT U10633 ( .A1(mem_reg_rs2[61]), .A2(io_fpu_store_data[61]), .S0(
        n2498), .Y(io_dmem_s1_data_data[61]) );
  MUX21X1_LVT U10634 ( .A1(mem_reg_rs2[62]), .A2(io_fpu_store_data[62]), .S0(
        n2498), .Y(io_dmem_s1_data_data[62]) );
  MUX21X1_LVT U10635 ( .A1(mem_reg_rs2[63]), .A2(io_fpu_store_data[63]), .S0(
        n2498), .Y(io_dmem_s1_data_data[63]) );
  NAND4X0_LVT U10636 ( .A1(n9306), .A2(n9305), .A3(n9304), .A4(n9303), .Y(
        n9317) );
  NAND4X0_LVT U10637 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .Y(
        n9316) );
  NOR4X1_LVT U10638 ( .A1(io_fpu_fromint_data[40]), .A2(
        io_fpu_fromint_data[42]), .A3(io_fpu_fromint_data[41]), .A4(
        io_fpu_fromint_data[43]), .Y(n9314) );
  NOR4X1_LVT U10639 ( .A1(io_fpu_fromint_data[45]), .A2(
        io_fpu_fromint_data[44]), .A3(io_fpu_fromint_data[46]), .A4(
        io_fpu_fromint_data[48]), .Y(n9313) );
  NOR4X1_LVT U10640 ( .A1(io_fpu_fromint_data[47]), .A2(
        io_fpu_fromint_data[49]), .A3(io_fpu_fromint_data[51]), .A4(
        io_fpu_fromint_data[50]), .Y(n9312) );
  NOR4X1_LVT U10641 ( .A1(io_fpu_fromint_data[52]), .A2(
        io_fpu_fromint_data[54]), .A3(io_fpu_fromint_data[53]), .A4(
        io_fpu_fromint_data[55]), .Y(n9311) );
  NAND4X0_LVT U10642 ( .A1(n9314), .A2(n9313), .A3(n9312), .A4(n9311), .Y(
        n9315) );
  OR3X1_LVT U10643 ( .A1(n9317), .A2(n9316), .A3(n9315), .Y(n9326) );
  NAND4X0_LVT U10644 ( .A1(io_fpu_fromint_data[57]), .A2(
        io_fpu_fromint_data[56]), .A3(io_fpu_fromint_data[58]), .A4(
        io_fpu_fromint_data[60]), .Y(n9324) );
  NAND4X0_LVT U10645 ( .A1(io_fpu_fromint_data[59]), .A2(
        io_fpu_fromint_data[61]), .A3(io_fpu_fromint_data[63]), .A4(
        io_fpu_fromint_data[62]), .Y(n9323) );
  AND4X1_LVT U10646 ( .A1(io_fpu_fromint_data[40]), .A2(
        io_fpu_fromint_data[42]), .A3(io_fpu_fromint_data[41]), .A4(
        io_fpu_fromint_data[43]), .Y(n9321) );
  AND4X1_LVT U10647 ( .A1(io_fpu_fromint_data[45]), .A2(
        io_fpu_fromint_data[44]), .A3(io_fpu_fromint_data[46]), .A4(
        io_fpu_fromint_data[48]), .Y(n9320) );
  AND4X1_LVT U10648 ( .A1(io_fpu_fromint_data[47]), .A2(
        io_fpu_fromint_data[49]), .A3(io_fpu_fromint_data[51]), .A4(
        io_fpu_fromint_data[50]), .Y(n9319) );
  AND4X1_LVT U10649 ( .A1(io_fpu_fromint_data[52]), .A2(
        io_fpu_fromint_data[54]), .A3(io_fpu_fromint_data[53]), .A4(
        io_fpu_fromint_data[55]), .Y(n9318) );
  NAND4X0_LVT U10650 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .Y(
        n9322) );
  OR3X1_LVT U10651 ( .A1(n9324), .A2(n9323), .A3(n9322), .Y(n9325) );
  MUX21X1_LVT U10652 ( .A1(n9326), .A2(n9325), .S0(io_fpu_fromint_data[39]), 
        .Y(n9327) );
  MUX21X1_LVT U10653 ( .A1(alu_io_adder_out_39_), .A2(n9328), .S0(n9327), .Y(
        io_dmem_req_bits_addr[39]) );
  NAND4X0_LVT U10654 ( .A1(n3310), .A2(n3104), .A3(
        io_imem_bht_update_bits_branch), .A4(n555), .Y(n9329) );
  INVX1_LVT U10655 ( .A(n9512), .Y(n9333) );
  AO222X1_LVT U10656 ( .A1(n4065), .A2(csr_io_evec[1]), .A3(n4062), .A4(
        csr_io_pc[1]), .A5(n9333), .A6(n4060), .Y(io_imem_req_bits_pc[1]) );
  AO22X1_LVT U10657 ( .A1(n4063), .A2(csr_io_pc[2]), .A3(n9334), .A4(n4060), 
        .Y(n9335) );
  AO21X1_LVT U10658 ( .A1(n4067), .A2(csr_io_evec[2]), .A3(n9335), .Y(
        io_imem_req_bits_pc[2]) );
  AO22X1_LVT U10659 ( .A1(n4064), .A2(csr_io_pc[3]), .A3(n9336), .A4(n4061), 
        .Y(n9337) );
  AO21X1_LVT U10660 ( .A1(n4067), .A2(csr_io_evec[3]), .A3(n9337), .Y(
        io_imem_req_bits_pc[3]) );
  AO22X1_LVT U10661 ( .A1(n4064), .A2(csr_io_pc[4]), .A3(n9338), .A4(n4061), 
        .Y(n9339) );
  AO21X1_LVT U10662 ( .A1(n4067), .A2(csr_io_evec[4]), .A3(n9339), .Y(
        io_imem_req_bits_pc[4]) );
  AO22X1_LVT U10663 ( .A1(n4064), .A2(csr_io_pc[5]), .A3(n9340), .A4(n4061), 
        .Y(n9341) );
  AO21X1_LVT U10664 ( .A1(n4067), .A2(csr_io_evec[5]), .A3(n9341), .Y(
        io_imem_req_bits_pc[5]) );
  AO22X1_LVT U10665 ( .A1(n4064), .A2(csr_io_pc[6]), .A3(n9342), .A4(n4061), 
        .Y(n9343) );
  AO21X1_LVT U10666 ( .A1(n4067), .A2(csr_io_evec[6]), .A3(n9343), .Y(
        io_imem_req_bits_pc[6]) );
  AO22X1_LVT U10667 ( .A1(n4064), .A2(csr_io_pc[7]), .A3(n9344), .A4(n4061), 
        .Y(n9345) );
  AO21X1_LVT U10668 ( .A1(n4067), .A2(csr_io_evec[7]), .A3(n9345), .Y(
        io_imem_req_bits_pc[7]) );
  AO22X1_LVT U10669 ( .A1(n4064), .A2(csr_io_pc[8]), .A3(n9346), .A4(n4061), 
        .Y(n9347) );
  AO21X1_LVT U10670 ( .A1(n4067), .A2(csr_io_evec[8]), .A3(n9347), .Y(
        io_imem_req_bits_pc[8]) );
  AO22X1_LVT U10671 ( .A1(n4064), .A2(csr_io_pc[9]), .A3(n9348), .A4(n4061), 
        .Y(n9349) );
  AO21X1_LVT U10672 ( .A1(n4067), .A2(csr_io_evec[9]), .A3(n9349), .Y(
        io_imem_req_bits_pc[9]) );
  INVX1_LVT U10673 ( .A(n9509), .Y(n9350) );
  AO222X1_LVT U10674 ( .A1(n4065), .A2(csr_io_evec[10]), .A3(n4064), .A4(
        csr_io_pc[10]), .A5(n9350), .A6(n4059), .Y(io_imem_req_bits_pc[10]) );
  INVX1_LVT U10675 ( .A(n9490), .Y(n9351) );
  AO222X1_LVT U10676 ( .A1(n4065), .A2(csr_io_evec[11]), .A3(n4064), .A4(
        csr_io_pc[11]), .A5(n9351), .A6(n4059), .Y(io_imem_req_bits_pc[11]) );
  INVX1_LVT U10677 ( .A(n9491), .Y(n9352) );
  AO222X1_LVT U10678 ( .A1(n4065), .A2(csr_io_evec[12]), .A3(n4064), .A4(
        csr_io_pc[12]), .A5(n9352), .A6(n4059), .Y(io_imem_req_bits_pc[12]) );
  INVX1_LVT U10679 ( .A(n9500), .Y(n9353) );
  AO222X1_LVT U10680 ( .A1(n4065), .A2(csr_io_evec[13]), .A3(n4064), .A4(
        csr_io_pc[13]), .A5(n9353), .A6(n4059), .Y(io_imem_req_bits_pc[13]) );
  INVX1_LVT U10681 ( .A(n9506), .Y(n9354) );
  AO222X1_LVT U10682 ( .A1(n4065), .A2(csr_io_evec[14]), .A3(n4064), .A4(
        csr_io_pc[14]), .A5(n9354), .A6(n4059), .Y(io_imem_req_bits_pc[14]) );
  AO222X1_LVT U10683 ( .A1(n4065), .A2(csr_io_evec[15]), .A3(n4064), .A4(
        csr_io_pc[15]), .A5(n9355), .A6(n4059), .Y(io_imem_req_bits_pc[15]) );
  AO222X1_LVT U10684 ( .A1(n4065), .A2(csr_io_evec[16]), .A3(n4063), .A4(
        csr_io_pc[16]), .A5(n9356), .A6(n4059), .Y(io_imem_req_bits_pc[16]) );
  INVX1_LVT U10685 ( .A(n9487), .Y(n9357) );
  AO222X1_LVT U10686 ( .A1(n4065), .A2(csr_io_evec[17]), .A3(n4063), .A4(
        csr_io_pc[17]), .A5(n9357), .A6(n4059), .Y(io_imem_req_bits_pc[17]) );
  INVX1_LVT U10687 ( .A(n9496), .Y(n9358) );
  AO222X1_LVT U10688 ( .A1(n4065), .A2(csr_io_evec[18]), .A3(n4063), .A4(
        csr_io_pc[18]), .A5(n9358), .A6(n4059), .Y(io_imem_req_bits_pc[18]) );
  INVX1_LVT U10689 ( .A(n9510), .Y(n9359) );
  AO222X1_LVT U10690 ( .A1(n4065), .A2(csr_io_evec[19]), .A3(n4063), .A4(
        csr_io_pc[19]), .A5(n9359), .A6(n4059), .Y(io_imem_req_bits_pc[19]) );
  INVX1_LVT U10691 ( .A(n9486), .Y(n9360) );
  AO222X1_LVT U10692 ( .A1(n4066), .A2(csr_io_evec[20]), .A3(n4063), .A4(
        csr_io_pc[20]), .A5(n9360), .A6(n4059), .Y(io_imem_req_bits_pc[20]) );
  AO222X1_LVT U10693 ( .A1(n4066), .A2(csr_io_evec[21]), .A3(n4063), .A4(
        csr_io_pc[21]), .A5(n9361), .A6(n4059), .Y(io_imem_req_bits_pc[21]) );
  INVX1_LVT U10694 ( .A(n9501), .Y(n9362) );
  AO222X1_LVT U10695 ( .A1(n4066), .A2(csr_io_evec[22]), .A3(n4063), .A4(
        csr_io_pc[22]), .A5(n9362), .A6(n4060), .Y(io_imem_req_bits_pc[22]) );
  INVX1_LVT U10696 ( .A(n9488), .Y(n9363) );
  AO222X1_LVT U10697 ( .A1(n4066), .A2(csr_io_evec[23]), .A3(n4063), .A4(
        csr_io_pc[23]), .A5(n9363), .A6(n4060), .Y(io_imem_req_bits_pc[23]) );
  AO222X1_LVT U10698 ( .A1(n4066), .A2(csr_io_evec[24]), .A3(n4063), .A4(
        csr_io_pc[24]), .A5(n9364), .A6(n4060), .Y(io_imem_req_bits_pc[24]) );
  INVX1_LVT U10699 ( .A(n9497), .Y(n9365) );
  AO222X1_LVT U10700 ( .A1(n4066), .A2(csr_io_evec[25]), .A3(n4063), .A4(
        csr_io_pc[25]), .A5(n9365), .A6(n4060), .Y(io_imem_req_bits_pc[25]) );
  INVX1_LVT U10701 ( .A(n9483), .Y(n9366) );
  AO222X1_LVT U10702 ( .A1(n4066), .A2(csr_io_evec[26]), .A3(n4063), .A4(
        csr_io_pc[26]), .A5(n9366), .A6(n4060), .Y(io_imem_req_bits_pc[26]) );
  INVX1_LVT U10703 ( .A(n9489), .Y(n9367) );
  AO222X1_LVT U10704 ( .A1(n4066), .A2(csr_io_evec[27]), .A3(n4063), .A4(
        csr_io_pc[27]), .A5(n9367), .A6(n4060), .Y(io_imem_req_bits_pc[27]) );
  AO222X1_LVT U10705 ( .A1(n4066), .A2(csr_io_evec[28]), .A3(n4062), .A4(
        csr_io_pc[28]), .A5(n9368), .A6(n4060), .Y(io_imem_req_bits_pc[28]) );
  INVX1_LVT U10706 ( .A(n9504), .Y(n9369) );
  AO222X1_LVT U10707 ( .A1(n4066), .A2(csr_io_evec[29]), .A3(n4062), .A4(
        csr_io_pc[29]), .A5(n9369), .A6(n4060), .Y(io_imem_req_bits_pc[29]) );
  INVX1_LVT U10708 ( .A(n9502), .Y(n9370) );
  AO222X1_LVT U10709 ( .A1(n4066), .A2(csr_io_evec[31]), .A3(n4062), .A4(
        csr_io_pc[31]), .A5(n9370), .A6(n4060), .Y(io_imem_req_bits_pc[31]) );
  INVX1_LVT U10710 ( .A(n9505), .Y(n9371) );
  AO222X1_LVT U10711 ( .A1(n4066), .A2(csr_io_evec[32]), .A3(n4062), .A4(
        csr_io_pc[32]), .A5(n9371), .A6(n4060), .Y(io_imem_req_bits_pc[32]) );
  INVX1_LVT U10712 ( .A(n9493), .Y(n9372) );
  AO222X1_LVT U10713 ( .A1(n4066), .A2(csr_io_evec[33]), .A3(n4062), .A4(
        csr_io_pc[33]), .A5(n9372), .A6(n4061), .Y(io_imem_req_bits_pc[33]) );
  AO222X1_LVT U10714 ( .A1(n4066), .A2(csr_io_evec[35]), .A3(n4062), .A4(
        csr_io_pc[35]), .A5(n9374), .A6(n4061), .Y(io_imem_req_bits_pc[35]) );
  INVX1_LVT U10715 ( .A(n9494), .Y(n9375) );
  AO222X1_LVT U10716 ( .A1(n4066), .A2(csr_io_evec[37]), .A3(n4062), .A4(
        csr_io_pc[37]), .A5(n9375), .A6(n4061), .Y(io_imem_req_bits_pc[37]) );
  INVX1_LVT U10717 ( .A(n9498), .Y(n9376) );
  AO222X1_LVT U10718 ( .A1(n4065), .A2(csr_io_evec[38]), .A3(n4062), .A4(
        csr_io_pc[38]), .A5(n9376), .A6(n4061), .Y(io_imem_req_bits_pc[38]) );
  OR2X1_LVT U10719 ( .A1(reset), .A2(n9379), .Y(N778) );
  AND3X1_LVT U10720 ( .A1(ex_ctrl_mem), .A2(N290), .A3(ex_ctrl_rxs2), .Y(N526)
         );
  NAND2X0_LVT U10721 ( .A1(n9417), .A2(n1822), .Y(n9384) );
  NAND2X0_LVT U10722 ( .A1(n9385), .A2(n9384), .Y(n_T_760) );
  AND2X1_LVT U10723 ( .A1(n9389), .A2(n2133), .Y(n9404) );
  AND2X1_LVT U10724 ( .A1(n9394), .A2(n9404), .Y(N238) );
  AND2X1_LVT U10725 ( .A1(n9394), .A2(n9405), .Y(N239) );
  AND2X1_LVT U10726 ( .A1(n9389), .A2(n9392), .Y(n9406) );
  AND2X1_LVT U10727 ( .A1(n9394), .A2(n9406), .Y(N240) );
  AND2X1_LVT U10728 ( .A1(n3042), .A2(n2574), .Y(n9391) );
  AND2X1_LVT U10729 ( .A1(n9391), .A2(n2133), .Y(n9407) );
  AND2X1_LVT U10730 ( .A1(n9394), .A2(n9407), .Y(N241) );
  AND2X1_LVT U10731 ( .A1(n9393), .A2(n2133), .Y(n9408) );
  AND2X1_LVT U10732 ( .A1(n9394), .A2(n9408), .Y(N242) );
  AND2X1_LVT U10733 ( .A1(n9391), .A2(n9392), .Y(n9409) );
  AND2X1_LVT U10734 ( .A1(n9394), .A2(n9409), .Y(N243) );
  AND2X1_LVT U10735 ( .A1(n9393), .A2(n9392), .Y(n9411) );
  AND2X1_LVT U10736 ( .A1(n9394), .A2(n9411), .Y(N244) );
  AND2X1_LVT U10737 ( .A1(n9396), .A2(n2150), .Y(N245) );
  AND2X1_LVT U10738 ( .A1(n9404), .A2(n9396), .Y(N246) );
  AND2X1_LVT U10739 ( .A1(n9405), .A2(n9396), .Y(N247) );
  AND2X1_LVT U10740 ( .A1(n9406), .A2(n9396), .Y(N248) );
  AND2X1_LVT U10741 ( .A1(n9407), .A2(n9396), .Y(N249) );
  AND2X1_LVT U10742 ( .A1(n9408), .A2(n9396), .Y(N250) );
  AND2X1_LVT U10743 ( .A1(n9409), .A2(n9396), .Y(N251) );
  AND2X1_LVT U10744 ( .A1(n9411), .A2(n9396), .Y(N252) );
  AND2X1_LVT U10745 ( .A1(n9401), .A2(n2150), .Y(N253) );
  AND2X1_LVT U10746 ( .A1(n9404), .A2(n9401), .Y(N254) );
  AND2X1_LVT U10747 ( .A1(n9401), .A2(n9405), .Y(N255) );
  AND2X1_LVT U10748 ( .A1(n9406), .A2(n9401), .Y(N256) );
  AND2X1_LVT U10749 ( .A1(n9407), .A2(n9401), .Y(N257) );
  AND2X1_LVT U10750 ( .A1(n9408), .A2(n9401), .Y(N258) );
  AND2X1_LVT U10751 ( .A1(n9409), .A2(n9401), .Y(N259) );
  AND2X1_LVT U10752 ( .A1(n9411), .A2(n9401), .Y(N260) );
  AND2X1_LVT U10753 ( .A1(n9410), .A2(n2150), .Y(N261) );
  AND2X1_LVT U10754 ( .A1(n9404), .A2(n9410), .Y(N262) );
  AND2X1_LVT U10755 ( .A1(n9410), .A2(n9405), .Y(N263) );
  AND2X1_LVT U10756 ( .A1(n9406), .A2(n9410), .Y(N264) );
  AND2X1_LVT U10757 ( .A1(n9407), .A2(n9410), .Y(N265) );
  AND2X1_LVT U10758 ( .A1(n9408), .A2(n9410), .Y(N266) );
  AND2X1_LVT U10759 ( .A1(n9409), .A2(n9410), .Y(N267) );
  AND2X1_LVT U10760 ( .A1(n9411), .A2(n9410), .Y(N268) );
  NAND2X0_LVT U10761 ( .A1(n9426), .A2(n9449), .Y(N271) );
  AOI22X1_LVT U10764 ( .A1(n_T_698[14]), .A2(n9506), .A3(n_T_698[8]), .A4(
        n9511), .Y(n9450) );
  AOI22X1_LVT U10765 ( .A1(n_T_698[12]), .A2(n9491), .A3(n_T_698[29]), .A4(
        n9504), .Y(n9451) );
  AOI22X1_LVT U10766 ( .A1(n_T_698[32]), .A2(n9505), .A3(n_T_698[27]), .A4(
        n9489), .Y(n9452) );
  AOI22X1_LVT U10767 ( .A1(n_T_698[6]), .A2(n9485), .A3(n_T_698[9]), .A4(n9507), .Y(n9453) );
  NAND4X0_LVT U10768 ( .A1(n_T_918[59]), .A2(n_T_918[48]), .A3(n_T_918[62]), 
        .A4(n_T_918[56]), .Y(n9469) );
  AND4X1_LVT U10769 ( .A1(n_T_918[39]), .A2(n_T_918[40]), .A3(n_T_918[47]), 
        .A4(n_T_918[60]), .Y(n9459) );
  NAND4X0_LVT U10770 ( .A1(n_T_918[55]), .A2(n_T_918[58]), .A3(n_T_918[44]), 
        .A4(n_T_918[43]), .Y(n9457) );
  NAND4X0_LVT U10771 ( .A1(n_T_918[49]), .A2(n_T_918[45]), .A3(n_T_918[61]), 
        .A4(n_T_918[57]), .Y(n9456) );
  NAND4X0_LVT U10772 ( .A1(n_T_918[41]), .A2(n_T_918[53]), .A3(n_T_918[54]), 
        .A4(n_T_918[50]), .Y(n9455) );
  NAND4X0_LVT U10773 ( .A1(n_T_918[63]), .A2(n_T_918[46]), .A3(n_T_918[42]), 
        .A4(n_T_918[52]), .Y(n9454) );
  NAND3X0_LVT U10774 ( .A1(n_T_918[51]), .A2(n9459), .A3(n9458), .Y(n9468) );
  NAND4X0_LVT U10775 ( .A1(n9463), .A2(n9462), .A3(n9461), .A4(n9460), .Y(
        n9467) );
  NAND3X0_LVT U10776 ( .A1(n9465), .A2(n9464), .A3(n3249), .Y(n9466) );
  OA22X1_LVT U10777 ( .A1(n9469), .A2(n9468), .A3(n9467), .A4(n9466), .Y(n9470) );
  AOI22X1_LVT U10778 ( .A1(n_T_698[3]), .A2(n9503), .A3(n_T_698[18]), .A4(
        n9496), .Y(n9471) );
  AOI22X1_LVT U10779 ( .A1(n_T_698[10]), .A2(n9509), .A3(n_T_698[13]), .A4(
        n9500), .Y(n9472) );
  OAI22X1_LVT U10780 ( .A1(n_T_698[38]), .A2(n9498), .A3(n_T_698[36]), .A4(
        n9508), .Y(n9473) );
  AO221X1_LVT U10781 ( .A1(n9498), .A2(n_T_698[38]), .A3(n_T_698[36]), .A4(
        n9508), .A5(n9473), .Y(n9482) );
  AOI22X1_LVT U10782 ( .A1(n_T_698[33]), .A2(n9493), .A3(n_T_698[5]), .A4(
        n9484), .Y(n9474) );
  OA221X1_LVT U10783 ( .A1(n_T_698[33]), .A2(n9493), .A3(n_T_698[5]), .A4(
        n9484), .A5(n9474), .Y(n9481) );
  AOI22X1_LVT U10784 ( .A1(n_T_698[37]), .A2(n9494), .A3(n_T_698[30]), .A4(
        n9492), .Y(n9475) );
  OA221X1_LVT U10785 ( .A1(n_T_698[37]), .A2(n9494), .A3(n_T_698[30]), .A4(
        n9492), .A5(n9475), .Y(n9480) );
  AOI22X1_LVT U10786 ( .A1(n_T_698[26]), .A2(n9483), .A3(n_T_698[20]), .A4(
        n9486), .Y(n9476) );
  OA221X1_LVT U10787 ( .A1(n_T_698[26]), .A2(n9483), .A3(n_T_698[20]), .A4(
        n9486), .A5(n9476), .Y(n9479) );
  AOI22X1_LVT U10788 ( .A1(n_T_698[11]), .A2(n9490), .A3(n_T_698[17]), .A4(
        n9487), .Y(n9477) );
  OA221X1_LVT U10789 ( .A1(n_T_698[11]), .A2(n9490), .A3(n_T_698[17]), .A4(
        n9487), .A5(n9477), .Y(n9478) );
  NAND2X0_LVT U10790 ( .A1(n555), .A2(n3104), .Y(n9514) );
  AND2X1_LVT U10791 ( .A1(n3202), .A2(n9514), .Y(
        io_imem_btb_update_bits_cfiType[0]) );
  AO22X1_LVT U10792 ( .A1(n_T_849[11]), .A2(n9514), .A3(n_T_904[3]), .A4(n9513), .Y(io_imem_btb_update_bits_cfiType[1]) );
  OR2X1_LVT U10793 ( .A1(io_imem_bht_update_bits_branch), .A2(n9514), .Y(
        io_imem_btb_update_bits_isValid) );
endmodule

